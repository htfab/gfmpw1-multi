magic
tech gf180mcuD
magscale 1 10
timestamp 1702448400
<< metal1 >>
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 1344 55466 58576 55500
rect 1344 55414 4478 55466
rect 4530 55414 4582 55466
rect 4634 55414 4686 55466
rect 4738 55414 35198 55466
rect 35250 55414 35302 55466
rect 35354 55414 35406 55466
rect 35458 55414 58576 55466
rect 1344 55380 58576 55414
rect 1344 54458 58576 54492
rect 1344 54406 19838 54458
rect 19890 54406 19942 54458
rect 19994 54406 20046 54458
rect 20098 54406 50558 54458
rect 50610 54406 50662 54458
rect 50714 54406 50766 54458
rect 50818 54406 58576 54458
rect 1344 54372 58576 54406
rect 55246 54178 55298 54190
rect 55246 54114 55298 54126
rect 1344 53450 58576 53484
rect 1344 53398 4478 53450
rect 4530 53398 4582 53450
rect 4634 53398 4686 53450
rect 4738 53398 35198 53450
rect 35250 53398 35302 53450
rect 35354 53398 35406 53450
rect 35458 53398 58576 53450
rect 1344 53364 58576 53398
rect 1344 52442 58576 52476
rect 1344 52390 19838 52442
rect 19890 52390 19942 52442
rect 19994 52390 20046 52442
rect 20098 52390 50558 52442
rect 50610 52390 50662 52442
rect 50714 52390 50766 52442
rect 50818 52390 58576 52442
rect 1344 52356 58576 52390
rect 5854 52162 5906 52174
rect 5854 52098 5906 52110
rect 1344 51434 58576 51468
rect 1344 51382 4478 51434
rect 4530 51382 4582 51434
rect 4634 51382 4686 51434
rect 4738 51382 35198 51434
rect 35250 51382 35302 51434
rect 35354 51382 35406 51434
rect 35458 51382 58576 51434
rect 1344 51348 58576 51382
rect 1344 50426 58576 50460
rect 1344 50374 19838 50426
rect 19890 50374 19942 50426
rect 19994 50374 20046 50426
rect 20098 50374 50558 50426
rect 50610 50374 50662 50426
rect 50714 50374 50766 50426
rect 50818 50374 58576 50426
rect 1344 50340 58576 50374
rect 36990 49810 37042 49822
rect 36990 49746 37042 49758
rect 41358 49810 41410 49822
rect 41358 49746 41410 49758
rect 41806 49810 41858 49822
rect 41806 49746 41858 49758
rect 42254 49810 42306 49822
rect 42254 49746 42306 49758
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 41694 49026 41746 49038
rect 41694 48962 41746 48974
rect 31278 48914 31330 48926
rect 31278 48850 31330 48862
rect 32734 48914 32786 48926
rect 32734 48850 32786 48862
rect 30830 48802 30882 48814
rect 30830 48738 30882 48750
rect 31950 48802 32002 48814
rect 31950 48738 32002 48750
rect 37438 48802 37490 48814
rect 37438 48738 37490 48750
rect 40798 48802 40850 48814
rect 40798 48738 40850 48750
rect 41246 48802 41298 48814
rect 41246 48738 41298 48750
rect 42142 48802 42194 48814
rect 42142 48738 42194 48750
rect 42366 48802 42418 48814
rect 42366 48738 42418 48750
rect 36430 48690 36482 48702
rect 34850 48638 34862 48690
rect 34914 48638 34926 48690
rect 36430 48626 36482 48638
rect 38110 48690 38162 48702
rect 38110 48626 38162 48638
rect 40126 48690 40178 48702
rect 40126 48626 40178 48638
rect 43374 48690 43426 48702
rect 43374 48626 43426 48638
rect 44158 48690 44210 48702
rect 44158 48626 44210 48638
rect 1344 48410 58576 48444
rect 1344 48358 19838 48410
rect 19890 48358 19942 48410
rect 19994 48358 20046 48410
rect 20098 48358 50558 48410
rect 50610 48358 50662 48410
rect 50714 48358 50766 48410
rect 50818 48358 58576 48410
rect 1344 48324 58576 48358
rect 41806 48130 41858 48142
rect 6178 48078 6190 48130
rect 6242 48078 6254 48130
rect 41806 48066 41858 48078
rect 43710 48130 43762 48142
rect 43710 48066 43762 48078
rect 37102 48018 37154 48030
rect 42814 48018 42866 48030
rect 39330 47966 39342 48018
rect 39394 47966 39406 48018
rect 37102 47954 37154 47966
rect 42814 47954 42866 47966
rect 3390 47906 3442 47918
rect 26014 47906 26066 47918
rect 3938 47854 3950 47906
rect 4002 47854 4014 47906
rect 3390 47842 3442 47854
rect 26014 47842 26066 47854
rect 26574 47906 26626 47918
rect 26574 47842 26626 47854
rect 36766 47906 36818 47918
rect 36766 47842 36818 47854
rect 40350 47906 40402 47918
rect 43486 47906 43538 47918
rect 40786 47854 40798 47906
rect 40850 47903 40862 47906
rect 41458 47903 41470 47906
rect 40850 47857 41470 47903
rect 40850 47854 40862 47857
rect 41458 47854 41470 47857
rect 41522 47854 41534 47906
rect 40350 47842 40402 47854
rect 43486 47842 43538 47854
rect 3054 47794 3106 47806
rect 3054 47730 3106 47742
rect 24670 47794 24722 47806
rect 24670 47730 24722 47742
rect 25566 47794 25618 47806
rect 35422 47794 35474 47806
rect 28690 47742 28702 47794
rect 28754 47742 28766 47794
rect 25566 47730 25618 47742
rect 35422 47730 35474 47742
rect 35870 47794 35922 47806
rect 35870 47730 35922 47742
rect 36318 47794 36370 47806
rect 36318 47730 36370 47742
rect 6514 47630 6526 47682
rect 6578 47630 6590 47682
rect 35410 47518 35422 47570
rect 35474 47567 35486 47570
rect 35858 47567 35870 47570
rect 35474 47521 35870 47567
rect 35474 47518 35486 47521
rect 35858 47518 35870 47521
rect 35922 47567 35934 47570
rect 36642 47567 36654 47570
rect 35922 47521 36654 47567
rect 35922 47518 35934 47521
rect 36642 47518 36654 47521
rect 36706 47518 36718 47570
rect 1344 47402 58576 47436
rect 1344 47350 4478 47402
rect 4530 47350 4582 47402
rect 4634 47350 4686 47402
rect 4738 47350 35198 47402
rect 35250 47350 35302 47402
rect 35354 47350 35406 47402
rect 35458 47350 58576 47402
rect 1344 47316 58576 47350
rect 34850 47182 34862 47234
rect 34914 47182 34926 47234
rect 6290 47119 6302 47122
rect 5969 47073 6302 47119
rect 5630 47010 5682 47022
rect 5730 46958 5742 47010
rect 5794 47007 5806 47010
rect 5969 47007 6015 47073
rect 6290 47070 6302 47073
rect 6354 47070 6366 47122
rect 38658 47070 38670 47122
rect 38722 47119 38734 47122
rect 39442 47119 39454 47122
rect 38722 47073 39454 47119
rect 38722 47070 38734 47073
rect 39442 47070 39454 47073
rect 39506 47119 39518 47122
rect 40002 47119 40014 47122
rect 39506 47073 40014 47119
rect 39506 47070 39518 47073
rect 40002 47070 40014 47073
rect 40066 47070 40078 47122
rect 5794 46961 6015 47007
rect 39454 47010 39506 47022
rect 5794 46958 5806 46961
rect 5630 46946 5682 46958
rect 39454 46946 39506 46958
rect 25006 46898 25058 46910
rect 5730 46846 5742 46898
rect 5794 46846 5806 46898
rect 22530 46846 22542 46898
rect 22594 46846 22606 46898
rect 22978 46846 22990 46898
rect 23042 46846 23054 46898
rect 25006 46834 25058 46846
rect 39006 46898 39058 46910
rect 39006 46834 39058 46846
rect 40238 46898 40290 46910
rect 40238 46834 40290 46846
rect 40686 46898 40738 46910
rect 40686 46834 40738 46846
rect 30494 46786 30546 46798
rect 31490 46734 31502 46786
rect 31554 46734 31566 46786
rect 30494 46722 30546 46734
rect 6190 46674 6242 46686
rect 6190 46610 6242 46622
rect 21646 46674 21698 46686
rect 21646 46610 21698 46622
rect 22094 46674 22146 46686
rect 22094 46610 22146 46622
rect 25790 46674 25842 46686
rect 25790 46610 25842 46622
rect 26350 46674 26402 46686
rect 26350 46610 26402 46622
rect 27582 46674 27634 46686
rect 27582 46610 27634 46622
rect 29262 46674 29314 46686
rect 29262 46610 29314 46622
rect 29710 46674 29762 46686
rect 29710 46610 29762 46622
rect 30158 46674 30210 46686
rect 30158 46610 30210 46622
rect 39902 46674 39954 46686
rect 39902 46610 39954 46622
rect 42926 46674 42978 46686
rect 42926 46610 42978 46622
rect 29250 46510 29262 46562
rect 29314 46559 29326 46562
rect 30146 46559 30158 46562
rect 29314 46513 30158 46559
rect 29314 46510 29326 46513
rect 30146 46510 30158 46513
rect 30210 46510 30222 46562
rect 38882 46510 38894 46562
rect 38946 46559 38958 46562
rect 39890 46559 39902 46562
rect 38946 46513 39902 46559
rect 38946 46510 38958 46513
rect 39890 46510 39902 46513
rect 39954 46510 39966 46562
rect 44034 46510 44046 46562
rect 44098 46510 44110 46562
rect 1344 46394 58576 46428
rect 1344 46342 19838 46394
rect 19890 46342 19942 46394
rect 19994 46342 20046 46394
rect 20098 46342 50558 46394
rect 50610 46342 50662 46394
rect 50714 46342 50766 46394
rect 50818 46342 58576 46394
rect 1344 46308 58576 46342
rect 7198 46114 7250 46126
rect 7198 46050 7250 46062
rect 27806 46114 27858 46126
rect 27806 46050 27858 46062
rect 30942 46114 30994 46126
rect 30942 46050 30994 46062
rect 41134 46114 41186 46126
rect 41134 46050 41186 46062
rect 41582 46114 41634 46126
rect 41582 46050 41634 46062
rect 28590 46002 28642 46014
rect 28590 45938 28642 45950
rect 4510 45890 4562 45902
rect 28142 45890 28194 45902
rect 5058 45838 5070 45890
rect 5122 45838 5134 45890
rect 8418 45838 8430 45890
rect 8482 45838 8494 45890
rect 11666 45838 11678 45890
rect 11730 45838 11742 45890
rect 4510 45826 4562 45838
rect 28142 45826 28194 45838
rect 35086 45890 35138 45902
rect 35086 45826 35138 45838
rect 35870 45890 35922 45902
rect 36418 45838 36430 45890
rect 36482 45838 36494 45890
rect 38546 45838 38558 45890
rect 38610 45838 38622 45890
rect 46050 45838 46062 45890
rect 46114 45838 46126 45890
rect 48178 45838 48190 45890
rect 48242 45838 48254 45890
rect 35870 45826 35922 45838
rect 1822 45778 1874 45790
rect 1822 45714 1874 45726
rect 4174 45778 4226 45790
rect 4174 45714 4226 45726
rect 9662 45778 9714 45790
rect 9662 45714 9714 45726
rect 26462 45778 26514 45790
rect 26462 45714 26514 45726
rect 26910 45778 26962 45790
rect 26910 45714 26962 45726
rect 27358 45778 27410 45790
rect 27358 45714 27410 45726
rect 33182 45778 33234 45790
rect 33182 45714 33234 45726
rect 34638 45778 34690 45790
rect 34638 45714 34690 45726
rect 35534 45778 35586 45790
rect 35534 45714 35586 45726
rect 7634 45614 7646 45666
rect 7698 45614 7710 45666
rect 26562 45614 26574 45666
rect 26626 45663 26638 45666
rect 26898 45663 26910 45666
rect 26626 45617 26910 45663
rect 26626 45614 26638 45617
rect 26898 45614 26910 45617
rect 26962 45663 26974 45666
rect 27346 45663 27358 45666
rect 26962 45617 27358 45663
rect 26962 45614 26974 45617
rect 27346 45614 27358 45617
rect 27410 45663 27422 45666
rect 28130 45663 28142 45666
rect 27410 45617 28142 45663
rect 27410 45614 27422 45617
rect 28130 45614 28142 45617
rect 28194 45614 28206 45666
rect 31826 45614 31838 45666
rect 31890 45614 31902 45666
rect 40002 45614 40014 45666
rect 40066 45614 40078 45666
rect 43138 45614 43150 45666
rect 43202 45614 43214 45666
rect 8306 45502 8318 45554
rect 8370 45502 8382 45554
rect 11554 45502 11566 45554
rect 11618 45502 11630 45554
rect 1344 45386 58576 45420
rect 1344 45334 4478 45386
rect 4530 45334 4582 45386
rect 4634 45334 4686 45386
rect 4738 45334 35198 45386
rect 35250 45334 35302 45386
rect 35354 45334 35406 45386
rect 35458 45334 58576 45386
rect 1344 45300 58576 45334
rect 5618 45166 5630 45218
rect 5682 45166 5694 45218
rect 22082 45166 22094 45218
rect 22146 45215 22158 45218
rect 22978 45215 22990 45218
rect 22146 45169 22990 45215
rect 22146 45166 22158 45169
rect 22978 45166 22990 45169
rect 23042 45166 23054 45218
rect 12786 45054 12798 45106
rect 12850 45054 12862 45106
rect 22206 44994 22258 45006
rect 22206 44930 22258 44942
rect 28590 44994 28642 45006
rect 28590 44930 28642 44942
rect 37662 44994 37714 45006
rect 37662 44930 37714 44942
rect 1822 44882 1874 44894
rect 6078 44882 6130 44894
rect 9662 44882 9714 44894
rect 23438 44882 23490 44894
rect 26350 44882 26402 44894
rect 29486 44882 29538 44894
rect 2370 44830 2382 44882
rect 2434 44830 2446 44882
rect 5730 44830 5742 44882
rect 5794 44830 5806 44882
rect 6626 44830 6638 44882
rect 6690 44830 6702 44882
rect 10210 44830 10222 44882
rect 10274 44830 10286 44882
rect 23986 44830 23998 44882
rect 24050 44830 24062 44882
rect 26674 44830 26686 44882
rect 26738 44830 26750 44882
rect 1822 44818 1874 44830
rect 6078 44818 6130 44830
rect 9662 44818 9714 44830
rect 23438 44818 23490 44830
rect 26350 44818 26402 44830
rect 29486 44818 29538 44830
rect 29934 44882 29986 44894
rect 29934 44818 29986 44830
rect 30270 44882 30322 44894
rect 33182 44882 33234 44894
rect 45614 44882 45666 44894
rect 32610 44830 32622 44882
rect 32674 44830 32686 44882
rect 41458 44830 41470 44882
rect 41522 44830 41534 44882
rect 30270 44818 30322 44830
rect 33182 44818 33234 44830
rect 45614 44818 45666 44830
rect 38334 44770 38386 44782
rect 38334 44706 38386 44718
rect 46510 44770 46562 44782
rect 46510 44706 46562 44718
rect 47294 44770 47346 44782
rect 47294 44706 47346 44718
rect 4510 44658 4562 44670
rect 4510 44594 4562 44606
rect 4958 44658 5010 44670
rect 4958 44594 5010 44606
rect 8766 44658 8818 44670
rect 8766 44594 8818 44606
rect 9214 44658 9266 44670
rect 9214 44594 9266 44606
rect 12350 44658 12402 44670
rect 12350 44594 12402 44606
rect 22654 44658 22706 44670
rect 22654 44594 22706 44606
rect 23102 44658 23154 44670
rect 23102 44594 23154 44606
rect 33630 44658 33682 44670
rect 33630 44594 33682 44606
rect 35646 44658 35698 44670
rect 35646 44594 35698 44606
rect 36430 44658 36482 44670
rect 36430 44594 36482 44606
rect 37214 44658 37266 44670
rect 37214 44594 37266 44606
rect 38894 44658 38946 44670
rect 38894 44594 38946 44606
rect 41134 44658 41186 44670
rect 41134 44594 41186 44606
rect 42254 44658 42306 44670
rect 42254 44594 42306 44606
rect 45166 44658 45218 44670
rect 45166 44594 45218 44606
rect 27794 44494 27806 44546
rect 27858 44494 27870 44546
rect 1344 44378 58576 44412
rect 1344 44326 19838 44378
rect 19890 44326 19942 44378
rect 19994 44326 20046 44378
rect 20098 44326 50558 44378
rect 50610 44326 50662 44378
rect 50714 44326 50766 44378
rect 50818 44326 58576 44378
rect 1344 44292 58576 44326
rect 10210 44158 10222 44210
rect 10274 44158 10286 44210
rect 1822 44098 1874 44110
rect 1822 44034 1874 44046
rect 4846 44098 4898 44110
rect 8878 44098 8930 44110
rect 8530 44046 8542 44098
rect 8594 44046 8606 44098
rect 4846 44034 4898 44046
rect 8878 44034 8930 44046
rect 9886 44098 9938 44110
rect 9886 44034 9938 44046
rect 10334 44098 10386 44110
rect 10334 44034 10386 44046
rect 13582 44098 13634 44110
rect 13582 44034 13634 44046
rect 27246 44098 27298 44110
rect 27246 44034 27298 44046
rect 33294 44098 33346 44110
rect 33294 44034 33346 44046
rect 35646 44098 35698 44110
rect 35646 44034 35698 44046
rect 38894 44098 38946 44110
rect 38894 44034 38946 44046
rect 43710 44098 43762 44110
rect 43710 44034 43762 44046
rect 45390 44098 45442 44110
rect 45390 44034 45442 44046
rect 48190 44098 48242 44110
rect 48190 44034 48242 44046
rect 14478 43986 14530 43998
rect 14478 43922 14530 43934
rect 18174 43986 18226 43998
rect 18174 43922 18226 43934
rect 27694 43986 27746 43998
rect 27694 43922 27746 43934
rect 28814 43986 28866 43998
rect 28814 43922 28866 43934
rect 34302 43986 34354 43998
rect 34302 43922 34354 43934
rect 35086 43986 35138 43998
rect 35086 43922 35138 43934
rect 40910 43986 40962 43998
rect 40910 43922 40962 43934
rect 41582 43986 41634 43998
rect 41582 43922 41634 43934
rect 43038 43986 43090 43998
rect 43038 43922 43090 43934
rect 2158 43874 2210 43886
rect 5742 43874 5794 43886
rect 10894 43874 10946 43886
rect 17390 43874 17442 43886
rect 2706 43822 2718 43874
rect 2770 43822 2782 43874
rect 6290 43822 6302 43874
rect 6354 43822 6366 43874
rect 11442 43822 11454 43874
rect 11506 43822 11518 43874
rect 14578 43822 14590 43874
rect 14642 43822 14654 43874
rect 2158 43810 2210 43822
rect 5742 43810 5794 43822
rect 10894 43810 10946 43822
rect 17390 43810 17442 43822
rect 28142 43874 28194 43886
rect 28142 43810 28194 43822
rect 33518 43874 33570 43886
rect 33518 43810 33570 43822
rect 36206 43874 36258 43886
rect 41246 43874 41298 43886
rect 36754 43822 36766 43874
rect 36818 43822 36830 43874
rect 36206 43810 36258 43822
rect 41246 43810 41298 43822
rect 41918 43874 41970 43886
rect 41918 43810 41970 43822
rect 42478 43874 42530 43886
rect 54114 43822 54126 43874
rect 54178 43822 54190 43874
rect 42478 43810 42530 43822
rect 16830 43762 16882 43774
rect 16830 43698 16882 43710
rect 20190 43762 20242 43774
rect 20190 43698 20242 43710
rect 32286 43762 32338 43774
rect 32286 43698 32338 43710
rect 45726 43762 45778 43774
rect 45726 43698 45778 43710
rect 46958 43762 47010 43774
rect 46958 43698 47010 43710
rect 47406 43762 47458 43774
rect 51762 43710 51774 43762
rect 51826 43710 51838 43762
rect 47406 43698 47458 43710
rect 5282 43598 5294 43650
rect 5346 43598 5358 43650
rect 14018 43598 14030 43650
rect 14082 43598 14094 43650
rect 31378 43598 31390 43650
rect 31442 43598 31454 43650
rect 39330 43598 39342 43650
rect 39394 43598 39406 43650
rect 1344 43370 58576 43404
rect 1344 43318 4478 43370
rect 4530 43318 4582 43370
rect 4634 43318 4686 43370
rect 4738 43318 35198 43370
rect 35250 43318 35302 43370
rect 35354 43318 35406 43370
rect 35458 43318 58576 43370
rect 1344 43284 58576 43318
rect 5618 43150 5630 43202
rect 5682 43150 5694 43202
rect 6066 43150 6078 43202
rect 6130 43150 6142 43202
rect 13458 43150 13470 43202
rect 13522 43150 13534 43202
rect 12786 43038 12798 43090
rect 12850 43038 12862 43090
rect 35870 42978 35922 42990
rect 35870 42914 35922 42926
rect 37102 42978 37154 42990
rect 37102 42914 37154 42926
rect 37886 42978 37938 42990
rect 37886 42914 37938 42926
rect 46734 42978 46786 42990
rect 46734 42914 46786 42926
rect 48078 42978 48130 42990
rect 48078 42914 48130 42926
rect 1822 42866 1874 42878
rect 9662 42866 9714 42878
rect 17054 42866 17106 42878
rect 2370 42814 2382 42866
rect 2434 42814 2446 42866
rect 5730 42814 5742 42866
rect 5794 42814 5806 42866
rect 6178 42814 6190 42866
rect 6242 42814 6254 42866
rect 10210 42814 10222 42866
rect 10274 42814 10286 42866
rect 13570 42814 13582 42866
rect 13634 42814 13646 42866
rect 1822 42802 1874 42814
rect 9662 42802 9714 42814
rect 17054 42802 17106 42814
rect 19854 42866 19906 42878
rect 19854 42802 19906 42814
rect 23774 42866 23826 42878
rect 23774 42802 23826 42814
rect 31726 42866 31778 42878
rect 31726 42802 31778 42814
rect 32398 42866 32450 42878
rect 32398 42802 32450 42814
rect 33854 42866 33906 42878
rect 33854 42802 33906 42814
rect 39678 42866 39730 42878
rect 39678 42802 39730 42814
rect 40350 42866 40402 42878
rect 40350 42802 40402 42814
rect 41806 42866 41858 42878
rect 41806 42802 41858 42814
rect 47966 42866 48018 42878
rect 47966 42802 48018 42814
rect 48190 42866 48242 42878
rect 48190 42802 48242 42814
rect 22318 42754 22370 42766
rect 22318 42690 22370 42702
rect 22542 42754 22594 42766
rect 22542 42690 22594 42702
rect 22766 42754 22818 42766
rect 22766 42690 22818 42702
rect 23438 42754 23490 42766
rect 23438 42690 23490 42702
rect 32062 42754 32114 42766
rect 32062 42690 32114 42702
rect 33294 42754 33346 42766
rect 33294 42690 33346 42702
rect 34526 42754 34578 42766
rect 34526 42690 34578 42702
rect 35310 42754 35362 42766
rect 35310 42690 35362 42702
rect 40014 42754 40066 42766
rect 42478 42754 42530 42766
rect 41122 42702 41134 42754
rect 41186 42702 41198 42754
rect 40014 42690 40066 42702
rect 42478 42690 42530 42702
rect 47518 42754 47570 42766
rect 47518 42690 47570 42702
rect 47742 42754 47794 42766
rect 47742 42690 47794 42702
rect 4958 42642 5010 42654
rect 4610 42590 4622 42642
rect 4674 42590 4686 42642
rect 4958 42578 5010 42590
rect 6638 42642 6690 42654
rect 6638 42578 6690 42590
rect 9326 42642 9378 42654
rect 9326 42578 9378 42590
rect 12350 42642 12402 42654
rect 12350 42578 12402 42590
rect 16718 42642 16770 42654
rect 16718 42578 16770 42590
rect 17838 42642 17890 42654
rect 17838 42578 17890 42590
rect 21422 42642 21474 42654
rect 21422 42578 21474 42590
rect 21870 42642 21922 42654
rect 21870 42578 21922 42590
rect 26350 42642 26402 42654
rect 26350 42578 26402 42590
rect 27358 42642 27410 42654
rect 27358 42578 27410 42590
rect 27806 42642 27858 42654
rect 27806 42578 27858 42590
rect 29374 42642 29426 42654
rect 29374 42578 29426 42590
rect 29822 42642 29874 42654
rect 29822 42578 29874 42590
rect 32734 42642 32786 42654
rect 32734 42578 32786 42590
rect 40686 42642 40738 42654
rect 40686 42578 40738 42590
rect 43934 42642 43986 42654
rect 43934 42578 43986 42590
rect 44942 42642 44994 42654
rect 44942 42578 44994 42590
rect 45390 42642 45442 42654
rect 45390 42578 45442 42590
rect 45838 42642 45890 42654
rect 45838 42578 45890 42590
rect 46286 42642 46338 42654
rect 46286 42578 46338 42590
rect 47182 42642 47234 42654
rect 47182 42578 47234 42590
rect 48638 42642 48690 42654
rect 48638 42578 48690 42590
rect 49086 42642 49138 42654
rect 49086 42578 49138 42590
rect 49534 42642 49586 42654
rect 49534 42578 49586 42590
rect 50878 42642 50930 42654
rect 50878 42578 50930 42590
rect 51214 42642 51266 42654
rect 51214 42578 51266 42590
rect 51662 42642 51714 42654
rect 51662 42578 51714 42590
rect 52110 42642 52162 42654
rect 52110 42578 52162 42590
rect 52782 42642 52834 42654
rect 52782 42578 52834 42590
rect 53342 42642 53394 42654
rect 53342 42578 53394 42590
rect 53790 42642 53842 42654
rect 53790 42578 53842 42590
rect 54238 42642 54290 42654
rect 54238 42578 54290 42590
rect 21858 42478 21870 42530
rect 21922 42527 21934 42530
rect 22418 42527 22430 42530
rect 21922 42481 22430 42527
rect 21922 42478 21934 42481
rect 22418 42478 22430 42481
rect 22482 42478 22494 42530
rect 44930 42478 44942 42530
rect 44994 42527 45006 42530
rect 46274 42527 46286 42530
rect 44994 42481 46286 42527
rect 44994 42478 45006 42481
rect 46274 42478 46286 42481
rect 46338 42527 46350 42530
rect 47282 42527 47294 42530
rect 46338 42481 47294 42527
rect 46338 42478 46350 42481
rect 47282 42478 47294 42481
rect 47346 42478 47358 42530
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 3502 42082 3554 42094
rect 13470 42082 13522 42094
rect 6626 42030 6638 42082
rect 6690 42030 6702 42082
rect 3502 42018 3554 42030
rect 13470 42018 13522 42030
rect 29262 42082 29314 42094
rect 52334 42082 52386 42094
rect 47170 42030 47182 42082
rect 47234 42030 47246 42082
rect 29262 42018 29314 42030
rect 52334 42018 52386 42030
rect 3390 41970 3442 41982
rect 3390 41906 3442 41918
rect 20526 41970 20578 41982
rect 20526 41906 20578 41918
rect 21870 41970 21922 41982
rect 21870 41906 21922 41918
rect 26126 41970 26178 41982
rect 26126 41906 26178 41918
rect 26462 41970 26514 41982
rect 26462 41906 26514 41918
rect 27134 41970 27186 41982
rect 27134 41906 27186 41918
rect 28030 41970 28082 41982
rect 28030 41906 28082 41918
rect 28590 41970 28642 41982
rect 28590 41906 28642 41918
rect 33406 41970 33458 41982
rect 33406 41906 33458 41918
rect 34638 41970 34690 41982
rect 34638 41906 34690 41918
rect 35198 41970 35250 41982
rect 35198 41906 35250 41918
rect 35870 41970 35922 41982
rect 35870 41906 35922 41918
rect 37998 41970 38050 41982
rect 37998 41906 38050 41918
rect 43934 41970 43986 41982
rect 43934 41906 43986 41918
rect 46734 41970 46786 41982
rect 48862 41970 48914 41982
rect 47506 41918 47518 41970
rect 47570 41918 47582 41970
rect 46734 41906 46786 41918
rect 48862 41906 48914 41918
rect 53118 41970 53170 41982
rect 53118 41906 53170 41918
rect 55582 41970 55634 41982
rect 55582 41906 55634 41918
rect 3838 41858 3890 41870
rect 10782 41858 10834 41870
rect 13918 41858 13970 41870
rect 18510 41858 18562 41870
rect 4386 41806 4398 41858
rect 4450 41806 4462 41858
rect 11330 41806 11342 41858
rect 11394 41806 11406 41858
rect 14466 41806 14478 41858
rect 14530 41806 14542 41858
rect 3838 41794 3890 41806
rect 10782 41794 10834 41806
rect 13918 41794 13970 41806
rect 18510 41794 18562 41806
rect 21310 41858 21362 41870
rect 21310 41794 21362 41806
rect 26798 41858 26850 41870
rect 26798 41794 26850 41806
rect 27470 41858 27522 41870
rect 27470 41794 27522 41806
rect 30046 41858 30098 41870
rect 30046 41794 30098 41806
rect 33070 41858 33122 41870
rect 33070 41794 33122 41806
rect 33742 41858 33794 41870
rect 33742 41794 33794 41806
rect 34078 41858 34130 41870
rect 34078 41794 34130 41806
rect 40910 41858 40962 41870
rect 40910 41794 40962 41806
rect 44270 41858 44322 41870
rect 44270 41794 44322 41806
rect 44494 41858 44546 41870
rect 44494 41794 44546 41806
rect 44718 41858 44770 41870
rect 44718 41794 44770 41806
rect 45614 41858 45666 41870
rect 45614 41794 45666 41806
rect 49198 41858 49250 41870
rect 49758 41858 49810 41870
rect 52782 41858 52834 41870
rect 49410 41806 49422 41858
rect 49474 41806 49486 41858
rect 49858 41806 49870 41858
rect 49922 41806 49934 41858
rect 49198 41794 49250 41806
rect 49758 41794 49810 41806
rect 52782 41794 52834 41806
rect 53454 41858 53506 41870
rect 53454 41794 53506 41806
rect 53790 41858 53842 41870
rect 53790 41794 53842 41806
rect 54350 41858 54402 41870
rect 54350 41794 54402 41806
rect 54910 41858 54962 41870
rect 54910 41794 54962 41806
rect 1822 41746 1874 41758
rect 1822 41682 1874 41694
rect 3054 41746 3106 41758
rect 3054 41682 3106 41694
rect 10446 41746 10498 41758
rect 10446 41682 10498 41694
rect 18174 41746 18226 41758
rect 18174 41682 18226 41694
rect 30494 41746 30546 41758
rect 30494 41682 30546 41694
rect 32510 41746 32562 41758
rect 32510 41682 32562 41694
rect 36766 41746 36818 41758
rect 36766 41682 36818 41694
rect 37102 41746 37154 41758
rect 37102 41682 37154 41694
rect 37550 41746 37602 41758
rect 37550 41682 37602 41694
rect 39902 41746 39954 41758
rect 39902 41682 39954 41694
rect 40462 41746 40514 41758
rect 40462 41682 40514 41694
rect 43038 41746 43090 41758
rect 43038 41682 43090 41694
rect 43486 41746 43538 41758
rect 43486 41682 43538 41694
rect 50878 41746 50930 41758
rect 50878 41682 50930 41694
rect 51550 41746 51602 41758
rect 51550 41682 51602 41694
rect 51998 41746 52050 41758
rect 51998 41682 52050 41694
rect 14366 41634 14418 41646
rect 6962 41582 6974 41634
rect 7026 41582 7038 41634
rect 50306 41582 50318 41634
rect 50370 41582 50382 41634
rect 14366 41570 14418 41582
rect 41346 41470 41358 41522
rect 41410 41470 41422 41522
rect 45042 41470 45054 41522
rect 45106 41470 45118 41522
rect 1344 41354 58576 41388
rect 1344 41302 4478 41354
rect 4530 41302 4582 41354
rect 4634 41302 4686 41354
rect 4738 41302 35198 41354
rect 35250 41302 35302 41354
rect 35354 41302 35406 41354
rect 35458 41302 58576 41354
rect 1344 41268 58576 41302
rect 5618 41134 5630 41186
rect 5682 41134 5694 41186
rect 17042 41134 17054 41186
rect 17106 41183 17118 41186
rect 17602 41183 17614 41186
rect 17106 41137 17614 41183
rect 17106 41134 17118 41137
rect 17602 41134 17614 41137
rect 17666 41134 17678 41186
rect 53330 41134 53342 41186
rect 53394 41134 53406 41186
rect 42590 41074 42642 41086
rect 21298 41022 21310 41074
rect 21362 41071 21374 41074
rect 22306 41071 22318 41074
rect 21362 41025 22318 41071
rect 21362 41022 21374 41025
rect 22306 41022 22318 41025
rect 22370 41022 22382 41074
rect 42590 41010 42642 41022
rect 6078 40962 6130 40974
rect 6078 40898 6130 40910
rect 17166 40962 17218 40974
rect 17166 40898 17218 40910
rect 17614 40962 17666 40974
rect 17614 40898 17666 40910
rect 23550 40962 23602 40974
rect 23550 40898 23602 40910
rect 31614 40962 31666 40974
rect 31614 40898 31666 40910
rect 34414 40962 34466 40974
rect 34414 40898 34466 40910
rect 34750 40962 34802 40974
rect 35858 40910 35870 40962
rect 35922 40910 35934 40962
rect 34750 40898 34802 40910
rect 1822 40850 1874 40862
rect 9662 40850 9714 40862
rect 17950 40850 18002 40862
rect 2370 40798 2382 40850
rect 2434 40798 2446 40850
rect 5730 40798 5742 40850
rect 5794 40798 5806 40850
rect 10210 40798 10222 40850
rect 10274 40798 10286 40850
rect 1822 40786 1874 40798
rect 9662 40786 9714 40798
rect 17950 40786 18002 40798
rect 20750 40850 20802 40862
rect 20750 40786 20802 40798
rect 24222 40850 24274 40862
rect 24222 40786 24274 40798
rect 26014 40850 26066 40862
rect 30494 40850 30546 40862
rect 27458 40798 27470 40850
rect 27522 40798 27534 40850
rect 26014 40786 26066 40798
rect 30494 40786 30546 40798
rect 30718 40850 30770 40862
rect 30718 40786 30770 40798
rect 37326 40850 37378 40862
rect 37326 40786 37378 40798
rect 37886 40850 37938 40862
rect 37886 40786 37938 40798
rect 38670 40850 38722 40862
rect 38670 40786 38722 40798
rect 41582 40850 41634 40862
rect 41582 40786 41634 40798
rect 42926 40850 42978 40862
rect 42926 40786 42978 40798
rect 44046 40850 44098 40862
rect 46174 40850 46226 40862
rect 54462 40850 54514 40862
rect 45378 40798 45390 40850
rect 45442 40798 45454 40850
rect 46722 40798 46734 40850
rect 46786 40798 46798 40850
rect 47506 40798 47518 40850
rect 47570 40798 47582 40850
rect 53218 40798 53230 40850
rect 53282 40798 53294 40850
rect 44046 40786 44098 40798
rect 46174 40786 46226 40798
rect 54462 40786 54514 40798
rect 13470 40738 13522 40750
rect 13470 40674 13522 40686
rect 23886 40738 23938 40750
rect 23886 40674 23938 40686
rect 29822 40738 29874 40750
rect 29822 40674 29874 40686
rect 31166 40738 31218 40750
rect 31166 40674 31218 40686
rect 37662 40738 37714 40750
rect 37662 40674 37714 40686
rect 41246 40738 41298 40750
rect 56142 40738 56194 40750
rect 43026 40686 43038 40738
rect 43090 40735 43102 40738
rect 43090 40689 43199 40735
rect 43090 40686 43102 40689
rect 41246 40674 41298 40686
rect 4510 40626 4562 40638
rect 4510 40562 4562 40574
rect 4958 40626 5010 40638
rect 4958 40562 5010 40574
rect 6190 40626 6242 40638
rect 6190 40562 6242 40574
rect 9326 40626 9378 40638
rect 9326 40562 9378 40574
rect 12350 40626 12402 40638
rect 12350 40562 12402 40574
rect 12798 40626 12850 40638
rect 12798 40562 12850 40574
rect 13582 40626 13634 40638
rect 13582 40562 13634 40574
rect 18734 40626 18786 40638
rect 18734 40562 18786 40574
rect 21422 40626 21474 40638
rect 21422 40562 21474 40574
rect 21870 40626 21922 40638
rect 21870 40562 21922 40574
rect 22318 40626 22370 40638
rect 22318 40562 22370 40574
rect 23102 40626 23154 40638
rect 23102 40562 23154 40574
rect 27582 40626 27634 40638
rect 27582 40562 27634 40574
rect 29374 40626 29426 40638
rect 29374 40562 29426 40574
rect 30270 40626 30322 40638
rect 30270 40562 30322 40574
rect 37102 40626 37154 40638
rect 37102 40562 37154 40574
rect 42366 40626 42418 40638
rect 42366 40562 42418 40574
rect 21858 40462 21870 40514
rect 21922 40511 21934 40514
rect 22418 40511 22430 40514
rect 21922 40465 22430 40511
rect 21922 40462 21934 40465
rect 22418 40462 22430 40465
rect 22482 40462 22494 40514
rect 27010 40462 27022 40514
rect 27074 40462 27086 40514
rect 43153 40511 43199 40689
rect 54562 40686 54574 40738
rect 54626 40686 54638 40738
rect 56142 40674 56194 40686
rect 43486 40626 43538 40638
rect 44930 40574 44942 40626
rect 44994 40574 45006 40626
rect 43486 40562 43538 40574
rect 43474 40511 43486 40514
rect 43153 40465 43486 40511
rect 43474 40462 43486 40465
rect 43538 40462 43550 40514
rect 49410 40462 49422 40514
rect 49474 40462 49486 40514
rect 1344 40346 58576 40380
rect 1344 40294 19838 40346
rect 19890 40294 19942 40346
rect 19994 40294 20046 40346
rect 20098 40294 50558 40346
rect 50610 40294 50662 40346
rect 50714 40294 50766 40346
rect 50818 40294 58576 40346
rect 1344 40260 58576 40294
rect 17378 40126 17390 40178
rect 17442 40126 17454 40178
rect 21970 40126 21982 40178
rect 22034 40126 22046 40178
rect 37538 40126 37550 40178
rect 37602 40126 37614 40178
rect 1822 40066 1874 40078
rect 1822 40002 1874 40014
rect 6862 40066 6914 40078
rect 6862 40002 6914 40014
rect 13470 40066 13522 40078
rect 13470 40002 13522 40014
rect 24222 40066 24274 40078
rect 24222 40002 24274 40014
rect 24670 40066 24722 40078
rect 24670 40002 24722 40014
rect 32286 40066 32338 40078
rect 32286 40002 32338 40014
rect 34078 40066 34130 40078
rect 43710 40066 43762 40078
rect 39890 40014 39902 40066
rect 39954 40014 39966 40066
rect 34078 40002 34130 40014
rect 43710 40002 43762 40014
rect 47854 40066 47906 40078
rect 47854 40002 47906 40014
rect 52334 40066 52386 40078
rect 52334 40002 52386 40014
rect 53118 40066 53170 40078
rect 54898 40014 54910 40066
rect 54962 40014 54974 40066
rect 53118 40002 53170 40014
rect 16830 39954 16882 39966
rect 16830 39890 16882 39902
rect 17838 39954 17890 39966
rect 17838 39890 17890 39902
rect 18398 39954 18450 39966
rect 18398 39890 18450 39902
rect 19742 39954 19794 39966
rect 19742 39890 19794 39902
rect 22430 39954 22482 39966
rect 22430 39890 22482 39902
rect 22878 39954 22930 39966
rect 22878 39890 22930 39902
rect 25118 39954 25170 39966
rect 25118 39890 25170 39902
rect 25454 39954 25506 39966
rect 25454 39890 25506 39902
rect 27134 39954 27186 39966
rect 27134 39890 27186 39902
rect 29262 39954 29314 39966
rect 29262 39890 29314 39902
rect 29822 39954 29874 39966
rect 29822 39890 29874 39902
rect 30382 39954 30434 39966
rect 30382 39890 30434 39902
rect 33070 39954 33122 39966
rect 33070 39890 33122 39902
rect 34974 39954 35026 39966
rect 34974 39890 35026 39902
rect 35534 39954 35586 39966
rect 35534 39890 35586 39902
rect 38334 39954 38386 39966
rect 38334 39890 38386 39902
rect 40910 39954 40962 39966
rect 40910 39890 40962 39902
rect 41582 39954 41634 39966
rect 41582 39890 41634 39902
rect 42478 39954 42530 39966
rect 42478 39890 42530 39902
rect 43038 39954 43090 39966
rect 43038 39890 43090 39902
rect 45054 39954 45106 39966
rect 45054 39890 45106 39902
rect 45726 39954 45778 39966
rect 47182 39954 47234 39966
rect 46498 39902 46510 39954
rect 46562 39902 46574 39954
rect 45726 39890 45778 39902
rect 47182 39890 47234 39902
rect 49198 39954 49250 39966
rect 49198 39890 49250 39902
rect 49534 39954 49586 39966
rect 49534 39890 49586 39902
rect 49870 39954 49922 39966
rect 49870 39890 49922 39902
rect 50206 39954 50258 39966
rect 50206 39890 50258 39902
rect 51102 39954 51154 39966
rect 51102 39890 51154 39902
rect 51662 39954 51714 39966
rect 51662 39890 51714 39902
rect 53230 39954 53282 39966
rect 54562 39902 54574 39954
rect 54626 39902 54638 39954
rect 55570 39902 55582 39954
rect 55634 39902 55646 39954
rect 53230 39890 53282 39902
rect 4174 39842 4226 39854
rect 10782 39842 10834 39854
rect 18958 39842 19010 39854
rect 36430 39842 36482 39854
rect 4722 39790 4734 39842
rect 4786 39790 4798 39842
rect 11330 39790 11342 39842
rect 11394 39790 11406 39842
rect 22642 39790 22654 39842
rect 22706 39790 22718 39842
rect 28466 39790 28478 39842
rect 28530 39790 28542 39842
rect 4174 39778 4226 39790
rect 10782 39778 10834 39790
rect 18958 39778 19010 39790
rect 36430 39778 36482 39790
rect 37886 39842 37938 39854
rect 37886 39778 37938 39790
rect 41246 39842 41298 39854
rect 41246 39778 41298 39790
rect 41918 39842 41970 39854
rect 41918 39778 41970 39790
rect 44494 39842 44546 39854
rect 44494 39778 44546 39790
rect 45390 39842 45442 39854
rect 45390 39778 45442 39790
rect 46062 39842 46114 39854
rect 46062 39778 46114 39790
rect 50542 39842 50594 39854
rect 50542 39778 50594 39790
rect 53006 39842 53058 39854
rect 53006 39778 53058 39790
rect 53454 39848 53506 39860
rect 53454 39784 53506 39796
rect 54014 39842 54066 39854
rect 54338 39790 54350 39842
rect 54402 39790 54414 39842
rect 55346 39790 55358 39842
rect 55410 39790 55422 39842
rect 54014 39778 54066 39790
rect 3838 39730 3890 39742
rect 3838 39666 3890 39678
rect 10446 39730 10498 39742
rect 10446 39666 10498 39678
rect 16494 39730 16546 39742
rect 16494 39666 16546 39678
rect 18510 39730 18562 39742
rect 18510 39666 18562 39678
rect 29934 39730 29986 39742
rect 29934 39666 29986 39678
rect 35646 39730 35698 39742
rect 35646 39666 35698 39678
rect 36990 39730 37042 39742
rect 36990 39666 37042 39678
rect 56702 39730 56754 39742
rect 56702 39666 56754 39678
rect 57150 39730 57202 39742
rect 57150 39666 57202 39678
rect 28366 39618 28418 39630
rect 7298 39566 7310 39618
rect 7362 39566 7374 39618
rect 13906 39566 13918 39618
rect 13970 39566 13982 39618
rect 21746 39566 21758 39618
rect 21810 39566 21822 39618
rect 27906 39566 27918 39618
rect 27970 39566 27982 39618
rect 28366 39554 28418 39566
rect 36094 39618 36146 39630
rect 36094 39554 36146 39566
rect 28802 39454 28814 39506
rect 28866 39454 28878 39506
rect 34514 39454 34526 39506
rect 34578 39454 34590 39506
rect 1344 39338 58576 39372
rect 1344 39286 4478 39338
rect 4530 39286 4582 39338
rect 4634 39286 4686 39338
rect 4738 39286 35198 39338
rect 35250 39286 35302 39338
rect 35354 39286 35406 39338
rect 35458 39286 58576 39338
rect 1344 39252 58576 39286
rect 4946 39118 4958 39170
rect 5010 39118 5022 39170
rect 12674 39118 12686 39170
rect 12738 39118 12750 39170
rect 18050 39118 18062 39170
rect 18114 39118 18126 39170
rect 19506 39118 19518 39170
rect 19570 39118 19582 39170
rect 37202 39118 37214 39170
rect 37266 39167 37278 39170
rect 38322 39167 38334 39170
rect 37266 39121 38334 39167
rect 37266 39118 37278 39121
rect 38322 39118 38334 39121
rect 38386 39118 38398 39170
rect 21646 39058 21698 39070
rect 39230 39058 39282 39070
rect 25442 39006 25454 39058
rect 25506 39006 25518 39058
rect 36978 39006 36990 39058
rect 37042 39055 37054 39058
rect 37762 39055 37774 39058
rect 37042 39009 37774 39055
rect 37042 39006 37054 39009
rect 37762 39006 37774 39009
rect 37826 39006 37838 39058
rect 21646 38994 21698 39006
rect 39230 38994 39282 39006
rect 17390 38946 17442 38958
rect 17390 38882 17442 38894
rect 28030 38946 28082 38958
rect 28030 38882 28082 38894
rect 29374 38946 29426 38958
rect 29374 38882 29426 38894
rect 30046 38946 30098 38958
rect 30046 38882 30098 38894
rect 32510 38946 32562 38958
rect 32510 38882 32562 38894
rect 34414 38946 34466 38958
rect 34414 38882 34466 38894
rect 37214 38946 37266 38958
rect 37214 38882 37266 38894
rect 37662 38946 37714 38958
rect 37662 38882 37714 38894
rect 38110 38946 38162 38958
rect 38110 38882 38162 38894
rect 38558 38946 38610 38958
rect 38558 38882 38610 38894
rect 43038 38946 43090 38958
rect 43038 38882 43090 38894
rect 50878 38946 50930 38958
rect 50878 38882 50930 38894
rect 51774 38946 51826 38958
rect 51774 38882 51826 38894
rect 52782 38946 52834 38958
rect 52782 38882 52834 38894
rect 54686 38946 54738 38958
rect 54686 38882 54738 38894
rect 8878 38834 8930 38846
rect 19966 38834 20018 38846
rect 8306 38782 8318 38834
rect 8370 38782 8382 38834
rect 12786 38782 12798 38834
rect 12850 38782 12862 38834
rect 18722 38782 18734 38834
rect 18786 38782 18798 38834
rect 8878 38770 8930 38782
rect 19966 38770 20018 38782
rect 22654 38834 22706 38846
rect 22654 38770 22706 38782
rect 26574 38834 26626 38846
rect 26574 38770 26626 38782
rect 27582 38834 27634 38846
rect 27582 38770 27634 38782
rect 28478 38834 28530 38846
rect 42254 38834 42306 38846
rect 33618 38782 33630 38834
rect 33682 38782 33694 38834
rect 28478 38770 28530 38782
rect 42254 38770 42306 38782
rect 46734 38834 46786 38846
rect 46734 38770 46786 38782
rect 55358 38834 55410 38846
rect 55358 38770 55410 38782
rect 56478 38834 56530 38846
rect 56478 38770 56530 38782
rect 4622 38722 4674 38734
rect 4622 38658 4674 38670
rect 5070 38722 5122 38734
rect 5070 38658 5122 38670
rect 5742 38722 5794 38734
rect 5742 38658 5794 38670
rect 13470 38722 13522 38734
rect 13470 38658 13522 38670
rect 16606 38722 16658 38734
rect 16606 38658 16658 38670
rect 17838 38722 17890 38734
rect 17838 38658 17890 38670
rect 18510 38722 18562 38734
rect 18510 38658 18562 38670
rect 18958 38722 19010 38734
rect 18958 38658 19010 38670
rect 20414 38722 20466 38734
rect 20414 38658 20466 38670
rect 20638 38722 20690 38734
rect 20638 38658 20690 38670
rect 21310 38722 21362 38734
rect 21310 38658 21362 38670
rect 27134 38722 27186 38734
rect 27134 38658 27186 38670
rect 27246 38722 27298 38734
rect 27246 38658 27298 38670
rect 33182 38722 33234 38734
rect 33182 38658 33234 38670
rect 33742 38722 33794 38734
rect 33742 38658 33794 38670
rect 38894 38722 38946 38734
rect 38894 38658 38946 38670
rect 40462 38722 40514 38734
rect 42702 38722 42754 38734
rect 41122 38670 41134 38722
rect 41186 38670 41198 38722
rect 40462 38658 40514 38670
rect 42702 38658 42754 38670
rect 47182 38722 47234 38734
rect 47182 38658 47234 38670
rect 47406 38722 47458 38734
rect 47406 38658 47458 38670
rect 13582 38610 13634 38622
rect 6066 38558 6078 38610
rect 6130 38558 6142 38610
rect 13582 38546 13634 38558
rect 17054 38610 17106 38622
rect 17054 38546 17106 38558
rect 22206 38610 22258 38622
rect 22206 38546 22258 38558
rect 23438 38610 23490 38622
rect 23438 38546 23490 38558
rect 27806 38610 27858 38622
rect 39790 38610 39842 38622
rect 28242 38558 28254 38610
rect 28306 38558 28318 38610
rect 27806 38546 27858 38558
rect 39790 38546 39842 38558
rect 41918 38610 41970 38622
rect 41918 38546 41970 38558
rect 44942 38610 44994 38622
rect 44942 38546 44994 38558
rect 49982 38610 50034 38622
rect 49982 38546 50034 38558
rect 50430 38610 50482 38622
rect 50430 38546 50482 38558
rect 51326 38610 51378 38622
rect 51326 38546 51378 38558
rect 53230 38610 53282 38622
rect 53230 38546 53282 38558
rect 53678 38610 53730 38622
rect 53678 38546 53730 38558
rect 57038 38610 57090 38622
rect 57038 38546 57090 38558
rect 26114 38446 26126 38498
rect 26178 38446 26190 38498
rect 32722 38446 32734 38498
rect 32786 38446 32798 38498
rect 46274 38446 46286 38498
rect 46338 38446 46350 38498
rect 49970 38446 49982 38498
rect 50034 38495 50046 38498
rect 51314 38495 51326 38498
rect 50034 38449 51326 38495
rect 50034 38446 50046 38449
rect 51314 38446 51326 38449
rect 51378 38446 51390 38498
rect 52546 38446 52558 38498
rect 52610 38495 52622 38498
rect 53218 38495 53230 38498
rect 52610 38449 53230 38495
rect 52610 38446 52622 38449
rect 53218 38446 53230 38449
rect 53282 38495 53294 38498
rect 53666 38495 53678 38498
rect 53282 38449 53678 38495
rect 53282 38446 53294 38449
rect 53666 38446 53678 38449
rect 53730 38446 53742 38498
rect 1344 38330 58576 38364
rect 1344 38278 19838 38330
rect 19890 38278 19942 38330
rect 19994 38278 20046 38330
rect 20098 38278 50558 38330
rect 50610 38278 50662 38330
rect 50714 38278 50766 38330
rect 50818 38278 58576 38330
rect 1344 38244 58576 38278
rect 7074 38110 7086 38162
rect 7138 38110 7150 38162
rect 7522 38110 7534 38162
rect 7586 38110 7598 38162
rect 18834 38110 18846 38162
rect 18898 38159 18910 38162
rect 19394 38159 19406 38162
rect 18898 38113 19406 38159
rect 18898 38110 18910 38113
rect 19394 38110 19406 38113
rect 19458 38110 19470 38162
rect 27458 38110 27470 38162
rect 27522 38110 27534 38162
rect 33730 38110 33742 38162
rect 33794 38110 33806 38162
rect 36306 38110 36318 38162
rect 36370 38110 36382 38162
rect 39218 38110 39230 38162
rect 39282 38159 39294 38162
rect 39778 38159 39790 38162
rect 39282 38113 39790 38159
rect 39282 38110 39294 38113
rect 39778 38110 39790 38113
rect 39842 38110 39854 38162
rect 49298 38110 49310 38162
rect 49362 38159 49374 38162
rect 49634 38159 49646 38162
rect 49362 38113 49646 38159
rect 49362 38110 49374 38113
rect 49634 38110 49646 38113
rect 49698 38159 49710 38162
rect 50642 38159 50654 38162
rect 49698 38113 50654 38159
rect 49698 38110 49710 38113
rect 50642 38110 50654 38113
rect 50706 38159 50718 38162
rect 51650 38159 51662 38162
rect 50706 38113 51662 38159
rect 50706 38110 50718 38113
rect 51650 38110 51662 38113
rect 51714 38110 51726 38162
rect 6190 38050 6242 38062
rect 6190 37986 6242 37998
rect 7198 38050 7250 38062
rect 7198 37986 7250 37998
rect 14366 38050 14418 38062
rect 14366 37986 14418 37998
rect 17502 38050 17554 38062
rect 17502 37986 17554 37998
rect 17950 38050 18002 38062
rect 17950 37986 18002 37998
rect 19518 38050 19570 38062
rect 19518 37986 19570 37998
rect 25454 38050 25506 38062
rect 25454 37986 25506 37998
rect 28142 38050 28194 38062
rect 28142 37986 28194 37998
rect 28590 38050 28642 38062
rect 28590 37986 28642 37998
rect 38782 38050 38834 38062
rect 38782 37986 38834 37998
rect 41918 38050 41970 38062
rect 41918 37986 41970 37998
rect 48190 38050 48242 38062
rect 48190 37986 48242 37998
rect 49310 38050 49362 38062
rect 49310 37986 49362 37998
rect 50206 38050 50258 38062
rect 50206 37986 50258 37998
rect 50654 38050 50706 38062
rect 50654 37986 50706 37998
rect 56030 38050 56082 38062
rect 56030 37986 56082 37998
rect 20414 37938 20466 37950
rect 20414 37874 20466 37886
rect 21534 37938 21586 37950
rect 21534 37874 21586 37886
rect 21758 37938 21810 37950
rect 21758 37874 21810 37886
rect 22094 37938 22146 37950
rect 22094 37874 22146 37886
rect 23550 37938 23602 37950
rect 26462 37938 26514 37950
rect 25778 37886 25790 37938
rect 25842 37886 25854 37938
rect 23550 37874 23602 37886
rect 26462 37874 26514 37886
rect 27022 37938 27074 37950
rect 27022 37874 27074 37886
rect 41246 37938 41298 37950
rect 41246 37874 41298 37886
rect 41582 37938 41634 37950
rect 41582 37874 41634 37886
rect 43710 37938 43762 37950
rect 43710 37874 43762 37886
rect 46846 37938 46898 37950
rect 46846 37874 46898 37886
rect 47294 37938 47346 37950
rect 47294 37874 47346 37886
rect 52558 37938 52610 37950
rect 52558 37874 52610 37886
rect 3502 37826 3554 37838
rect 11678 37826 11730 37838
rect 18398 37826 18450 37838
rect 4050 37774 4062 37826
rect 4114 37774 4126 37826
rect 7634 37774 7646 37826
rect 7698 37774 7710 37826
rect 12226 37774 12238 37826
rect 12290 37774 12302 37826
rect 3502 37762 3554 37774
rect 11678 37762 11730 37774
rect 18398 37762 18450 37774
rect 19406 37826 19458 37838
rect 19406 37762 19458 37774
rect 19966 37826 20018 37838
rect 21086 37826 21138 37838
rect 20290 37774 20302 37826
rect 20354 37774 20366 37826
rect 19966 37762 20018 37774
rect 21086 37762 21138 37774
rect 21310 37826 21362 37838
rect 25118 37826 25170 37838
rect 22642 37774 22654 37826
rect 22706 37774 22718 37826
rect 21310 37762 21362 37774
rect 25118 37762 25170 37774
rect 26014 37826 26066 37838
rect 36654 37826 36706 37838
rect 35298 37774 35310 37826
rect 35362 37774 35374 37826
rect 26014 37762 26066 37774
rect 36654 37762 36706 37774
rect 40910 37826 40962 37838
rect 40910 37762 40962 37774
rect 42478 37826 42530 37838
rect 42478 37762 42530 37774
rect 43038 37826 43090 37838
rect 43038 37762 43090 37774
rect 45278 37826 45330 37838
rect 45278 37762 45330 37774
rect 51550 37826 51602 37838
rect 53790 37826 53842 37838
rect 52714 37774 52726 37826
rect 52778 37774 52790 37826
rect 51550 37762 51602 37774
rect 53790 37762 53842 37774
rect 3166 37714 3218 37726
rect 3166 37650 3218 37662
rect 11342 37714 11394 37726
rect 11342 37650 11394 37662
rect 16830 37714 16882 37726
rect 16830 37650 16882 37662
rect 18846 37714 18898 37726
rect 18846 37650 18898 37662
rect 23214 37714 23266 37726
rect 23214 37650 23266 37662
rect 25566 37714 25618 37726
rect 25566 37650 25618 37662
rect 26350 37714 26402 37726
rect 26350 37650 26402 37662
rect 32510 37714 32562 37726
rect 32510 37650 32562 37662
rect 39230 37714 39282 37726
rect 39230 37650 39282 37662
rect 39678 37714 39730 37726
rect 39678 37650 39730 37662
rect 40350 37714 40402 37726
rect 40350 37650 40402 37662
rect 44942 37714 44994 37726
rect 44942 37650 44994 37662
rect 47518 37714 47570 37726
rect 47518 37650 47570 37662
rect 48862 37714 48914 37726
rect 48862 37650 48914 37662
rect 49758 37714 49810 37726
rect 49758 37650 49810 37662
rect 51102 37714 51154 37726
rect 51102 37650 51154 37662
rect 55582 37714 55634 37726
rect 55582 37650 55634 37662
rect 56702 37714 56754 37726
rect 56702 37650 56754 37662
rect 57150 37714 57202 37726
rect 57150 37650 57202 37662
rect 57598 37714 57650 37726
rect 57598 37650 57650 37662
rect 6626 37550 6638 37602
rect 6690 37550 6702 37602
rect 14802 37550 14814 37602
rect 14866 37550 14878 37602
rect 51090 37550 51102 37602
rect 51154 37599 51166 37602
rect 51314 37599 51326 37602
rect 51154 37553 51326 37599
rect 51154 37550 51166 37553
rect 51314 37550 51326 37553
rect 51378 37550 51390 37602
rect 21186 37438 21198 37490
rect 21250 37438 21262 37490
rect 22194 37438 22206 37490
rect 22258 37438 22270 37490
rect 22530 37438 22542 37490
rect 22594 37438 22606 37490
rect 46386 37438 46398 37490
rect 46450 37438 46462 37490
rect 49746 37438 49758 37490
rect 49810 37487 49822 37490
rect 50194 37487 50206 37490
rect 49810 37441 50206 37487
rect 49810 37438 49822 37441
rect 50194 37438 50206 37441
rect 50258 37438 50270 37490
rect 54338 37438 54350 37490
rect 54402 37438 54414 37490
rect 1344 37322 58576 37356
rect 1344 37270 4478 37322
rect 4530 37270 4582 37322
rect 4634 37270 4686 37322
rect 4738 37270 35198 37322
rect 35250 37270 35302 37322
rect 35354 37270 35406 37322
rect 35458 37270 58576 37322
rect 1344 37236 58576 37270
rect 4386 37102 4398 37154
rect 4450 37102 4462 37154
rect 23090 37102 23102 37154
rect 23154 37102 23166 37154
rect 33058 37102 33070 37154
rect 33122 37102 33134 37154
rect 43810 37102 43822 37154
rect 43874 37102 43886 37154
rect 8766 36930 8818 36942
rect 8766 36866 8818 36878
rect 14702 36930 14754 36942
rect 14702 36866 14754 36878
rect 19182 36930 19234 36942
rect 19182 36866 19234 36878
rect 20750 36930 20802 36942
rect 20750 36866 20802 36878
rect 24782 36930 24834 36942
rect 24782 36866 24834 36878
rect 37326 36930 37378 36942
rect 37326 36866 37378 36878
rect 37998 36930 38050 36942
rect 50418 36878 50430 36930
rect 50482 36878 50494 36930
rect 51538 36927 51550 36930
rect 50881 36881 51550 36927
rect 37998 36866 38050 36878
rect 5630 36818 5682 36830
rect 15038 36818 15090 36830
rect 4498 36766 4510 36818
rect 4562 36766 4574 36818
rect 6178 36766 6190 36818
rect 6242 36766 6254 36818
rect 5630 36754 5682 36766
rect 15038 36754 15090 36766
rect 17838 36818 17890 36830
rect 17838 36754 17890 36766
rect 20414 36818 20466 36830
rect 20414 36754 20466 36766
rect 21310 36818 21362 36830
rect 21310 36754 21362 36766
rect 23550 36818 23602 36830
rect 23550 36754 23602 36766
rect 30718 36818 30770 36830
rect 42926 36818 42978 36830
rect 32498 36766 32510 36818
rect 32562 36766 32574 36818
rect 30718 36754 30770 36766
rect 42926 36754 42978 36766
rect 43038 36818 43090 36830
rect 43038 36754 43090 36766
rect 43934 36818 43986 36830
rect 43934 36754 43986 36766
rect 44046 36818 44098 36830
rect 44046 36754 44098 36766
rect 46174 36818 46226 36830
rect 49870 36818 49922 36830
rect 49634 36766 49646 36818
rect 49698 36766 49710 36818
rect 46174 36754 46226 36766
rect 49870 36754 49922 36766
rect 50094 36818 50146 36830
rect 50094 36754 50146 36766
rect 50318 36818 50370 36830
rect 50642 36766 50654 36818
rect 50706 36815 50718 36818
rect 50881 36815 50927 36881
rect 51538 36878 51550 36881
rect 51602 36878 51614 36930
rect 53678 36818 53730 36830
rect 50706 36769 50927 36815
rect 50706 36766 50718 36769
rect 51426 36766 51438 36818
rect 51490 36766 51502 36818
rect 50318 36754 50370 36766
rect 53678 36754 53730 36766
rect 56926 36818 56978 36830
rect 56926 36754 56978 36766
rect 57486 36818 57538 36830
rect 57486 36754 57538 36766
rect 18510 36706 18562 36718
rect 18510 36642 18562 36654
rect 19070 36706 19122 36718
rect 19070 36642 19122 36654
rect 20078 36706 20130 36718
rect 20078 36642 20130 36654
rect 21982 36706 22034 36718
rect 21982 36642 22034 36654
rect 22206 36706 22258 36718
rect 22206 36642 22258 36654
rect 22430 36706 22482 36718
rect 22430 36642 22482 36654
rect 22654 36706 22706 36718
rect 22654 36642 22706 36654
rect 23998 36706 24050 36718
rect 23998 36642 24050 36654
rect 24222 36706 24274 36718
rect 24222 36642 24274 36654
rect 29262 36706 29314 36718
rect 29262 36642 29314 36654
rect 29374 36706 29426 36718
rect 29374 36642 29426 36654
rect 29934 36706 29986 36718
rect 29934 36642 29986 36654
rect 37662 36706 37714 36718
rect 37662 36642 37714 36654
rect 38334 36706 38386 36718
rect 38334 36642 38386 36654
rect 38670 36706 38722 36718
rect 38670 36642 38722 36654
rect 39006 36706 39058 36718
rect 39006 36642 39058 36654
rect 39902 36706 39954 36718
rect 39902 36642 39954 36654
rect 40462 36706 40514 36718
rect 40462 36642 40514 36654
rect 45502 36706 45554 36718
rect 45502 36642 45554 36654
rect 46062 36706 46114 36718
rect 46062 36642 46114 36654
rect 46734 36706 46786 36718
rect 46734 36642 46786 36654
rect 47070 36706 47122 36718
rect 47070 36642 47122 36654
rect 47742 36706 47794 36718
rect 47742 36642 47794 36654
rect 50542 36706 50594 36718
rect 50542 36642 50594 36654
rect 50878 36706 50930 36718
rect 50878 36642 50930 36654
rect 51214 36706 51266 36718
rect 51214 36642 51266 36654
rect 52110 36706 52162 36718
rect 52110 36642 52162 36654
rect 53006 36706 53058 36718
rect 53006 36642 53058 36654
rect 53342 36706 53394 36718
rect 55134 36706 55186 36718
rect 54450 36654 54462 36706
rect 54514 36654 54526 36706
rect 53342 36642 53394 36654
rect 55134 36642 55186 36654
rect 57150 36706 57202 36718
rect 57150 36642 57202 36654
rect 57934 36706 57986 36718
rect 57934 36642 57986 36654
rect 4062 36594 4114 36606
rect 4062 36530 4114 36542
rect 4958 36594 5010 36606
rect 4958 36530 5010 36542
rect 8318 36594 8370 36606
rect 8318 36530 8370 36542
rect 11006 36594 11058 36606
rect 11006 36530 11058 36542
rect 13582 36594 13634 36606
rect 13582 36530 13634 36542
rect 15822 36594 15874 36606
rect 15822 36530 15874 36542
rect 18062 36594 18114 36606
rect 18062 36530 18114 36542
rect 21646 36594 21698 36606
rect 21646 36530 21698 36542
rect 28590 36594 28642 36606
rect 28590 36530 28642 36542
rect 32174 36594 32226 36606
rect 32174 36530 32226 36542
rect 35982 36594 36034 36606
rect 35982 36530 36034 36542
rect 36430 36594 36482 36606
rect 36430 36530 36482 36542
rect 39342 36594 39394 36606
rect 39342 36530 39394 36542
rect 41134 36594 41186 36606
rect 41134 36530 41186 36542
rect 41918 36594 41970 36606
rect 41918 36530 41970 36542
rect 51662 36594 51714 36606
rect 51662 36530 51714 36542
rect 54014 36594 54066 36606
rect 54014 36530 54066 36542
rect 55806 36594 55858 36606
rect 55806 36530 55858 36542
rect 56590 36594 56642 36606
rect 56590 36530 56642 36542
rect 4834 36430 4846 36482
rect 4898 36430 4910 36482
rect 13458 36430 13470 36482
rect 13522 36430 13534 36482
rect 22754 36430 22766 36482
rect 22818 36430 22830 36482
rect 30370 36430 30382 36482
rect 30434 36430 30446 36482
rect 45042 36430 45054 36482
rect 45106 36430 45118 36482
rect 48850 36430 48862 36482
rect 48914 36430 48926 36482
rect 1344 36314 58576 36348
rect 1344 36262 19838 36314
rect 19890 36262 19942 36314
rect 19994 36262 20046 36314
rect 20098 36262 50558 36314
rect 50610 36262 50662 36314
rect 50714 36262 50766 36314
rect 50818 36262 58576 36314
rect 1344 36228 58576 36262
rect 3714 36094 3726 36146
rect 3778 36143 3790 36146
rect 4498 36143 4510 36146
rect 3778 36097 4510 36143
rect 3778 36094 3790 36097
rect 4498 36094 4510 36097
rect 4562 36094 4574 36146
rect 37986 36094 37998 36146
rect 38050 36094 38062 36146
rect 39778 36094 39790 36146
rect 39842 36094 39854 36146
rect 2718 36034 2770 36046
rect 6190 36034 6242 36046
rect 5842 35982 5854 36034
rect 5906 35982 5918 36034
rect 2718 35970 2770 35982
rect 6190 35970 6242 35982
rect 21310 36034 21362 36046
rect 21310 35970 21362 35982
rect 21758 36034 21810 36046
rect 21758 35970 21810 35982
rect 21982 36034 22034 36046
rect 21982 35970 22034 35982
rect 24782 36034 24834 36046
rect 30158 36034 30210 36046
rect 25330 35982 25342 36034
rect 25394 35982 25406 36034
rect 24782 35970 24834 35982
rect 30158 35970 30210 35982
rect 36318 36034 36370 36046
rect 36318 35970 36370 35982
rect 40798 36034 40850 36046
rect 40798 35970 40850 35982
rect 44382 36034 44434 36046
rect 44382 35970 44434 35982
rect 44830 36034 44882 36046
rect 44830 35970 44882 35982
rect 45614 36034 45666 36046
rect 45614 35970 45666 35982
rect 46734 36034 46786 36046
rect 46734 35970 46786 35982
rect 48302 36034 48354 36046
rect 48302 35970 48354 35982
rect 51550 36034 51602 36046
rect 51550 35970 51602 35982
rect 52334 36034 52386 36046
rect 52334 35970 52386 35982
rect 56702 36034 56754 36046
rect 56702 35970 56754 35982
rect 12126 35922 12178 35934
rect 12126 35858 12178 35870
rect 14478 35922 14530 35934
rect 14478 35858 14530 35870
rect 18958 35922 19010 35934
rect 18958 35858 19010 35870
rect 19070 35922 19122 35934
rect 19070 35858 19122 35870
rect 19742 35922 19794 35934
rect 19742 35858 19794 35870
rect 22878 35922 22930 35934
rect 22878 35858 22930 35870
rect 23774 35922 23826 35934
rect 23774 35858 23826 35870
rect 25566 35922 25618 35934
rect 25566 35858 25618 35870
rect 25790 35922 25842 35934
rect 25790 35858 25842 35870
rect 27022 35922 27074 35934
rect 27022 35858 27074 35870
rect 43150 35922 43202 35934
rect 43150 35858 43202 35870
rect 49086 35922 49138 35934
rect 49086 35858 49138 35870
rect 49422 35922 49474 35934
rect 49422 35858 49474 35870
rect 50318 35922 50370 35934
rect 50318 35858 50370 35870
rect 54238 35922 54290 35934
rect 54238 35858 54290 35870
rect 3054 35810 3106 35822
rect 10782 35810 10834 35822
rect 3602 35758 3614 35810
rect 3666 35758 3678 35810
rect 3054 35746 3106 35758
rect 10782 35746 10834 35758
rect 11342 35810 11394 35822
rect 18398 35810 18450 35822
rect 14578 35758 14590 35810
rect 14642 35758 14654 35810
rect 11342 35746 11394 35758
rect 18398 35746 18450 35758
rect 19518 35810 19570 35822
rect 19518 35746 19570 35758
rect 19630 35810 19682 35822
rect 19630 35746 19682 35758
rect 19966 35810 20018 35822
rect 24334 35810 24386 35822
rect 24098 35758 24110 35810
rect 24162 35758 24174 35810
rect 19966 35746 20018 35758
rect 24334 35746 24386 35758
rect 25118 35810 25170 35822
rect 25118 35746 25170 35758
rect 25902 35810 25954 35822
rect 25902 35746 25954 35758
rect 26238 35810 26290 35822
rect 26238 35746 26290 35758
rect 29374 35810 29426 35822
rect 29374 35746 29426 35758
rect 32174 35810 32226 35822
rect 32174 35746 32226 35758
rect 34974 35810 35026 35822
rect 34974 35746 35026 35758
rect 36766 35810 36818 35822
rect 36766 35746 36818 35758
rect 37326 35810 37378 35822
rect 37326 35746 37378 35758
rect 38894 35810 38946 35822
rect 38894 35746 38946 35758
rect 39230 35810 39282 35822
rect 43486 35810 43538 35822
rect 41234 35758 41246 35810
rect 41298 35758 41310 35810
rect 39230 35746 39282 35758
rect 43486 35746 43538 35758
rect 48750 35810 48802 35822
rect 48750 35746 48802 35758
rect 49758 35810 49810 35822
rect 49758 35746 49810 35758
rect 50878 35810 50930 35822
rect 50878 35746 50930 35758
rect 53454 35810 53506 35822
rect 53454 35746 53506 35758
rect 53678 35810 53730 35822
rect 54574 35810 54626 35822
rect 54002 35758 54014 35810
rect 54066 35758 54078 35810
rect 53678 35746 53730 35758
rect 54574 35746 54626 35758
rect 55918 35810 55970 35822
rect 55918 35746 55970 35758
rect 10894 35698 10946 35710
rect 10894 35634 10946 35646
rect 20526 35698 20578 35710
rect 20526 35634 20578 35646
rect 22542 35698 22594 35710
rect 22542 35634 22594 35646
rect 23214 35698 23266 35710
rect 23214 35634 23266 35646
rect 40350 35698 40402 35710
rect 40350 35634 40402 35646
rect 43934 35698 43986 35710
rect 43934 35634 43986 35646
rect 57150 35698 57202 35710
rect 57150 35634 57202 35646
rect 57598 35698 57650 35710
rect 57598 35634 57650 35646
rect 34638 35586 34690 35598
rect 10098 35534 10110 35586
rect 10162 35534 10174 35586
rect 14130 35534 14142 35586
rect 14194 35534 14206 35586
rect 29026 35534 29038 35586
rect 29090 35534 29102 35586
rect 53554 35534 53566 35586
rect 53618 35534 53630 35586
rect 34638 35522 34690 35534
rect 17938 35422 17950 35474
rect 18002 35422 18014 35474
rect 22082 35422 22094 35474
rect 22146 35422 22158 35474
rect 22306 35422 22318 35474
rect 22370 35471 22382 35474
rect 22642 35471 22654 35474
rect 22370 35425 22654 35471
rect 22370 35422 22382 35425
rect 22642 35422 22654 35425
rect 22706 35471 22718 35474
rect 22866 35471 22878 35474
rect 22706 35425 22878 35471
rect 22706 35422 22718 35425
rect 22866 35422 22878 35425
rect 22930 35422 22942 35474
rect 55570 35422 55582 35474
rect 55634 35422 55646 35474
rect 56690 35422 56702 35474
rect 56754 35471 56766 35474
rect 57362 35471 57374 35474
rect 56754 35425 57374 35471
rect 56754 35422 56766 35425
rect 57362 35422 57374 35425
rect 57426 35422 57438 35474
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 55458 35086 55470 35138
rect 55522 35086 55534 35138
rect 13582 35026 13634 35038
rect 13582 34962 13634 34974
rect 5630 34914 5682 34926
rect 5630 34850 5682 34862
rect 15486 34914 15538 34926
rect 15486 34850 15538 34862
rect 19182 34914 19234 34926
rect 34750 34914 34802 34926
rect 22866 34862 22878 34914
rect 22930 34862 22942 34914
rect 19182 34850 19234 34862
rect 34750 34850 34802 34862
rect 35646 34914 35698 34926
rect 35646 34850 35698 34862
rect 38782 34914 38834 34926
rect 38782 34850 38834 34862
rect 44270 34914 44322 34926
rect 44270 34850 44322 34862
rect 46398 34914 46450 34926
rect 46398 34850 46450 34862
rect 53902 34914 53954 34926
rect 53902 34850 53954 34862
rect 1822 34802 1874 34814
rect 10446 34802 10498 34814
rect 2370 34750 2382 34802
rect 2434 34750 2446 34802
rect 9762 34750 9774 34802
rect 9826 34750 9838 34802
rect 1822 34738 1874 34750
rect 10446 34738 10498 34750
rect 13470 34802 13522 34814
rect 13470 34738 13522 34750
rect 13694 34802 13746 34814
rect 13694 34738 13746 34750
rect 15822 34802 15874 34814
rect 15822 34738 15874 34750
rect 18622 34802 18674 34814
rect 22542 34802 22594 34814
rect 20178 34750 20190 34802
rect 20242 34750 20254 34802
rect 18622 34738 18674 34750
rect 22542 34738 22594 34750
rect 23326 34802 23378 34814
rect 23326 34738 23378 34750
rect 23550 34802 23602 34814
rect 23550 34738 23602 34750
rect 24446 34802 24498 34814
rect 29262 34802 29314 34814
rect 27346 34750 27358 34802
rect 27410 34750 27422 34802
rect 24446 34738 24498 34750
rect 29262 34738 29314 34750
rect 32062 34802 32114 34814
rect 36094 34802 36146 34814
rect 33058 34750 33070 34802
rect 33122 34750 33134 34802
rect 32062 34738 32114 34750
rect 36094 34738 36146 34750
rect 37102 34802 37154 34814
rect 37102 34738 37154 34750
rect 37886 34802 37938 34814
rect 37886 34738 37938 34750
rect 40126 34802 40178 34814
rect 40126 34738 40178 34750
rect 41582 34802 41634 34814
rect 49646 34802 49698 34814
rect 52782 34802 52834 34814
rect 47730 34750 47742 34802
rect 47794 34750 47806 34802
rect 51538 34750 51550 34802
rect 51602 34750 51614 34802
rect 41582 34738 41634 34750
rect 49646 34738 49698 34750
rect 52782 34738 52834 34750
rect 53006 34802 53058 34814
rect 53006 34738 53058 34750
rect 53454 34802 53506 34814
rect 53454 34738 53506 34750
rect 55470 34802 55522 34814
rect 55470 34738 55522 34750
rect 57598 34802 57650 34814
rect 57598 34738 57650 34750
rect 58046 34802 58098 34814
rect 58046 34738 58098 34750
rect 8542 34690 8594 34702
rect 8542 34626 8594 34638
rect 9886 34690 9938 34702
rect 9886 34626 9938 34638
rect 12126 34690 12178 34702
rect 12126 34626 12178 34638
rect 16606 34690 16658 34702
rect 16606 34626 16658 34638
rect 19854 34690 19906 34702
rect 19854 34626 19906 34638
rect 20302 34690 20354 34702
rect 20302 34626 20354 34638
rect 22878 34690 22930 34702
rect 27134 34690 27186 34702
rect 23762 34638 23774 34690
rect 23826 34638 23838 34690
rect 22878 34626 22930 34638
rect 27134 34626 27186 34638
rect 27582 34690 27634 34702
rect 27582 34626 27634 34638
rect 30046 34690 30098 34702
rect 30046 34626 30098 34638
rect 33406 34690 33458 34702
rect 33406 34626 33458 34638
rect 34078 34690 34130 34702
rect 34078 34626 34130 34638
rect 35198 34690 35250 34702
rect 39454 34690 39506 34702
rect 37650 34638 37662 34690
rect 37714 34638 37726 34690
rect 35198 34626 35250 34638
rect 39454 34626 39506 34638
rect 42254 34690 42306 34702
rect 42254 34626 42306 34638
rect 45054 34690 45106 34702
rect 49758 34690 49810 34702
rect 48514 34638 48526 34690
rect 48578 34638 48590 34690
rect 45054 34626 45106 34638
rect 49758 34626 49810 34638
rect 50318 34690 50370 34702
rect 50318 34626 50370 34638
rect 51326 34690 51378 34702
rect 51326 34626 51378 34638
rect 51886 34690 51938 34702
rect 51886 34626 51938 34638
rect 55806 34690 55858 34702
rect 55806 34626 55858 34638
rect 57374 34690 57426 34702
rect 57374 34626 57426 34638
rect 4958 34578 5010 34590
rect 4610 34526 4622 34578
rect 4674 34526 4686 34578
rect 4958 34514 5010 34526
rect 5742 34578 5794 34590
rect 5742 34514 5794 34526
rect 8990 34578 9042 34590
rect 8990 34514 9042 34526
rect 9326 34578 9378 34590
rect 9326 34514 9378 34526
rect 10110 34578 10162 34590
rect 10110 34514 10162 34526
rect 23102 34578 23154 34590
rect 23102 34514 23154 34526
rect 23998 34578 24050 34590
rect 23998 34514 24050 34526
rect 24222 34578 24274 34590
rect 24222 34514 24274 34526
rect 25902 34578 25954 34590
rect 25902 34514 25954 34526
rect 28590 34578 28642 34590
rect 28590 34514 28642 34526
rect 32734 34578 32786 34590
rect 32734 34514 32786 34526
rect 33182 34578 33234 34590
rect 33182 34514 33234 34526
rect 40798 34578 40850 34590
rect 40798 34514 40850 34526
rect 43486 34578 43538 34590
rect 43486 34514 43538 34526
rect 50766 34578 50818 34590
rect 50766 34514 50818 34526
rect 52894 34578 52946 34590
rect 52894 34514 52946 34526
rect 9426 34414 9438 34466
rect 9490 34414 9502 34466
rect 12898 34414 12910 34466
rect 12962 34414 12974 34466
rect 19394 34414 19406 34466
rect 19458 34414 19470 34466
rect 28018 34414 28030 34466
rect 28082 34414 28094 34466
rect 50866 34414 50878 34466
rect 50930 34414 50942 34466
rect 1344 34298 58576 34332
rect 1344 34246 19838 34298
rect 19890 34246 19942 34298
rect 19994 34246 20046 34298
rect 20098 34246 50558 34298
rect 50610 34246 50662 34298
rect 50714 34246 50766 34298
rect 50818 34246 58576 34298
rect 1344 34212 58576 34246
rect 1810 34078 1822 34130
rect 1874 34127 1886 34130
rect 2706 34127 2718 34130
rect 1874 34081 2718 34127
rect 1874 34078 1886 34081
rect 2706 34078 2718 34081
rect 2770 34078 2782 34130
rect 12114 34078 12126 34130
rect 12178 34078 12190 34130
rect 12562 34078 12574 34130
rect 12626 34078 12638 34130
rect 46610 34078 46622 34130
rect 46674 34078 46686 34130
rect 50530 34078 50542 34130
rect 50594 34078 50606 34130
rect 15038 34018 15090 34030
rect 5506 33966 5518 34018
rect 5570 33966 5582 34018
rect 15038 33954 15090 33966
rect 22654 34018 22706 34030
rect 22654 33954 22706 33966
rect 25566 34018 25618 34030
rect 25566 33954 25618 33966
rect 26798 34018 26850 34030
rect 26798 33954 26850 33966
rect 28142 34018 28194 34030
rect 28142 33954 28194 33966
rect 29486 34018 29538 34030
rect 29486 33954 29538 33966
rect 36542 34018 36594 34030
rect 36542 33954 36594 33966
rect 36990 34018 37042 34030
rect 36990 33954 37042 33966
rect 37550 34018 37602 34030
rect 37550 33954 37602 33966
rect 38782 34018 38834 34030
rect 38782 33954 38834 33966
rect 39230 34018 39282 34030
rect 39230 33954 39282 33966
rect 39678 34018 39730 34030
rect 39678 33954 39730 33966
rect 40350 34018 40402 34030
rect 40350 33954 40402 33966
rect 41022 34018 41074 34030
rect 41022 33954 41074 33966
rect 41470 34018 41522 34030
rect 41470 33954 41522 33966
rect 42366 34018 42418 34030
rect 42366 33954 42418 33966
rect 53230 34018 53282 34030
rect 53230 33954 53282 33966
rect 55022 34018 55074 34030
rect 55022 33954 55074 33966
rect 55806 34018 55858 34030
rect 55806 33954 55858 33966
rect 58158 34018 58210 34030
rect 58158 33954 58210 33966
rect 10334 33906 10386 33918
rect 10334 33842 10386 33854
rect 11006 33906 11058 33918
rect 11006 33842 11058 33854
rect 13022 33906 13074 33918
rect 13022 33842 13074 33854
rect 13582 33906 13634 33918
rect 13582 33842 13634 33854
rect 13694 33906 13746 33918
rect 13694 33842 13746 33854
rect 14142 33906 14194 33918
rect 14142 33842 14194 33854
rect 14702 33906 14754 33918
rect 14702 33842 14754 33854
rect 16158 33906 16210 33918
rect 16158 33842 16210 33854
rect 18958 33906 19010 33918
rect 18958 33842 19010 33854
rect 19070 33906 19122 33918
rect 19070 33842 19122 33854
rect 25230 33906 25282 33918
rect 25230 33842 25282 33854
rect 27134 33906 27186 33918
rect 27134 33842 27186 33854
rect 34078 33906 34130 33918
rect 34078 33842 34130 33854
rect 35870 33906 35922 33918
rect 35870 33842 35922 33854
rect 36206 33906 36258 33918
rect 36206 33842 36258 33854
rect 42814 33906 42866 33918
rect 42814 33842 42866 33854
rect 43486 33906 43538 33918
rect 45614 33906 45666 33918
rect 44258 33854 44270 33906
rect 44322 33854 44334 33906
rect 43486 33842 43538 33854
rect 45614 33842 45666 33854
rect 46286 33906 46338 33918
rect 46286 33842 46338 33854
rect 47070 33906 47122 33918
rect 47070 33842 47122 33854
rect 47518 33906 47570 33918
rect 47518 33842 47570 33854
rect 49086 33906 49138 33918
rect 49086 33842 49138 33854
rect 49646 33906 49698 33918
rect 49646 33842 49698 33854
rect 52558 33906 52610 33918
rect 52558 33842 52610 33854
rect 52894 33906 52946 33918
rect 52894 33842 52946 33854
rect 54350 33906 54402 33918
rect 57710 33906 57762 33918
rect 56914 33854 56926 33906
rect 56978 33854 56990 33906
rect 54350 33842 54402 33854
rect 57710 33842 57762 33854
rect 2718 33794 2770 33806
rect 14478 33794 14530 33806
rect 3266 33742 3278 33794
rect 3330 33742 3342 33794
rect 2718 33730 2770 33742
rect 14478 33730 14530 33742
rect 15934 33794 15986 33806
rect 15934 33730 15986 33742
rect 16382 33794 16434 33806
rect 16382 33730 16434 33742
rect 18398 33794 18450 33806
rect 18398 33730 18450 33742
rect 21982 33794 22034 33806
rect 21982 33730 22034 33742
rect 27694 33794 27746 33806
rect 27694 33730 27746 33742
rect 28702 33794 28754 33806
rect 33518 33794 33570 33806
rect 32386 33742 32398 33794
rect 32450 33742 32462 33794
rect 28702 33730 28754 33742
rect 33518 33730 33570 33742
rect 34862 33794 34914 33806
rect 43150 33794 43202 33806
rect 35186 33742 35198 33794
rect 35250 33742 35262 33794
rect 34862 33730 34914 33742
rect 43150 33730 43202 33742
rect 43822 33794 43874 33806
rect 43822 33730 43874 33742
rect 44942 33794 44994 33806
rect 50206 33794 50258 33806
rect 49410 33742 49422 33794
rect 49474 33742 49486 33794
rect 44942 33730 44994 33742
rect 50206 33730 50258 33742
rect 51102 33794 51154 33806
rect 51102 33730 51154 33742
rect 51326 33794 51378 33806
rect 51326 33730 51378 33742
rect 51774 33794 51826 33806
rect 51774 33730 51826 33742
rect 52222 33794 52274 33806
rect 52222 33730 52274 33742
rect 53790 33794 53842 33806
rect 56018 33742 56030 33794
rect 56082 33742 56094 33794
rect 56690 33742 56702 33794
rect 56754 33742 56766 33794
rect 53790 33730 53842 33742
rect 1822 33682 1874 33694
rect 1822 33618 1874 33630
rect 2382 33682 2434 33694
rect 2382 33618 2434 33630
rect 5854 33682 5906 33694
rect 5854 33618 5906 33630
rect 14366 33682 14418 33694
rect 14366 33618 14418 33630
rect 21534 33682 21586 33694
rect 21534 33618 21586 33630
rect 24670 33682 24722 33694
rect 24670 33618 24722 33630
rect 26462 33682 26514 33694
rect 26462 33618 26514 33630
rect 32062 33682 32114 33694
rect 32062 33618 32114 33630
rect 34190 33682 34242 33694
rect 34190 33618 34242 33630
rect 35534 33682 35586 33694
rect 35534 33618 35586 33630
rect 41918 33682 41970 33694
rect 41918 33618 41970 33630
rect 48190 33682 48242 33694
rect 57362 33630 57374 33682
rect 57426 33630 57438 33682
rect 48190 33618 48242 33630
rect 27906 33518 27918 33570
rect 27970 33518 27982 33570
rect 31490 33518 31502 33570
rect 31554 33518 31566 33570
rect 16034 33406 16046 33458
rect 16098 33406 16110 33458
rect 17938 33406 17950 33458
rect 18002 33406 18014 33458
rect 27234 33406 27246 33458
rect 27298 33455 27310 33458
rect 27921 33455 27967 33518
rect 27298 33409 27967 33455
rect 27298 33406 27310 33409
rect 32498 33406 32510 33458
rect 32562 33406 32574 33458
rect 33058 33406 33070 33458
rect 33122 33406 33134 33458
rect 48626 33406 48638 33458
rect 48690 33406 48702 33458
rect 1344 33290 58576 33324
rect 1344 33238 4478 33290
rect 4530 33238 4582 33290
rect 4634 33238 4686 33290
rect 4738 33238 35198 33290
rect 35250 33238 35302 33290
rect 35354 33238 35406 33290
rect 35458 33238 58576 33290
rect 1344 33204 58576 33238
rect 4834 33070 4846 33122
rect 4898 33070 4910 33122
rect 34738 33070 34750 33122
rect 34802 33119 34814 33122
rect 35186 33119 35198 33122
rect 34802 33073 35198 33119
rect 34802 33070 34814 33073
rect 35186 33070 35198 33073
rect 35250 33070 35262 33122
rect 40786 33070 40798 33122
rect 40850 33070 40862 33122
rect 12462 33010 12514 33022
rect 12462 32946 12514 32958
rect 14702 33010 14754 33022
rect 14702 32946 14754 32958
rect 20414 33010 20466 33022
rect 20414 32946 20466 32958
rect 46062 33010 46114 33022
rect 50642 32958 50654 33010
rect 50706 33007 50718 33010
rect 51202 33007 51214 33010
rect 50706 32961 51214 33007
rect 50706 32958 50718 32961
rect 51202 32958 51214 32961
rect 51266 32958 51278 33010
rect 46062 32946 46114 32958
rect 22430 32898 22482 32910
rect 22430 32834 22482 32846
rect 28366 32898 28418 32910
rect 28366 32834 28418 32846
rect 31950 32898 32002 32910
rect 31950 32834 32002 32846
rect 34190 32898 34242 32910
rect 34190 32834 34242 32846
rect 34750 32898 34802 32910
rect 34750 32834 34802 32846
rect 35198 32898 35250 32910
rect 35198 32834 35250 32846
rect 35758 32898 35810 32910
rect 35758 32834 35810 32846
rect 37326 32898 37378 32910
rect 37326 32834 37378 32846
rect 39118 32898 39170 32910
rect 39118 32834 39170 32846
rect 43262 32898 43314 32910
rect 43262 32834 43314 32846
rect 45614 32898 45666 32910
rect 45614 32834 45666 32846
rect 50654 32898 50706 32910
rect 50654 32834 50706 32846
rect 51102 32898 51154 32910
rect 51102 32834 51154 32846
rect 56366 32898 56418 32910
rect 56366 32834 56418 32846
rect 57710 32898 57762 32910
rect 57710 32834 57762 32846
rect 58158 32898 58210 32910
rect 58158 32834 58210 32846
rect 15150 32786 15202 32798
rect 17278 32786 17330 32798
rect 4498 32734 4510 32786
rect 4562 32734 4574 32786
rect 11890 32734 11902 32786
rect 11954 32734 11966 32786
rect 15362 32734 15374 32786
rect 15426 32734 15438 32786
rect 15150 32722 15202 32734
rect 17278 32722 17330 32734
rect 17614 32786 17666 32798
rect 17614 32722 17666 32734
rect 18510 32786 18562 32798
rect 18510 32722 18562 32734
rect 23214 32786 23266 32798
rect 23214 32722 23266 32734
rect 26014 32786 26066 32798
rect 26014 32722 26066 32734
rect 27022 32786 27074 32798
rect 27022 32722 27074 32734
rect 27246 32786 27298 32798
rect 27246 32722 27298 32734
rect 27806 32786 27858 32798
rect 27806 32722 27858 32734
rect 32174 32786 32226 32798
rect 32174 32722 32226 32734
rect 33518 32786 33570 32798
rect 33518 32722 33570 32734
rect 37886 32786 37938 32798
rect 37886 32722 37938 32734
rect 38110 32786 38162 32798
rect 38110 32722 38162 32734
rect 40238 32786 40290 32798
rect 40238 32722 40290 32734
rect 42814 32786 42866 32798
rect 48974 32786 49026 32798
rect 46610 32734 46622 32786
rect 46674 32734 46686 32786
rect 42814 32722 42866 32734
rect 48974 32722 49026 32734
rect 49310 32786 49362 32798
rect 49310 32722 49362 32734
rect 53230 32786 53282 32798
rect 53230 32722 53282 32734
rect 53566 32786 53618 32798
rect 53566 32722 53618 32734
rect 53902 32786 53954 32798
rect 57262 32786 57314 32798
rect 56690 32734 56702 32786
rect 56754 32734 56766 32786
rect 53902 32722 53954 32734
rect 57262 32722 57314 32734
rect 4398 32674 4450 32686
rect 4398 32610 4450 32622
rect 12798 32674 12850 32686
rect 12798 32610 12850 32622
rect 14142 32674 14194 32686
rect 14142 32610 14194 32622
rect 15710 32674 15762 32686
rect 15710 32610 15762 32622
rect 16942 32674 16994 32686
rect 16942 32610 16994 32622
rect 19070 32674 19122 32686
rect 19070 32610 19122 32622
rect 20750 32674 20802 32686
rect 20750 32610 20802 32622
rect 23998 32674 24050 32686
rect 23998 32610 24050 32622
rect 26350 32674 26402 32686
rect 26350 32610 26402 32622
rect 26686 32674 26738 32686
rect 26686 32610 26738 32622
rect 27582 32674 27634 32686
rect 27582 32610 27634 32622
rect 32510 32674 32562 32686
rect 32510 32610 32562 32622
rect 34078 32674 34130 32686
rect 34078 32610 34130 32622
rect 40126 32674 40178 32686
rect 40126 32610 40178 32622
rect 41918 32674 41970 32686
rect 52894 32674 52946 32686
rect 55022 32674 55074 32686
rect 46946 32622 46958 32674
rect 47010 32622 47022 32674
rect 54338 32622 54350 32674
rect 54402 32622 54414 32674
rect 41918 32610 41970 32622
rect 52894 32610 52946 32622
rect 55022 32610 55074 32622
rect 55694 32674 55746 32686
rect 55694 32610 55746 32622
rect 56814 32674 56866 32686
rect 57138 32622 57150 32674
rect 57202 32622 57214 32674
rect 56814 32610 56866 32622
rect 4958 32562 5010 32574
rect 4958 32498 5010 32510
rect 14478 32562 14530 32574
rect 14478 32498 14530 32510
rect 17950 32562 18002 32574
rect 17950 32498 18002 32510
rect 19742 32562 19794 32574
rect 19742 32498 19794 32510
rect 22766 32562 22818 32574
rect 22766 32498 22818 32510
rect 22878 32562 22930 32574
rect 22878 32498 22930 32510
rect 26798 32562 26850 32574
rect 32846 32562 32898 32574
rect 31938 32510 31950 32562
rect 32002 32510 32014 32562
rect 26798 32498 26850 32510
rect 32846 32498 32898 32510
rect 43710 32562 43762 32574
rect 43710 32498 43762 32510
rect 44158 32562 44210 32574
rect 44158 32498 44210 32510
rect 45166 32562 45218 32574
rect 45166 32498 45218 32510
rect 52110 32562 52162 32574
rect 52110 32498 52162 32510
rect 56254 32562 56306 32574
rect 56254 32498 56306 32510
rect 11778 32398 11790 32450
rect 11842 32398 11854 32450
rect 27682 32398 27694 32450
rect 27746 32398 27758 32450
rect 33058 32398 33070 32450
rect 33122 32398 33134 32450
rect 38434 32398 38446 32450
rect 38498 32398 38510 32450
rect 1344 32282 58576 32316
rect 1344 32230 19838 32282
rect 19890 32230 19942 32282
rect 19994 32230 20046 32282
rect 20098 32230 50558 32282
rect 50610 32230 50662 32282
rect 50714 32230 50766 32282
rect 50818 32230 58576 32282
rect 1344 32196 58576 32230
rect 41234 32062 41246 32114
rect 41298 32062 41310 32114
rect 13470 32002 13522 32014
rect 5506 31950 5518 32002
rect 5570 31950 5582 32002
rect 13470 31938 13522 31950
rect 19742 32002 19794 32014
rect 19742 31938 19794 31950
rect 22878 32002 22930 32014
rect 22878 31938 22930 31950
rect 23662 32002 23714 32014
rect 23662 31938 23714 31950
rect 27918 32002 27970 32014
rect 27918 31938 27970 31950
rect 28366 32002 28418 32014
rect 28366 31938 28418 31950
rect 32174 32002 32226 32014
rect 32174 31938 32226 31950
rect 44382 32002 44434 32014
rect 44382 31938 44434 31950
rect 51550 32002 51602 32014
rect 52882 31950 52894 32002
rect 52946 31950 52958 32002
rect 51550 31938 51602 31950
rect 2382 31890 2434 31902
rect 2382 31826 2434 31838
rect 5854 31890 5906 31902
rect 5854 31826 5906 31838
rect 14366 31890 14418 31902
rect 14366 31826 14418 31838
rect 15934 31890 15986 31902
rect 15934 31826 15986 31838
rect 16046 31890 16098 31902
rect 16046 31826 16098 31838
rect 20974 31890 21026 31902
rect 20974 31826 21026 31838
rect 21086 31890 21138 31902
rect 21086 31826 21138 31838
rect 21870 31890 21922 31902
rect 21870 31826 21922 31838
rect 22542 31890 22594 31902
rect 22542 31826 22594 31838
rect 23886 31890 23938 31902
rect 23886 31826 23938 31838
rect 24110 31890 24162 31902
rect 24110 31826 24162 31838
rect 25342 31890 25394 31902
rect 25342 31826 25394 31838
rect 25566 31890 25618 31902
rect 26238 31890 26290 31902
rect 25890 31838 25902 31890
rect 25954 31838 25966 31890
rect 25566 31826 25618 31838
rect 26238 31826 26290 31838
rect 26350 31890 26402 31902
rect 27582 31890 27634 31902
rect 26350 31826 26402 31838
rect 27022 31834 27074 31846
rect 2718 31778 2770 31790
rect 10782 31778 10834 31790
rect 13918 31778 13970 31790
rect 15374 31778 15426 31790
rect 3266 31726 3278 31778
rect 3330 31726 3342 31778
rect 11330 31726 11342 31778
rect 11394 31726 11406 31778
rect 14466 31726 14478 31778
rect 14530 31726 14542 31778
rect 2718 31714 2770 31726
rect 10782 31714 10834 31726
rect 13918 31714 13970 31726
rect 15374 31714 15426 31726
rect 20414 31778 20466 31790
rect 20414 31714 20466 31726
rect 20862 31778 20914 31790
rect 20862 31714 20914 31726
rect 21310 31784 21362 31796
rect 23214 31778 23266 31790
rect 27582 31826 27634 31838
rect 31278 31890 31330 31902
rect 31278 31826 31330 31838
rect 31838 31890 31890 31902
rect 31838 31826 31890 31838
rect 32510 31890 32562 31902
rect 32510 31826 32562 31838
rect 33294 31890 33346 31902
rect 33294 31826 33346 31838
rect 35758 31890 35810 31902
rect 38446 31890 38498 31902
rect 37762 31838 37774 31890
rect 37826 31838 37838 31890
rect 35758 31826 35810 31838
rect 38446 31826 38498 31838
rect 39118 31890 39170 31902
rect 39118 31826 39170 31838
rect 41694 31890 41746 31902
rect 41694 31826 41746 31838
rect 42814 31890 42866 31902
rect 42814 31826 42866 31838
rect 43374 31890 43426 31902
rect 43374 31826 43426 31838
rect 44046 31890 44098 31902
rect 44046 31826 44098 31838
rect 45390 31890 45442 31902
rect 47182 31890 47234 31902
rect 46610 31838 46622 31890
rect 46674 31838 46686 31890
rect 45390 31826 45442 31838
rect 47182 31826 47234 31838
rect 51998 31890 52050 31902
rect 51998 31826 52050 31838
rect 53342 31890 53394 31902
rect 53342 31826 53394 31838
rect 33518 31790 33570 31802
rect 21310 31720 21362 31732
rect 21746 31726 21758 31778
rect 21810 31726 21822 31778
rect 24322 31726 24334 31778
rect 24386 31726 24398 31778
rect 25218 31726 25230 31778
rect 25282 31726 25294 31778
rect 27022 31770 27074 31782
rect 27246 31778 27298 31790
rect 23214 31714 23266 31726
rect 27246 31714 27298 31726
rect 31614 31778 31666 31790
rect 31614 31714 31666 31726
rect 33070 31778 33122 31790
rect 34750 31778 34802 31790
rect 33518 31726 33570 31738
rect 34402 31726 34414 31778
rect 34466 31726 34478 31778
rect 33070 31714 33122 31726
rect 34750 31714 34802 31726
rect 36318 31778 36370 31790
rect 36318 31714 36370 31726
rect 36654 31778 36706 31790
rect 36654 31714 36706 31726
rect 36990 31778 37042 31790
rect 36990 31714 37042 31726
rect 37326 31778 37378 31790
rect 37326 31714 37378 31726
rect 40910 31778 40962 31790
rect 46398 31778 46450 31790
rect 43474 31726 43486 31778
rect 43538 31726 43550 31778
rect 40910 31714 40962 31726
rect 46398 31714 46450 31726
rect 47966 31778 48018 31790
rect 47966 31714 48018 31726
rect 49870 31778 49922 31790
rect 49870 31714 49922 31726
rect 53454 31778 53506 31790
rect 55010 31753 55022 31805
rect 55074 31753 55086 31805
rect 53454 31714 53506 31726
rect 10446 31666 10498 31678
rect 10446 31602 10498 31614
rect 14926 31666 14978 31678
rect 14926 31602 14978 31614
rect 16830 31666 16882 31678
rect 30830 31666 30882 31678
rect 23650 31614 23662 31666
rect 23714 31663 23726 31666
rect 24546 31663 24558 31666
rect 23714 31617 24558 31663
rect 23714 31614 23726 31617
rect 24546 31614 24558 31617
rect 24610 31614 24622 31666
rect 16830 31602 16882 31614
rect 30830 31602 30882 31614
rect 39902 31666 39954 31678
rect 39902 31602 39954 31614
rect 40350 31666 40402 31678
rect 46846 31666 46898 31678
rect 45378 31614 45390 31666
rect 45442 31614 45454 31666
rect 40350 31602 40402 31614
rect 46846 31602 46898 31614
rect 47518 31666 47570 31678
rect 47518 31602 47570 31614
rect 49534 31666 49586 31678
rect 49534 31602 49586 31614
rect 50206 31666 50258 31678
rect 50206 31602 50258 31614
rect 51102 31666 51154 31678
rect 51102 31602 51154 31614
rect 52446 31666 52498 31678
rect 52446 31602 52498 31614
rect 55806 31666 55858 31678
rect 55806 31602 55858 31614
rect 56702 31666 56754 31678
rect 56702 31602 56754 31614
rect 57150 31666 57202 31678
rect 57150 31602 57202 31614
rect 25790 31554 25842 31566
rect 17714 31502 17726 31554
rect 17778 31502 17790 31554
rect 25790 31490 25842 31502
rect 31502 31554 31554 31566
rect 45714 31502 45726 31554
rect 45778 31502 45790 31554
rect 31502 31490 31554 31502
rect 26898 31390 26910 31442
rect 26962 31390 26974 31442
rect 33394 31390 33406 31442
rect 33458 31390 33470 31442
rect 42466 31390 42478 31442
rect 42530 31390 42542 31442
rect 1344 31274 58576 31308
rect 1344 31222 4478 31274
rect 4530 31222 4582 31274
rect 4634 31222 4686 31274
rect 4738 31222 35198 31274
rect 35250 31222 35302 31274
rect 35354 31222 35406 31274
rect 35458 31222 58576 31274
rect 1344 31188 58576 31222
rect 17266 31054 17278 31106
rect 17330 31054 17342 31106
rect 18722 31054 18734 31106
rect 18786 31054 18798 31106
rect 23874 31054 23886 31106
rect 23938 31054 23950 31106
rect 25106 31054 25118 31106
rect 25170 31054 25182 31106
rect 27570 31054 27582 31106
rect 27634 31054 27646 31106
rect 32946 31054 32958 31106
rect 33010 31054 33022 31106
rect 15038 30994 15090 31006
rect 15038 30930 15090 30942
rect 26126 30994 26178 31006
rect 32961 30991 33007 31054
rect 32961 30945 33221 30991
rect 26126 30930 26178 30942
rect 5630 30882 5682 30894
rect 5630 30818 5682 30830
rect 16158 30882 16210 30894
rect 31166 30882 31218 30894
rect 32846 30882 32898 30894
rect 28242 30830 28254 30882
rect 28306 30830 28318 30882
rect 32274 30830 32286 30882
rect 32338 30879 32350 30882
rect 32722 30879 32734 30882
rect 32338 30833 32734 30879
rect 32338 30830 32350 30833
rect 32722 30830 32734 30833
rect 32786 30830 32798 30882
rect 33175 30879 33221 30945
rect 36306 30942 36318 30994
rect 36370 30942 36382 30994
rect 33854 30882 33906 30894
rect 33506 30879 33518 30882
rect 33175 30833 33518 30879
rect 33506 30830 33518 30833
rect 33570 30830 33582 30882
rect 16158 30818 16210 30830
rect 31166 30818 31218 30830
rect 32846 30818 32898 30830
rect 33854 30818 33906 30830
rect 35534 30882 35586 30894
rect 35534 30818 35586 30830
rect 40574 30882 40626 30894
rect 40574 30818 40626 30830
rect 43598 30882 43650 30894
rect 43598 30818 43650 30830
rect 44046 30882 44098 30894
rect 53678 30882 53730 30894
rect 45602 30830 45614 30882
rect 45666 30879 45678 30882
rect 46386 30879 46398 30882
rect 45666 30833 46398 30879
rect 45666 30830 45678 30833
rect 46386 30830 46398 30833
rect 46450 30830 46462 30882
rect 44046 30818 44098 30830
rect 53678 30818 53730 30830
rect 55582 30882 55634 30894
rect 55582 30818 55634 30830
rect 1822 30770 1874 30782
rect 9662 30770 9714 30782
rect 19182 30770 19234 30782
rect 23550 30770 23602 30782
rect 2370 30718 2382 30770
rect 2434 30718 2446 30770
rect 10210 30718 10222 30770
rect 10274 30718 10286 30770
rect 14578 30718 14590 30770
rect 14642 30718 14654 30770
rect 17938 30718 17950 30770
rect 18002 30718 18014 30770
rect 19394 30718 19406 30770
rect 19458 30718 19470 30770
rect 1822 30706 1874 30718
rect 9662 30706 9714 30718
rect 19182 30706 19234 30718
rect 23550 30706 23602 30718
rect 23774 30770 23826 30782
rect 23774 30706 23826 30718
rect 23998 30770 24050 30782
rect 23998 30706 24050 30718
rect 24222 30770 24274 30782
rect 24222 30706 24274 30718
rect 24558 30770 24610 30782
rect 24558 30706 24610 30718
rect 24782 30770 24834 30782
rect 24782 30706 24834 30718
rect 26462 30770 26514 30782
rect 26462 30706 26514 30718
rect 27358 30770 27410 30782
rect 27358 30706 27410 30718
rect 27918 30770 27970 30782
rect 27918 30706 27970 30718
rect 28590 30770 28642 30782
rect 32734 30770 32786 30782
rect 30706 30718 30718 30770
rect 30770 30718 30782 30770
rect 28590 30706 28642 30718
rect 32734 30706 32786 30718
rect 33182 30770 33234 30782
rect 33182 30706 33234 30718
rect 33518 30770 33570 30782
rect 33518 30706 33570 30718
rect 33966 30770 34018 30782
rect 33966 30706 34018 30718
rect 35646 30770 35698 30782
rect 35646 30706 35698 30718
rect 37662 30770 37714 30782
rect 37662 30706 37714 30718
rect 39678 30770 39730 30782
rect 39678 30706 39730 30718
rect 41134 30770 41186 30782
rect 41134 30706 41186 30718
rect 41358 30770 41410 30782
rect 41358 30706 41410 30718
rect 41806 30770 41858 30782
rect 41806 30706 41858 30718
rect 44942 30770 44994 30782
rect 44942 30706 44994 30718
rect 45166 30770 45218 30782
rect 45166 30706 45218 30718
rect 45390 30770 45442 30782
rect 45390 30706 45442 30718
rect 45950 30770 46002 30782
rect 45950 30706 46002 30718
rect 46174 30770 46226 30782
rect 46174 30706 46226 30718
rect 14030 30658 14082 30670
rect 14030 30594 14082 30606
rect 14478 30658 14530 30670
rect 14478 30594 14530 30606
rect 15486 30658 15538 30670
rect 15486 30594 15538 30606
rect 16046 30658 16098 30670
rect 16046 30594 16098 30606
rect 17726 30658 17778 30670
rect 17726 30594 17778 30606
rect 18286 30658 18338 30670
rect 18286 30594 18338 30606
rect 19630 30658 19682 30670
rect 19630 30594 19682 30606
rect 22766 30658 22818 30670
rect 22766 30594 22818 30606
rect 25006 30658 25058 30670
rect 25006 30594 25058 30606
rect 25566 30658 25618 30670
rect 25566 30594 25618 30606
rect 25678 30658 25730 30670
rect 25678 30594 25730 30606
rect 26350 30658 26402 30670
rect 26350 30594 26402 30606
rect 26910 30658 26962 30670
rect 26910 30594 26962 30606
rect 27022 30658 27074 30670
rect 27022 30594 27074 30606
rect 27694 30658 27746 30670
rect 27694 30594 27746 30606
rect 28366 30658 28418 30670
rect 28366 30594 28418 30606
rect 30830 30658 30882 30670
rect 30830 30594 30882 30606
rect 31390 30658 31442 30670
rect 31390 30594 31442 30606
rect 32062 30658 32114 30670
rect 32062 30594 32114 30606
rect 32958 30658 33010 30670
rect 32958 30594 33010 30606
rect 33742 30658 33794 30670
rect 33742 30594 33794 30606
rect 34414 30658 34466 30670
rect 34414 30594 34466 30606
rect 36990 30658 37042 30670
rect 36990 30594 37042 30606
rect 39230 30658 39282 30670
rect 39230 30594 39282 30606
rect 45614 30658 45666 30670
rect 45614 30594 45666 30606
rect 46622 30658 46674 30670
rect 46622 30594 46674 30606
rect 49310 30658 49362 30670
rect 49310 30594 49362 30606
rect 53006 30658 53058 30670
rect 53006 30594 53058 30606
rect 53566 30658 53618 30670
rect 53566 30594 53618 30606
rect 54238 30658 54290 30670
rect 54238 30594 54290 30606
rect 54686 30658 54738 30670
rect 54686 30594 54738 30606
rect 4958 30546 5010 30558
rect 4610 30494 4622 30546
rect 4674 30494 4686 30546
rect 4958 30482 5010 30494
rect 5742 30546 5794 30558
rect 5742 30482 5794 30494
rect 6078 30546 6130 30558
rect 6078 30482 6130 30494
rect 9326 30546 9378 30558
rect 12798 30546 12850 30558
rect 12450 30494 12462 30546
rect 12514 30494 12526 30546
rect 9326 30482 9378 30494
rect 12798 30482 12850 30494
rect 23102 30546 23154 30558
rect 26686 30546 26738 30558
rect 26002 30494 26014 30546
rect 26066 30494 26078 30546
rect 23102 30482 23154 30494
rect 26686 30482 26738 30494
rect 29262 30546 29314 30558
rect 29262 30482 29314 30494
rect 29710 30546 29762 30558
rect 29710 30482 29762 30494
rect 31726 30546 31778 30558
rect 31726 30482 31778 30494
rect 34750 30546 34802 30558
rect 34750 30482 34802 30494
rect 37326 30546 37378 30558
rect 43150 30546 43202 30558
rect 39106 30494 39118 30546
rect 39170 30494 39182 30546
rect 37326 30482 37378 30494
rect 43150 30482 43202 30494
rect 45054 30546 45106 30558
rect 45054 30482 45106 30494
rect 47070 30546 47122 30558
rect 47070 30482 47122 30494
rect 48302 30546 48354 30558
rect 48302 30482 48354 30494
rect 48750 30546 48802 30558
rect 48750 30482 48802 30494
rect 49982 30546 50034 30558
rect 49982 30482 50034 30494
rect 55134 30546 55186 30558
rect 55134 30482 55186 30494
rect 56030 30546 56082 30558
rect 56030 30482 56082 30494
rect 6178 30382 6190 30434
rect 6242 30382 6254 30434
rect 13570 30382 13582 30434
rect 13634 30382 13646 30434
rect 31042 30382 31054 30434
rect 31106 30382 31118 30434
rect 37986 30382 37998 30434
rect 38050 30382 38062 30434
rect 51874 30382 51886 30434
rect 51938 30382 51950 30434
rect 52546 30382 52558 30434
rect 52610 30382 52622 30434
rect 54898 30382 54910 30434
rect 54962 30431 54974 30434
rect 55794 30431 55806 30434
rect 54962 30385 55806 30431
rect 54962 30382 54974 30385
rect 55794 30382 55806 30385
rect 55858 30382 55870 30434
rect 1344 30266 58576 30300
rect 1344 30214 19838 30266
rect 19890 30214 19942 30266
rect 19994 30214 20046 30266
rect 20098 30214 50558 30266
rect 50610 30214 50662 30266
rect 50714 30214 50766 30266
rect 50818 30214 58576 30266
rect 1344 30180 58576 30214
rect 3826 30046 3838 30098
rect 3890 30046 3902 30098
rect 10322 30046 10334 30098
rect 10386 30046 10398 30098
rect 14242 30046 14254 30098
rect 14306 30046 14318 30098
rect 24434 30046 24446 30098
rect 24498 30046 24510 30098
rect 25554 30046 25566 30098
rect 25618 30046 25630 30098
rect 26450 30046 26462 30098
rect 26514 30046 26526 30098
rect 28130 30046 28142 30098
rect 28194 30046 28206 30098
rect 48626 30046 48638 30098
rect 48690 30046 48702 30098
rect 50530 30046 50542 30098
rect 50594 30095 50606 30098
rect 51090 30095 51102 30098
rect 50594 30049 51102 30095
rect 50594 30046 50606 30049
rect 51090 30046 51102 30049
rect 51154 30046 51166 30098
rect 4734 29986 4786 29998
rect 4734 29922 4786 29934
rect 5182 29986 5234 29998
rect 5182 29922 5234 29934
rect 8542 29986 8594 29998
rect 8542 29922 8594 29934
rect 13470 29986 13522 29998
rect 13470 29922 13522 29934
rect 13918 29986 13970 29998
rect 13918 29922 13970 29934
rect 24334 29986 24386 29998
rect 24334 29922 24386 29934
rect 27806 29986 27858 29998
rect 27806 29922 27858 29934
rect 30158 29986 30210 29998
rect 30158 29922 30210 29934
rect 31726 29986 31778 29998
rect 31726 29922 31778 29934
rect 32174 29986 32226 29998
rect 32174 29922 32226 29934
rect 34190 29986 34242 29998
rect 34190 29922 34242 29934
rect 36654 29986 36706 29998
rect 36654 29922 36706 29934
rect 37998 29986 38050 29998
rect 37998 29922 38050 29934
rect 38446 29986 38498 29998
rect 38446 29922 38498 29934
rect 38894 29986 38946 29998
rect 38894 29922 38946 29934
rect 39902 29986 39954 29998
rect 39902 29922 39954 29934
rect 40350 29986 40402 29998
rect 40350 29922 40402 29934
rect 43374 29986 43426 29998
rect 43374 29922 43426 29934
rect 45166 29986 45218 29998
rect 45166 29922 45218 29934
rect 46398 29986 46450 29998
rect 46398 29922 46450 29934
rect 15262 29874 15314 29886
rect 15262 29810 15314 29822
rect 23886 29874 23938 29886
rect 23886 29810 23938 29822
rect 24222 29874 24274 29886
rect 24222 29810 24274 29822
rect 24782 29874 24834 29886
rect 24782 29810 24834 29822
rect 25230 29874 25282 29886
rect 25230 29810 25282 29822
rect 25566 29874 25618 29886
rect 25566 29810 25618 29822
rect 25678 29874 25730 29886
rect 26910 29874 26962 29886
rect 26562 29822 26574 29874
rect 26626 29822 26638 29874
rect 25678 29810 25730 29822
rect 26910 29810 26962 29822
rect 27022 29874 27074 29886
rect 27022 29810 27074 29822
rect 27470 29874 27522 29886
rect 30494 29874 30546 29886
rect 29586 29822 29598 29874
rect 29650 29822 29662 29874
rect 27470 29810 27522 29822
rect 30494 29810 30546 29822
rect 31054 29874 31106 29886
rect 31054 29810 31106 29822
rect 31390 29874 31442 29886
rect 31390 29810 31442 29822
rect 32510 29874 32562 29886
rect 32510 29810 32562 29822
rect 34526 29874 34578 29886
rect 34526 29810 34578 29822
rect 35758 29874 35810 29886
rect 35758 29810 35810 29822
rect 36206 29874 36258 29886
rect 36206 29810 36258 29822
rect 41246 29874 41298 29886
rect 41246 29810 41298 29822
rect 41694 29874 41746 29886
rect 41694 29810 41746 29822
rect 42366 29874 42418 29886
rect 42366 29810 42418 29822
rect 42702 29874 42754 29886
rect 42702 29810 42754 29822
rect 43038 29874 43090 29886
rect 49646 29874 49698 29886
rect 43810 29822 43822 29874
rect 43874 29822 43886 29874
rect 43038 29810 43090 29822
rect 49646 29810 49698 29822
rect 51326 29874 51378 29886
rect 51326 29810 51378 29822
rect 51662 29874 51714 29886
rect 51662 29810 51714 29822
rect 51998 29874 52050 29886
rect 54126 29874 54178 29886
rect 52770 29822 52782 29874
rect 52834 29822 52846 29874
rect 51998 29810 52050 29822
rect 54126 29810 54178 29822
rect 7870 29762 7922 29774
rect 10782 29762 10834 29774
rect 14702 29762 14754 29774
rect 26126 29762 26178 29774
rect 3378 29710 3390 29762
rect 3442 29710 3454 29762
rect 3714 29710 3726 29762
rect 3778 29710 3790 29762
rect 4162 29710 4174 29762
rect 4226 29710 4238 29762
rect 7298 29710 7310 29762
rect 7362 29710 7374 29762
rect 8978 29710 8990 29762
rect 9042 29710 9054 29762
rect 9986 29710 9998 29762
rect 10050 29710 10062 29762
rect 10434 29710 10446 29762
rect 10498 29710 10510 29762
rect 11330 29710 11342 29762
rect 11394 29710 11406 29762
rect 14914 29710 14926 29762
rect 14978 29710 14990 29762
rect 7870 29698 7922 29710
rect 10782 29698 10834 29710
rect 14702 29698 14754 29710
rect 26126 29698 26178 29710
rect 26238 29762 26290 29774
rect 26238 29698 26290 29710
rect 28478 29762 28530 29774
rect 28478 29698 28530 29710
rect 29262 29762 29314 29774
rect 29262 29698 29314 29710
rect 29934 29762 29986 29774
rect 29934 29698 29986 29710
rect 33070 29762 33122 29774
rect 33070 29698 33122 29710
rect 33182 29762 33234 29774
rect 33182 29698 33234 29710
rect 33294 29762 33346 29774
rect 33294 29698 33346 29710
rect 33518 29762 33570 29774
rect 33518 29698 33570 29710
rect 33742 29762 33794 29774
rect 33742 29698 33794 29710
rect 34862 29762 34914 29774
rect 34862 29698 34914 29710
rect 35422 29762 35474 29774
rect 35422 29698 35474 29710
rect 35534 29762 35586 29774
rect 44494 29762 44546 29774
rect 41458 29710 41470 29762
rect 41522 29710 41534 29762
rect 35534 29698 35586 29710
rect 44494 29698 44546 29710
rect 49086 29762 49138 29774
rect 52334 29762 52386 29774
rect 49298 29710 49310 29762
rect 49362 29710 49374 29762
rect 49086 29698 49138 29710
rect 52334 29698 52386 29710
rect 53454 29762 53506 29774
rect 53454 29698 53506 29710
rect 1822 29650 1874 29662
rect 1822 29586 1874 29598
rect 2942 29650 2994 29662
rect 2942 29586 2994 29598
rect 28926 29650 28978 29662
rect 28926 29586 28978 29598
rect 29598 29650 29650 29662
rect 29598 29586 29650 29598
rect 37102 29650 37154 29662
rect 37102 29586 37154 29598
rect 37550 29650 37602 29662
rect 37550 29586 37602 29598
rect 39454 29650 39506 29662
rect 39454 29586 39506 29598
rect 45950 29650 46002 29662
rect 45950 29586 46002 29598
rect 48190 29650 48242 29662
rect 48190 29586 48242 29598
rect 50542 29650 50594 29662
rect 50542 29586 50594 29598
rect 50990 29650 51042 29662
rect 50990 29586 51042 29598
rect 54910 29650 54962 29662
rect 54910 29586 54962 29598
rect 55806 29650 55858 29662
rect 55806 29586 55858 29598
rect 35198 29538 35250 29550
rect 35198 29474 35250 29486
rect 3266 29374 3278 29426
rect 3330 29374 3342 29426
rect 4274 29374 4286 29426
rect 4338 29374 4350 29426
rect 8866 29374 8878 29426
rect 8930 29374 8942 29426
rect 9874 29374 9886 29426
rect 9938 29374 9950 29426
rect 40786 29374 40798 29426
rect 40850 29374 40862 29426
rect 1344 29258 58576 29292
rect 1344 29206 4478 29258
rect 4530 29206 4582 29258
rect 4634 29206 4686 29258
rect 4738 29206 35198 29258
rect 35250 29206 35302 29258
rect 35354 29206 35406 29258
rect 35458 29206 58576 29258
rect 1344 29172 58576 29206
rect 13458 29038 13470 29090
rect 13522 29038 13534 29090
rect 27122 29038 27134 29090
rect 27186 29087 27198 29090
rect 27682 29087 27694 29090
rect 27186 29041 27694 29087
rect 27186 29038 27198 29041
rect 27682 29038 27694 29041
rect 27746 29038 27758 29090
rect 40114 29038 40126 29090
rect 40178 29038 40190 29090
rect 50866 29038 50878 29090
rect 50930 29038 50942 29090
rect 54002 29038 54014 29090
rect 54066 29038 54078 29090
rect 1922 28926 1934 28978
rect 1986 28926 1998 28978
rect 8754 28926 8766 28978
rect 8818 28926 8830 28978
rect 12786 28926 12798 28978
rect 12850 28926 12862 28978
rect 35634 28926 35646 28978
rect 35698 28975 35710 28978
rect 36418 28975 36430 28978
rect 35698 28929 36430 28975
rect 35698 28926 35710 28929
rect 36418 28926 36430 28929
rect 36482 28926 36494 28978
rect 9326 28866 9378 28878
rect 9326 28802 9378 28814
rect 15150 28866 15202 28878
rect 15150 28802 15202 28814
rect 24782 28866 24834 28878
rect 27582 28866 27634 28878
rect 25218 28814 25230 28866
rect 25282 28863 25294 28866
rect 26002 28863 26014 28866
rect 25282 28817 26014 28863
rect 25282 28814 25294 28817
rect 26002 28814 26014 28817
rect 26066 28814 26078 28866
rect 24782 28802 24834 28814
rect 27582 28802 27634 28814
rect 31502 28866 31554 28878
rect 31502 28802 31554 28814
rect 35198 28866 35250 28878
rect 35198 28802 35250 28814
rect 35646 28866 35698 28878
rect 35646 28802 35698 28814
rect 36094 28866 36146 28878
rect 36094 28802 36146 28814
rect 37102 28866 37154 28878
rect 37102 28802 37154 28814
rect 39118 28866 39170 28878
rect 39118 28802 39170 28814
rect 39902 28866 39954 28878
rect 39902 28802 39954 28814
rect 41246 28866 41298 28878
rect 41246 28802 41298 28814
rect 43374 28866 43426 28878
rect 43374 28802 43426 28814
rect 43822 28866 43874 28878
rect 43822 28802 43874 28814
rect 44270 28866 44322 28878
rect 54014 28866 54066 28878
rect 46162 28814 46174 28866
rect 46226 28814 46238 28866
rect 49858 28814 49870 28866
rect 49922 28814 49934 28866
rect 44270 28802 44322 28814
rect 54014 28802 54066 28814
rect 5070 28754 5122 28766
rect 4498 28702 4510 28754
rect 4562 28702 4574 28754
rect 5070 28690 5122 28702
rect 5630 28754 5682 28766
rect 9662 28754 9714 28766
rect 14030 28754 14082 28766
rect 6178 28702 6190 28754
rect 6242 28702 6254 28754
rect 10210 28702 10222 28754
rect 10274 28702 10286 28754
rect 13570 28702 13582 28754
rect 13634 28702 13646 28754
rect 5630 28690 5682 28702
rect 9662 28690 9714 28702
rect 14030 28690 14082 28702
rect 14478 28754 14530 28766
rect 14478 28690 14530 28702
rect 20302 28754 20354 28766
rect 20302 28690 20354 28702
rect 21310 28754 21362 28766
rect 21310 28690 21362 28702
rect 22318 28754 22370 28766
rect 22318 28690 22370 28702
rect 24446 28754 24498 28766
rect 26350 28754 26402 28766
rect 25106 28702 25118 28754
rect 25170 28702 25182 28754
rect 24446 28690 24498 28702
rect 26350 28690 26402 28702
rect 29486 28754 29538 28766
rect 30158 28754 30210 28766
rect 29698 28702 29710 28754
rect 29762 28702 29774 28754
rect 29486 28690 29538 28702
rect 30158 28690 30210 28702
rect 30382 28754 30434 28766
rect 31054 28754 31106 28766
rect 30594 28702 30606 28754
rect 30658 28702 30670 28754
rect 30382 28690 30434 28702
rect 31054 28690 31106 28702
rect 32062 28754 32114 28766
rect 32846 28754 32898 28766
rect 32498 28702 32510 28754
rect 32562 28702 32574 28754
rect 32062 28690 32114 28702
rect 32846 28690 32898 28702
rect 32958 28754 33010 28766
rect 32958 28690 33010 28702
rect 33070 28754 33122 28766
rect 33070 28690 33122 28702
rect 33294 28754 33346 28766
rect 33294 28690 33346 28702
rect 33518 28754 33570 28766
rect 33518 28690 33570 28702
rect 33966 28754 34018 28766
rect 33966 28690 34018 28702
rect 34190 28754 34242 28766
rect 34190 28690 34242 28702
rect 34414 28754 34466 28766
rect 34414 28690 34466 28702
rect 34638 28754 34690 28766
rect 34638 28690 34690 28702
rect 40574 28754 40626 28766
rect 40574 28690 40626 28702
rect 46846 28754 46898 28766
rect 46846 28690 46898 28702
rect 49086 28754 49138 28766
rect 56926 28754 56978 28766
rect 51538 28702 51550 28754
rect 51602 28702 51614 28754
rect 55122 28702 55134 28754
rect 55186 28702 55198 28754
rect 49086 28690 49138 28702
rect 56926 28690 56978 28702
rect 15038 28642 15090 28654
rect 15038 28578 15090 28590
rect 20750 28642 20802 28654
rect 20750 28578 20802 28590
rect 25454 28642 25506 28654
rect 25454 28578 25506 28590
rect 25678 28642 25730 28654
rect 25678 28578 25730 28590
rect 27134 28642 27186 28654
rect 31278 28642 31330 28654
rect 29810 28590 29822 28642
rect 29874 28590 29886 28642
rect 30706 28590 30718 28642
rect 30770 28590 30782 28642
rect 27134 28578 27186 28590
rect 31278 28578 31330 28590
rect 34078 28642 34130 28654
rect 34078 28578 34130 28590
rect 38782 28642 38834 28654
rect 38782 28578 38834 28590
rect 41022 28642 41074 28654
rect 41022 28578 41074 28590
rect 44830 28642 44882 28654
rect 51326 28642 51378 28654
rect 48178 28590 48190 28642
rect 48242 28590 48254 28642
rect 44830 28578 44882 28590
rect 51326 28578 51378 28590
rect 51886 28642 51938 28654
rect 51886 28578 51938 28590
rect 52782 28642 52834 28654
rect 52782 28578 52834 28590
rect 54238 28642 54290 28654
rect 54238 28578 54290 28590
rect 57038 28642 57090 28654
rect 57038 28578 57090 28590
rect 2382 28530 2434 28542
rect 22766 28530 22818 28542
rect 8418 28478 8430 28530
rect 8482 28478 8494 28530
rect 12450 28478 12462 28530
rect 12514 28478 12526 28530
rect 21634 28478 21646 28530
rect 21698 28478 21710 28530
rect 2382 28466 2434 28478
rect 22766 28466 22818 28478
rect 24558 28530 24610 28542
rect 25902 28530 25954 28542
rect 24994 28478 25006 28530
rect 25058 28478 25070 28530
rect 24558 28466 24610 28478
rect 25902 28466 25954 28478
rect 26798 28530 26850 28542
rect 32398 28530 32450 28542
rect 31490 28478 31502 28530
rect 31554 28478 31566 28530
rect 26798 28466 26850 28478
rect 32398 28466 32450 28478
rect 45166 28530 45218 28542
rect 45166 28466 45218 28478
rect 50654 28530 50706 28542
rect 50654 28466 50706 28478
rect 25778 28366 25790 28418
rect 25842 28366 25854 28418
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 5618 28030 5630 28082
rect 5682 28079 5694 28082
rect 6290 28079 6302 28082
rect 5682 28033 6302 28079
rect 5682 28030 5694 28033
rect 6290 28030 6302 28033
rect 6354 28030 6366 28082
rect 22642 28030 22654 28082
rect 22706 28030 22718 28082
rect 33394 28030 33406 28082
rect 33458 28030 33470 28082
rect 35522 28030 35534 28082
rect 35586 28030 35598 28082
rect 38434 28030 38446 28082
rect 38498 28079 38510 28082
rect 39442 28079 39454 28082
rect 38498 28033 39454 28079
rect 38498 28030 38510 28033
rect 39442 28030 39454 28033
rect 39506 28030 39518 28082
rect 49746 28030 49758 28082
rect 49810 28030 49822 28082
rect 3838 27970 3890 27982
rect 3838 27906 3890 27918
rect 4286 27970 4338 27982
rect 4286 27906 4338 27918
rect 8990 27970 9042 27982
rect 12798 27970 12850 27982
rect 12450 27918 12462 27970
rect 12514 27918 12526 27970
rect 8990 27906 9042 27918
rect 12798 27906 12850 27918
rect 22990 27970 23042 27982
rect 22990 27906 23042 27918
rect 23438 27970 23490 27982
rect 23438 27906 23490 27918
rect 25230 27970 25282 27982
rect 25230 27906 25282 27918
rect 26686 27970 26738 27982
rect 26686 27906 26738 27918
rect 27470 27970 27522 27982
rect 27470 27906 27522 27918
rect 29710 27970 29762 27982
rect 29710 27906 29762 27918
rect 30830 27970 30882 27982
rect 30830 27906 30882 27918
rect 31838 27970 31890 27982
rect 31838 27906 31890 27918
rect 34526 27970 34578 27982
rect 34526 27906 34578 27918
rect 35198 27970 35250 27982
rect 35198 27906 35250 27918
rect 38558 27970 38610 27982
rect 38558 27906 38610 27918
rect 39454 27970 39506 27982
rect 39454 27906 39506 27918
rect 45166 27970 45218 27982
rect 45166 27906 45218 27918
rect 45614 27970 45666 27982
rect 45614 27906 45666 27918
rect 51550 27970 51602 27982
rect 51550 27906 51602 27918
rect 53118 27970 53170 27982
rect 53118 27906 53170 27918
rect 57710 27970 57762 27982
rect 57710 27906 57762 27918
rect 1822 27858 1874 27870
rect 1822 27794 1874 27806
rect 3390 27858 3442 27870
rect 3390 27794 3442 27806
rect 21646 27858 21698 27870
rect 21646 27794 21698 27806
rect 25566 27858 25618 27870
rect 25566 27794 25618 27806
rect 26126 27858 26178 27870
rect 26126 27794 26178 27806
rect 27022 27858 27074 27870
rect 27022 27794 27074 27806
rect 32174 27858 32226 27870
rect 32174 27794 32226 27806
rect 33406 27858 33458 27870
rect 33406 27794 33458 27806
rect 33518 27858 33570 27870
rect 33518 27794 33570 27806
rect 33854 27858 33906 27870
rect 33854 27794 33906 27806
rect 34190 27858 34242 27870
rect 34190 27794 34242 27806
rect 46622 27858 46674 27870
rect 46622 27794 46674 27806
rect 48302 27858 48354 27870
rect 48302 27794 48354 27806
rect 48750 27858 48802 27870
rect 48750 27794 48802 27806
rect 49422 27858 49474 27870
rect 49422 27794 49474 27806
rect 52110 27858 52162 27870
rect 54910 27858 54962 27870
rect 56926 27858 56978 27870
rect 53554 27806 53566 27858
rect 53618 27806 53630 27858
rect 56690 27806 56702 27858
rect 56754 27806 56766 27858
rect 52110 27794 52162 27806
rect 54910 27794 54962 27806
rect 56926 27794 56978 27806
rect 57150 27858 57202 27870
rect 57150 27794 57202 27806
rect 6974 27746 7026 27758
rect 6402 27694 6414 27746
rect 6466 27694 6478 27746
rect 6974 27682 7026 27694
rect 9662 27746 9714 27758
rect 17390 27746 17442 27758
rect 10210 27694 10222 27746
rect 10274 27694 10286 27746
rect 9662 27682 9714 27694
rect 17390 27682 17442 27694
rect 19518 27746 19570 27758
rect 19518 27682 19570 27694
rect 20862 27746 20914 27758
rect 22206 27746 22258 27758
rect 21746 27694 21758 27746
rect 21810 27694 21822 27746
rect 20862 27682 20914 27694
rect 22206 27682 22258 27694
rect 23998 27746 24050 27758
rect 23998 27682 24050 27694
rect 24222 27746 24274 27758
rect 24222 27682 24274 27694
rect 24446 27746 24498 27758
rect 24446 27682 24498 27694
rect 24670 27746 24722 27758
rect 24670 27682 24722 27694
rect 26350 27746 26402 27758
rect 26350 27682 26402 27694
rect 29598 27746 29650 27758
rect 29598 27682 29650 27694
rect 29822 27746 29874 27758
rect 29822 27682 29874 27694
rect 30046 27746 30098 27758
rect 30046 27682 30098 27694
rect 30270 27746 30322 27758
rect 30270 27682 30322 27694
rect 30718 27746 30770 27758
rect 30718 27682 30770 27694
rect 30942 27746 30994 27758
rect 30942 27682 30994 27694
rect 31166 27746 31218 27758
rect 31166 27682 31218 27694
rect 31390 27746 31442 27758
rect 35086 27746 35138 27758
rect 33058 27694 33070 27746
rect 33122 27694 33134 27746
rect 31390 27682 31442 27694
rect 35086 27682 35138 27694
rect 35310 27746 35362 27758
rect 35310 27682 35362 27694
rect 35646 27746 35698 27758
rect 35646 27682 35698 27694
rect 35870 27746 35922 27758
rect 35870 27682 35922 27694
rect 41806 27746 41858 27758
rect 50318 27746 50370 27758
rect 51214 27746 51266 27758
rect 52446 27746 52498 27758
rect 42130 27694 42142 27746
rect 42194 27694 42206 27746
rect 50530 27694 50542 27746
rect 50594 27694 50606 27746
rect 51538 27694 51550 27746
rect 51602 27694 51614 27746
rect 41806 27682 41858 27694
rect 50318 27682 50370 27694
rect 51214 27682 51266 27694
rect 52446 27682 52498 27694
rect 52782 27746 52834 27758
rect 52782 27682 52834 27694
rect 54238 27746 54290 27758
rect 54238 27682 54290 27694
rect 55694 27746 55746 27758
rect 57262 27746 57314 27758
rect 56578 27694 56590 27746
rect 56642 27694 56654 27746
rect 55694 27682 55746 27694
rect 57262 27682 57314 27694
rect 58158 27746 58210 27758
rect 58158 27682 58210 27694
rect 17726 27634 17778 27646
rect 39006 27634 39058 27646
rect 26002 27582 26014 27634
rect 26066 27582 26078 27634
rect 17726 27570 17778 27582
rect 39006 27570 39058 27582
rect 40350 27634 40402 27646
rect 40350 27570 40402 27582
rect 41022 27634 41074 27646
rect 41022 27570 41074 27582
rect 46062 27634 46114 27646
rect 46062 27570 46114 27582
rect 47742 27634 47794 27646
rect 47742 27570 47794 27582
rect 23886 27522 23938 27534
rect 23886 27458 23938 27470
rect 46958 27522 47010 27534
rect 46958 27458 47010 27470
rect 49086 27522 49138 27534
rect 49086 27458 49138 27470
rect 22866 27358 22878 27410
rect 22930 27358 22942 27410
rect 34514 27358 34526 27410
rect 34578 27407 34590 27410
rect 34738 27407 34750 27410
rect 34578 27361 34750 27407
rect 34578 27358 34590 27361
rect 34738 27358 34750 27361
rect 34802 27358 34814 27410
rect 42690 27358 42702 27410
rect 42754 27358 42766 27410
rect 1344 27242 58576 27276
rect 1344 27190 4478 27242
rect 4530 27190 4582 27242
rect 4634 27190 4686 27242
rect 4738 27190 35198 27242
rect 35250 27190 35302 27242
rect 35354 27190 35406 27242
rect 35458 27190 58576 27242
rect 1344 27156 58576 27190
rect 30706 27022 30718 27074
rect 30770 27022 30782 27074
rect 48850 27022 48862 27074
rect 48914 27071 48926 27074
rect 49410 27071 49422 27074
rect 48914 27025 49422 27071
rect 48914 27022 48926 27025
rect 49410 27022 49422 27025
rect 49474 27071 49486 27074
rect 50082 27071 50094 27074
rect 49474 27025 50094 27071
rect 49474 27022 49486 27025
rect 50082 27022 50094 27025
rect 50146 27022 50158 27074
rect 23886 26962 23938 26974
rect 33170 26910 33182 26962
rect 33234 26910 33246 26962
rect 23886 26898 23938 26910
rect 5742 26850 5794 26862
rect 5742 26786 5794 26798
rect 22542 26850 22594 26862
rect 22542 26786 22594 26798
rect 25118 26850 25170 26862
rect 25118 26786 25170 26798
rect 26126 26850 26178 26862
rect 26126 26786 26178 26798
rect 27022 26850 27074 26862
rect 27022 26786 27074 26798
rect 33742 26850 33794 26862
rect 37102 26850 37154 26862
rect 34066 26798 34078 26850
rect 34130 26847 34142 26850
rect 34850 26847 34862 26850
rect 34130 26801 34862 26847
rect 34130 26798 34142 26801
rect 34850 26798 34862 26801
rect 34914 26798 34926 26850
rect 33742 26786 33794 26798
rect 37102 26786 37154 26798
rect 42030 26850 42082 26862
rect 42030 26786 42082 26798
rect 15934 26738 15986 26750
rect 23774 26738 23826 26750
rect 21858 26686 21870 26738
rect 21922 26686 21934 26738
rect 15934 26674 15986 26686
rect 23774 26674 23826 26686
rect 24446 26738 24498 26750
rect 24446 26674 24498 26686
rect 24670 26738 24722 26750
rect 24670 26674 24722 26686
rect 25566 26738 25618 26750
rect 25566 26674 25618 26686
rect 25678 26738 25730 26750
rect 25678 26674 25730 26686
rect 26574 26738 26626 26750
rect 26574 26674 26626 26686
rect 29934 26738 29986 26750
rect 29934 26674 29986 26686
rect 30158 26738 30210 26750
rect 30158 26674 30210 26686
rect 30382 26738 30434 26750
rect 30382 26674 30434 26686
rect 30606 26738 30658 26750
rect 30606 26674 30658 26686
rect 31166 26738 31218 26750
rect 31166 26674 31218 26686
rect 31502 26738 31554 26750
rect 31502 26674 31554 26686
rect 31726 26738 31778 26750
rect 31726 26674 31778 26686
rect 32286 26738 32338 26750
rect 32846 26738 32898 26750
rect 39454 26738 39506 26750
rect 32498 26686 32510 26738
rect 32562 26686 32574 26738
rect 33954 26686 33966 26738
rect 34018 26735 34030 26738
rect 34962 26735 34974 26738
rect 34018 26689 34974 26735
rect 34018 26686 34030 26689
rect 34962 26686 34974 26689
rect 35026 26686 35038 26738
rect 32286 26674 32338 26686
rect 32846 26674 32898 26686
rect 39454 26674 39506 26686
rect 42702 26738 42754 26750
rect 48862 26738 48914 26750
rect 42914 26686 42926 26738
rect 42978 26686 42990 26738
rect 42702 26674 42754 26686
rect 48862 26674 48914 26686
rect 50094 26738 50146 26750
rect 50094 26674 50146 26686
rect 50766 26738 50818 26750
rect 50766 26674 50818 26686
rect 50990 26738 51042 26750
rect 50990 26674 51042 26686
rect 51214 26738 51266 26750
rect 51214 26674 51266 26686
rect 51662 26738 51714 26750
rect 51662 26674 51714 26686
rect 51886 26738 51938 26750
rect 54126 26738 54178 26750
rect 53554 26686 53566 26738
rect 53618 26686 53630 26738
rect 51886 26674 51938 26686
rect 54126 26674 54178 26686
rect 55806 26738 55858 26750
rect 57250 26686 57262 26738
rect 57314 26686 57326 26738
rect 55806 26674 55858 26686
rect 16382 26626 16434 26638
rect 16382 26562 16434 26574
rect 16942 26626 16994 26638
rect 16942 26562 16994 26574
rect 17054 26626 17106 26638
rect 17054 26562 17106 26574
rect 17726 26626 17778 26638
rect 19854 26626 19906 26638
rect 17826 26574 17838 26626
rect 17890 26574 17902 26626
rect 17726 26562 17778 26574
rect 19854 26562 19906 26574
rect 21646 26626 21698 26638
rect 21646 26562 21698 26574
rect 22094 26626 22146 26638
rect 22094 26562 22146 26574
rect 23550 26626 23602 26638
rect 23550 26562 23602 26574
rect 24222 26626 24274 26638
rect 24222 26562 24274 26574
rect 25006 26626 25058 26638
rect 25006 26562 25058 26574
rect 25230 26626 25282 26638
rect 33518 26626 33570 26638
rect 26338 26574 26350 26626
rect 26402 26574 26414 26626
rect 25230 26562 25282 26574
rect 33518 26562 33570 26574
rect 34190 26626 34242 26638
rect 34190 26562 34242 26574
rect 34302 26626 34354 26638
rect 34302 26562 34354 26574
rect 34750 26626 34802 26638
rect 34750 26562 34802 26574
rect 34974 26626 35026 26638
rect 34974 26562 35026 26574
rect 35534 26626 35586 26638
rect 35534 26562 35586 26574
rect 38446 26626 38498 26638
rect 38446 26562 38498 26574
rect 38782 26626 38834 26638
rect 38782 26562 38834 26574
rect 39118 26626 39170 26638
rect 40574 26626 40626 26638
rect 39890 26574 39902 26626
rect 39954 26574 39966 26626
rect 39118 26562 39170 26574
rect 40574 26562 40626 26574
rect 43150 26626 43202 26638
rect 43150 26562 43202 26574
rect 51438 26626 51490 26638
rect 51438 26562 51490 26574
rect 56926 26626 56978 26638
rect 56926 26562 56978 26574
rect 20750 26514 20802 26526
rect 20750 26450 20802 26462
rect 23326 26514 23378 26526
rect 23326 26450 23378 26462
rect 25902 26514 25954 26526
rect 25902 26450 25954 26462
rect 27358 26514 27410 26526
rect 27358 26450 27410 26462
rect 28590 26514 28642 26526
rect 28590 26450 28642 26462
rect 29598 26514 29650 26526
rect 29598 26450 29650 26462
rect 32062 26514 32114 26526
rect 35198 26514 35250 26526
rect 33842 26462 33854 26514
rect 33906 26462 33918 26514
rect 32062 26450 32114 26462
rect 35198 26450 35250 26462
rect 35870 26514 35922 26526
rect 35870 26450 35922 26462
rect 35982 26514 36034 26526
rect 35982 26450 36034 26462
rect 36430 26514 36482 26526
rect 36430 26450 36482 26462
rect 37550 26514 37602 26526
rect 37550 26450 37602 26462
rect 37998 26514 38050 26526
rect 37998 26450 38050 26462
rect 41246 26514 41298 26526
rect 41246 26450 41298 26462
rect 43934 26514 43986 26526
rect 43934 26450 43986 26462
rect 45502 26514 45554 26526
rect 45502 26450 45554 26462
rect 49310 26514 49362 26526
rect 49310 26450 49362 26462
rect 49758 26514 49810 26526
rect 52782 26514 52834 26526
rect 51986 26462 51998 26514
rect 52050 26462 52062 26514
rect 54338 26462 54350 26514
rect 54402 26462 54414 26514
rect 49758 26450 49810 26462
rect 52782 26450 52834 26462
rect 24322 26350 24334 26402
rect 24386 26350 24398 26402
rect 35074 26350 35086 26402
rect 35138 26350 35150 26402
rect 36978 26350 36990 26402
rect 37042 26399 37054 26402
rect 38098 26399 38110 26402
rect 37042 26353 38110 26399
rect 37042 26350 37054 26353
rect 38098 26350 38110 26353
rect 38162 26350 38174 26402
rect 42242 26350 42254 26402
rect 42306 26350 42318 26402
rect 48514 26350 48526 26402
rect 48578 26350 48590 26402
rect 50418 26350 50430 26402
rect 50482 26350 50494 26402
rect 1344 26234 58576 26268
rect 1344 26182 19838 26234
rect 19890 26182 19942 26234
rect 19994 26182 20046 26234
rect 20098 26182 50558 26234
rect 50610 26182 50662 26234
rect 50714 26182 50766 26234
rect 50818 26182 58576 26234
rect 1344 26148 58576 26182
rect 22754 26014 22766 26066
rect 22818 26014 22830 26066
rect 41122 26014 41134 26066
rect 41186 26014 41198 26066
rect 43138 26014 43150 26066
rect 43202 26014 43214 26066
rect 45826 26014 45838 26066
rect 45890 26014 45902 26066
rect 49746 26014 49758 26066
rect 49810 26063 49822 26066
rect 50978 26063 50990 26066
rect 49810 26017 50990 26063
rect 49810 26014 49822 26017
rect 50978 26014 50990 26017
rect 51042 26063 51054 26066
rect 52098 26063 52110 26066
rect 51042 26017 52110 26063
rect 51042 26014 51054 26017
rect 52098 26014 52110 26017
rect 52162 26063 52174 26066
rect 52658 26063 52670 26066
rect 52162 26017 52670 26063
rect 52162 26014 52174 26017
rect 52658 26014 52670 26017
rect 52722 26014 52734 26066
rect 16718 25954 16770 25966
rect 16718 25890 16770 25902
rect 20526 25954 20578 25966
rect 20526 25890 20578 25902
rect 25230 25954 25282 25966
rect 25230 25890 25282 25902
rect 26014 25954 26066 25966
rect 26014 25890 26066 25902
rect 26910 25954 26962 25966
rect 26910 25890 26962 25902
rect 28478 25954 28530 25966
rect 28478 25890 28530 25902
rect 29374 25954 29426 25966
rect 29374 25890 29426 25902
rect 32510 25954 32562 25966
rect 36542 25954 36594 25966
rect 33170 25902 33182 25954
rect 33234 25902 33246 25954
rect 34402 25902 34414 25954
rect 34466 25902 34478 25954
rect 32510 25890 32562 25902
rect 36542 25890 36594 25902
rect 36990 25954 37042 25966
rect 36990 25890 37042 25902
rect 49310 25954 49362 25966
rect 49310 25890 49362 25902
rect 49758 25954 49810 25966
rect 49758 25890 49810 25902
rect 51550 25954 51602 25966
rect 51550 25890 51602 25902
rect 52110 25954 52162 25966
rect 52110 25890 52162 25902
rect 53342 25954 53394 25966
rect 53342 25890 53394 25902
rect 55022 25954 55074 25966
rect 55022 25890 55074 25902
rect 55358 25954 55410 25966
rect 55358 25890 55410 25902
rect 17614 25842 17666 25854
rect 17614 25778 17666 25790
rect 18174 25842 18226 25854
rect 18174 25778 18226 25790
rect 21870 25842 21922 25854
rect 21870 25778 21922 25790
rect 23438 25842 23490 25854
rect 23438 25778 23490 25790
rect 24446 25842 24498 25854
rect 24446 25778 24498 25790
rect 25566 25842 25618 25854
rect 25566 25778 25618 25790
rect 26126 25842 26178 25854
rect 26126 25778 26178 25790
rect 27022 25842 27074 25854
rect 30830 25842 30882 25854
rect 29698 25790 29710 25842
rect 29762 25790 29774 25842
rect 27022 25778 27074 25790
rect 30830 25778 30882 25790
rect 31390 25842 31442 25854
rect 31390 25778 31442 25790
rect 31614 25842 31666 25854
rect 41246 25842 41298 25854
rect 35410 25790 35422 25842
rect 35474 25790 35486 25842
rect 31614 25778 31666 25790
rect 41246 25778 41298 25790
rect 46846 25842 46898 25854
rect 46846 25778 46898 25790
rect 54014 25842 54066 25854
rect 54014 25778 54066 25790
rect 22430 25730 22482 25742
rect 13458 25678 13470 25730
rect 13522 25678 13534 25730
rect 17938 25678 17950 25730
rect 18002 25678 18014 25730
rect 22430 25666 22482 25678
rect 23102 25730 23154 25742
rect 23102 25666 23154 25678
rect 23886 25730 23938 25742
rect 23886 25666 23938 25678
rect 25902 25730 25954 25742
rect 25902 25666 25954 25678
rect 26350 25730 26402 25742
rect 26350 25666 26402 25678
rect 26798 25730 26850 25742
rect 26798 25666 26850 25678
rect 27246 25730 27298 25742
rect 27246 25666 27298 25678
rect 30270 25730 30322 25742
rect 30270 25666 30322 25678
rect 30494 25730 30546 25742
rect 30494 25666 30546 25678
rect 30606 25730 30658 25742
rect 30606 25666 30658 25678
rect 31726 25730 31778 25742
rect 31726 25666 31778 25678
rect 31950 25730 32002 25742
rect 31950 25666 32002 25678
rect 32174 25730 32226 25742
rect 35870 25730 35922 25742
rect 33618 25678 33630 25730
rect 33682 25678 33694 25730
rect 32174 25666 32226 25678
rect 35870 25666 35922 25678
rect 36206 25730 36258 25742
rect 36206 25666 36258 25678
rect 37550 25730 37602 25742
rect 37886 25730 37938 25742
rect 37762 25678 37774 25730
rect 37826 25678 37838 25730
rect 37550 25666 37602 25678
rect 37886 25666 37938 25678
rect 38110 25730 38162 25742
rect 41022 25730 41074 25742
rect 46286 25730 46338 25742
rect 54462 25730 54514 25742
rect 39106 25678 39118 25730
rect 39170 25678 39182 25730
rect 39330 25678 39342 25730
rect 39394 25678 39406 25730
rect 39666 25678 39678 25730
rect 39730 25678 39742 25730
rect 44818 25678 44830 25730
rect 44882 25678 44894 25730
rect 46498 25678 46510 25730
rect 46562 25678 46574 25730
rect 38110 25666 38162 25678
rect 41022 25666 41074 25678
rect 46286 25666 46338 25678
rect 54462 25666 54514 25678
rect 18958 25618 19010 25630
rect 18958 25554 19010 25566
rect 20974 25618 21026 25630
rect 20974 25554 21026 25566
rect 21422 25618 21474 25630
rect 21422 25554 21474 25566
rect 24558 25618 24610 25630
rect 24558 25554 24610 25566
rect 28030 25618 28082 25630
rect 28030 25554 28082 25566
rect 28926 25618 28978 25630
rect 28926 25554 28978 25566
rect 29934 25618 29986 25630
rect 29934 25554 29986 25566
rect 31166 25618 31218 25630
rect 31166 25554 31218 25566
rect 34974 25618 35026 25630
rect 38558 25618 38610 25630
rect 35634 25566 35646 25618
rect 35698 25566 35710 25618
rect 34974 25554 35026 25566
rect 38558 25554 38610 25566
rect 50206 25618 50258 25630
rect 50206 25554 50258 25566
rect 50654 25618 50706 25630
rect 50654 25554 50706 25566
rect 51102 25618 51154 25630
rect 51102 25554 51154 25566
rect 52558 25618 52610 25630
rect 52558 25554 52610 25566
rect 55582 25618 55634 25630
rect 55582 25554 55634 25566
rect 56030 25618 56082 25630
rect 56030 25554 56082 25566
rect 56702 25618 56754 25630
rect 56702 25554 56754 25566
rect 57150 25618 57202 25630
rect 57150 25554 57202 25566
rect 57598 25618 57650 25630
rect 57598 25554 57650 25566
rect 30146 25454 30158 25506
rect 30210 25454 30222 25506
rect 49858 25454 49870 25506
rect 49922 25503 49934 25506
rect 50642 25503 50654 25506
rect 49922 25457 50654 25503
rect 49922 25454 49934 25457
rect 50642 25454 50654 25457
rect 50706 25454 50718 25506
rect 56690 25454 56702 25506
rect 56754 25503 56766 25506
rect 57586 25503 57598 25506
rect 56754 25457 57598 25503
rect 56754 25454 56766 25457
rect 57586 25454 57598 25457
rect 57650 25454 57662 25506
rect 18610 25342 18622 25394
rect 18674 25342 18686 25394
rect 50418 25342 50430 25394
rect 50482 25391 50494 25394
rect 51090 25391 51102 25394
rect 50482 25345 51102 25391
rect 50482 25342 50494 25345
rect 51090 25342 51102 25345
rect 51154 25342 51166 25394
rect 51314 25342 51326 25394
rect 51378 25391 51390 25394
rect 51650 25391 51662 25394
rect 51378 25345 51662 25391
rect 51378 25342 51390 25345
rect 51650 25342 51662 25345
rect 51714 25391 51726 25394
rect 52546 25391 52558 25394
rect 51714 25345 52558 25391
rect 51714 25342 51726 25345
rect 52546 25342 52558 25345
rect 52610 25342 52622 25394
rect 1344 25226 58576 25260
rect 1344 25174 4478 25226
rect 4530 25174 4582 25226
rect 4634 25174 4686 25226
rect 4738 25174 35198 25226
rect 35250 25174 35302 25226
rect 35354 25174 35406 25226
rect 35458 25174 58576 25226
rect 1344 25140 58576 25174
rect 24882 25006 24894 25058
rect 24946 25006 24958 25058
rect 26786 25006 26798 25058
rect 26850 25006 26862 25058
rect 47394 25006 47406 25058
rect 47458 25006 47470 25058
rect 49186 25006 49198 25058
rect 49250 25055 49262 25058
rect 50082 25055 50094 25058
rect 49250 25009 50094 25055
rect 49250 25006 49262 25009
rect 50082 25006 50094 25009
rect 50146 25006 50158 25058
rect 29934 24946 29986 24958
rect 29934 24882 29986 24894
rect 30830 24946 30882 24958
rect 30830 24882 30882 24894
rect 31390 24946 31442 24958
rect 50206 24946 50258 24958
rect 34962 24894 34974 24946
rect 35026 24894 35038 24946
rect 31390 24882 31442 24894
rect 50206 24882 50258 24894
rect 19182 24834 19234 24846
rect 16930 24782 16942 24834
rect 16994 24782 17006 24834
rect 19182 24770 19234 24782
rect 20302 24834 20354 24846
rect 20302 24770 20354 24782
rect 21646 24834 21698 24846
rect 21646 24770 21698 24782
rect 22094 24834 22146 24846
rect 27918 24834 27970 24846
rect 22866 24782 22878 24834
rect 22930 24782 22942 24834
rect 22094 24770 22146 24782
rect 27918 24770 27970 24782
rect 28590 24834 28642 24846
rect 28590 24770 28642 24782
rect 36430 24834 36482 24846
rect 36430 24770 36482 24782
rect 45726 24834 45778 24846
rect 45726 24770 45778 24782
rect 13470 24722 13522 24734
rect 13470 24658 13522 24670
rect 22430 24722 22482 24734
rect 22430 24658 22482 24670
rect 23214 24722 23266 24734
rect 23214 24658 23266 24670
rect 23326 24722 23378 24734
rect 23326 24658 23378 24670
rect 24110 24722 24162 24734
rect 26462 24722 26514 24734
rect 24658 24670 24670 24722
rect 24722 24670 24734 24722
rect 25554 24670 25566 24722
rect 25618 24670 25630 24722
rect 24110 24658 24162 24670
rect 26462 24658 26514 24670
rect 26910 24722 26962 24734
rect 26910 24658 26962 24670
rect 29374 24722 29426 24734
rect 29374 24658 29426 24670
rect 32734 24722 32786 24734
rect 32734 24658 32786 24670
rect 37998 24722 38050 24734
rect 37998 24658 38050 24670
rect 38670 24722 38722 24734
rect 53454 24722 53506 24734
rect 39778 24670 39790 24722
rect 39842 24670 39854 24722
rect 40338 24670 40350 24722
rect 40402 24670 40414 24722
rect 48402 24670 48414 24722
rect 48466 24670 48478 24722
rect 50978 24670 50990 24722
rect 51042 24670 51054 24722
rect 38670 24658 38722 24670
rect 53454 24658 53506 24670
rect 53790 24722 53842 24734
rect 53790 24658 53842 24670
rect 55246 24722 55298 24734
rect 55246 24658 55298 24670
rect 57150 24722 57202 24734
rect 57150 24658 57202 24670
rect 24334 24610 24386 24622
rect 25342 24610 25394 24622
rect 23874 24558 23886 24610
rect 23938 24558 23950 24610
rect 24546 24558 24558 24610
rect 24610 24558 24622 24610
rect 24334 24546 24386 24558
rect 25342 24546 25394 24558
rect 25790 24610 25842 24622
rect 25790 24546 25842 24558
rect 26686 24610 26738 24622
rect 26686 24546 26738 24558
rect 27470 24610 27522 24622
rect 27470 24546 27522 24558
rect 29598 24610 29650 24622
rect 29598 24546 29650 24558
rect 30270 24610 30322 24622
rect 30270 24546 30322 24558
rect 30494 24610 30546 24622
rect 30494 24546 30546 24558
rect 31054 24610 31106 24622
rect 31054 24546 31106 24558
rect 31278 24610 31330 24622
rect 31278 24546 31330 24558
rect 31838 24610 31890 24622
rect 31838 24546 31890 24558
rect 31950 24610 32002 24622
rect 38894 24610 38946 24622
rect 43598 24610 43650 24622
rect 32834 24558 32846 24610
rect 32898 24558 32910 24610
rect 33170 24558 33182 24610
rect 33234 24558 33246 24610
rect 33506 24558 33518 24610
rect 33570 24558 33582 24610
rect 42354 24558 42366 24610
rect 42418 24558 42430 24610
rect 31950 24546 32002 24558
rect 38894 24546 38946 24558
rect 43598 24546 43650 24558
rect 47854 24610 47906 24622
rect 47854 24546 47906 24558
rect 48302 24610 48354 24622
rect 48302 24546 48354 24558
rect 50654 24610 50706 24622
rect 50654 24546 50706 24558
rect 51214 24610 51266 24622
rect 51214 24546 51266 24558
rect 53118 24610 53170 24622
rect 56814 24610 56866 24622
rect 54562 24558 54574 24610
rect 54626 24558 54638 24610
rect 53118 24546 53170 24558
rect 56814 24546 56866 24558
rect 19854 24498 19906 24510
rect 19854 24434 19906 24446
rect 20750 24498 20802 24510
rect 20750 24434 20802 24446
rect 22542 24498 22594 24510
rect 22542 24434 22594 24446
rect 22878 24498 22930 24510
rect 22878 24434 22930 24446
rect 23550 24498 23602 24510
rect 23550 24434 23602 24446
rect 29822 24498 29874 24510
rect 29822 24434 29874 24446
rect 30606 24498 30658 24510
rect 35534 24498 35586 24510
rect 31490 24446 31502 24498
rect 31554 24446 31566 24498
rect 30606 24434 30658 24446
rect 35534 24434 35586 24446
rect 35982 24498 36034 24510
rect 49086 24498 49138 24510
rect 37314 24446 37326 24498
rect 37378 24446 37390 24498
rect 35982 24434 36034 24446
rect 49086 24434 49138 24446
rect 49534 24498 49586 24510
rect 49534 24434 49586 24446
rect 49982 24498 50034 24510
rect 49982 24434 50034 24446
rect 52110 24498 52162 24510
rect 52110 24434 52162 24446
rect 52782 24498 52834 24510
rect 52782 24434 52834 24446
rect 54126 24498 54178 24510
rect 54126 24434 54178 24446
rect 55918 24498 55970 24510
rect 55918 24434 55970 24446
rect 56702 24498 56754 24510
rect 56702 24434 56754 24446
rect 57822 24498 57874 24510
rect 57822 24434 57874 24446
rect 19842 24334 19854 24386
rect 19906 24383 19918 24386
rect 20738 24383 20750 24386
rect 19906 24337 20750 24383
rect 19906 24334 19918 24337
rect 20738 24334 20750 24337
rect 20802 24334 20814 24386
rect 41458 24334 41470 24386
rect 41522 24334 41534 24386
rect 49074 24334 49086 24386
rect 49138 24383 49150 24386
rect 49970 24383 49982 24386
rect 49138 24337 49982 24383
rect 49138 24334 49150 24337
rect 49970 24334 49982 24337
rect 50034 24334 50046 24386
rect 1344 24218 58576 24252
rect 1344 24166 19838 24218
rect 19890 24166 19942 24218
rect 19994 24166 20046 24218
rect 20098 24166 50558 24218
rect 50610 24166 50662 24218
rect 50714 24166 50766 24218
rect 50818 24166 58576 24218
rect 1344 24132 58576 24166
rect 26338 23998 26350 24050
rect 26402 23998 26414 24050
rect 30594 23998 30606 24050
rect 30658 23998 30670 24050
rect 49970 23998 49982 24050
rect 50034 24047 50046 24050
rect 50642 24047 50654 24050
rect 50034 24001 50654 24047
rect 50034 23998 50046 24001
rect 50642 23998 50654 24001
rect 50706 23998 50718 24050
rect 56690 23998 56702 24050
rect 56754 24047 56766 24050
rect 57474 24047 57486 24050
rect 56754 24001 57486 24047
rect 56754 23998 56766 24001
rect 57474 23998 57486 24001
rect 57538 23998 57550 24050
rect 21086 23938 21138 23950
rect 21086 23874 21138 23886
rect 21758 23938 21810 23950
rect 24558 23938 24610 23950
rect 24098 23886 24110 23938
rect 24162 23886 24174 23938
rect 21758 23874 21810 23886
rect 24558 23874 24610 23886
rect 26462 23938 26514 23950
rect 26462 23874 26514 23886
rect 27246 23938 27298 23950
rect 33742 23938 33794 23950
rect 31378 23886 31390 23938
rect 31442 23886 31454 23938
rect 27246 23874 27298 23886
rect 33742 23874 33794 23886
rect 38222 23938 38274 23950
rect 38222 23874 38274 23886
rect 44830 23938 44882 23950
rect 44830 23874 44882 23886
rect 45278 23938 45330 23950
rect 45278 23874 45330 23886
rect 47518 23938 47570 23950
rect 47518 23874 47570 23886
rect 49982 23938 50034 23950
rect 56702 23938 56754 23950
rect 55682 23886 55694 23938
rect 55746 23886 55758 23938
rect 49982 23874 50034 23886
rect 56702 23874 56754 23886
rect 19182 23826 19234 23838
rect 14578 23774 14590 23826
rect 14642 23774 14654 23826
rect 19182 23762 19234 23774
rect 19406 23826 19458 23838
rect 19406 23762 19458 23774
rect 23102 23826 23154 23838
rect 27470 23826 27522 23838
rect 25442 23774 25454 23826
rect 25506 23774 25518 23826
rect 25778 23774 25790 23826
rect 25842 23774 25854 23826
rect 23102 23762 23154 23774
rect 27470 23762 27522 23774
rect 27582 23826 27634 23838
rect 27582 23762 27634 23774
rect 34190 23826 34242 23838
rect 34190 23762 34242 23774
rect 37214 23826 37266 23838
rect 37214 23762 37266 23774
rect 37550 23826 37602 23838
rect 37550 23762 37602 23774
rect 38782 23826 38834 23838
rect 38782 23762 38834 23774
rect 40014 23826 40066 23838
rect 40014 23762 40066 23774
rect 42814 23826 42866 23838
rect 42814 23762 42866 23774
rect 45726 23826 45778 23838
rect 45726 23762 45778 23774
rect 47070 23826 47122 23838
rect 52334 23826 52386 23838
rect 47730 23774 47742 23826
rect 47794 23774 47806 23826
rect 48738 23774 48750 23826
rect 48802 23774 48814 23826
rect 53218 23774 53230 23826
rect 53282 23774 53294 23826
rect 47070 23762 47122 23774
rect 52334 23762 52386 23774
rect 17502 23714 17554 23726
rect 11666 23662 11678 23714
rect 11730 23662 11742 23714
rect 17502 23650 17554 23662
rect 18846 23714 18898 23726
rect 18846 23650 18898 23662
rect 22654 23714 22706 23726
rect 29486 23714 29538 23726
rect 23538 23662 23550 23714
rect 23602 23662 23614 23714
rect 26674 23662 26686 23714
rect 26738 23662 26750 23714
rect 22654 23650 22706 23662
rect 29486 23650 29538 23662
rect 31726 23714 31778 23726
rect 31726 23650 31778 23662
rect 31950 23714 32002 23726
rect 33070 23714 33122 23726
rect 32386 23662 32398 23714
rect 32450 23662 32462 23714
rect 31950 23650 32002 23662
rect 33070 23650 33122 23662
rect 33406 23714 33458 23726
rect 33406 23650 33458 23662
rect 37886 23714 37938 23726
rect 37886 23650 37938 23662
rect 39342 23714 39394 23726
rect 41358 23714 41410 23726
rect 41122 23662 41134 23714
rect 41186 23662 41198 23714
rect 39342 23650 39394 23662
rect 41358 23650 41410 23662
rect 41470 23714 41522 23726
rect 41470 23650 41522 23662
rect 51662 23714 51714 23726
rect 51662 23650 51714 23662
rect 51774 23714 51826 23726
rect 51774 23650 51826 23662
rect 54574 23714 54626 23726
rect 54574 23650 54626 23662
rect 54686 23714 54738 23726
rect 54686 23650 54738 23662
rect 34638 23602 34690 23614
rect 34638 23538 34690 23550
rect 36430 23602 36482 23614
rect 36430 23538 36482 23550
rect 36878 23602 36930 23614
rect 48638 23602 48690 23614
rect 41906 23550 41918 23602
rect 41970 23550 41982 23602
rect 36878 23538 36930 23550
rect 48638 23538 48690 23550
rect 48974 23602 49026 23614
rect 48974 23538 49026 23550
rect 50430 23602 50482 23614
rect 57150 23602 57202 23614
rect 51202 23550 51214 23602
rect 51266 23550 51278 23602
rect 50430 23538 50482 23550
rect 57150 23538 57202 23550
rect 57598 23602 57650 23614
rect 57598 23538 57650 23550
rect 40798 23490 40850 23502
rect 24658 23438 24670 23490
rect 24722 23438 24734 23490
rect 40798 23426 40850 23438
rect 49534 23490 49586 23502
rect 57138 23438 57150 23490
rect 57202 23487 57214 23490
rect 57586 23487 57598 23490
rect 57202 23441 57598 23487
rect 57202 23438 57214 23441
rect 57586 23438 57598 23441
rect 57650 23438 57662 23490
rect 49534 23426 49586 23438
rect 46610 23326 46622 23378
rect 46674 23326 46686 23378
rect 1344 23210 58576 23244
rect 1344 23158 4478 23210
rect 4530 23158 4582 23210
rect 4634 23158 4686 23210
rect 4738 23158 35198 23210
rect 35250 23158 35302 23210
rect 35354 23158 35406 23210
rect 35458 23158 58576 23210
rect 1344 23124 58576 23158
rect 16594 22990 16606 23042
rect 16658 22990 16670 23042
rect 25890 22990 25902 23042
rect 25954 22990 25966 23042
rect 37314 22990 37326 23042
rect 37378 22990 37390 23042
rect 40114 22990 40126 23042
rect 40178 22990 40190 23042
rect 41346 22990 41358 23042
rect 41410 23039 41422 23042
rect 41794 23039 41806 23042
rect 41410 22993 41806 23039
rect 41410 22990 41422 22993
rect 41794 22990 41806 22993
rect 41858 22990 41870 23042
rect 50866 22990 50878 23042
rect 50930 22990 50942 23042
rect 41906 22927 41918 22930
rect 41249 22881 41918 22927
rect 17614 22818 17666 22830
rect 17614 22754 17666 22766
rect 19406 22818 19458 22830
rect 19406 22754 19458 22766
rect 19854 22818 19906 22830
rect 19854 22754 19906 22766
rect 20302 22818 20354 22830
rect 20302 22754 20354 22766
rect 20750 22818 20802 22830
rect 20750 22754 20802 22766
rect 21646 22818 21698 22830
rect 21646 22754 21698 22766
rect 22094 22818 22146 22830
rect 22094 22754 22146 22766
rect 22542 22818 22594 22830
rect 22542 22754 22594 22766
rect 33966 22818 34018 22830
rect 33966 22754 34018 22766
rect 36206 22818 36258 22830
rect 36206 22754 36258 22766
rect 38894 22818 38946 22830
rect 40898 22766 40910 22818
rect 40962 22815 40974 22818
rect 41249 22815 41295 22881
rect 41906 22878 41918 22881
rect 41970 22878 41982 22930
rect 40962 22769 41295 22815
rect 41358 22818 41410 22830
rect 40962 22766 40974 22769
rect 38894 22754 38946 22766
rect 41358 22754 41410 22766
rect 41806 22818 41858 22830
rect 41806 22754 41858 22766
rect 42254 22818 42306 22830
rect 42254 22754 42306 22766
rect 42702 22818 42754 22830
rect 42702 22754 42754 22766
rect 52782 22818 52834 22830
rect 52782 22754 52834 22766
rect 58158 22818 58210 22830
rect 58158 22754 58210 22766
rect 25678 22706 25730 22718
rect 15138 22654 15150 22706
rect 15202 22654 15214 22706
rect 24658 22654 24670 22706
rect 24722 22654 24734 22706
rect 25678 22642 25730 22654
rect 26350 22706 26402 22718
rect 29262 22706 29314 22718
rect 30718 22706 30770 22718
rect 26786 22654 26798 22706
rect 26850 22654 26862 22706
rect 29474 22654 29486 22706
rect 29538 22703 29550 22706
rect 30034 22703 30046 22706
rect 29538 22657 30046 22703
rect 29538 22654 29550 22657
rect 30034 22654 30046 22657
rect 30098 22654 30110 22706
rect 26350 22642 26402 22654
rect 29262 22642 29314 22654
rect 30718 22642 30770 22654
rect 30942 22706 30994 22718
rect 30942 22642 30994 22654
rect 31278 22706 31330 22718
rect 31278 22642 31330 22654
rect 31390 22706 31442 22718
rect 31390 22642 31442 22654
rect 37886 22706 37938 22718
rect 37886 22642 37938 22654
rect 40462 22706 40514 22718
rect 40462 22642 40514 22654
rect 40686 22706 40738 22718
rect 40686 22642 40738 22654
rect 40910 22706 40962 22718
rect 40910 22642 40962 22654
rect 46622 22706 46674 22718
rect 46622 22642 46674 22654
rect 46958 22706 47010 22718
rect 46958 22642 47010 22654
rect 47630 22706 47682 22718
rect 47630 22642 47682 22654
rect 48190 22706 48242 22718
rect 54014 22706 54066 22718
rect 51538 22654 51550 22706
rect 51602 22654 51614 22706
rect 48190 22642 48242 22654
rect 54014 22642 54066 22654
rect 55806 22706 55858 22718
rect 55806 22642 55858 22654
rect 57486 22706 57538 22718
rect 57486 22642 57538 22654
rect 57710 22706 57762 22718
rect 57710 22642 57762 22654
rect 24334 22594 24386 22606
rect 26910 22594 26962 22606
rect 25554 22542 25566 22594
rect 25618 22542 25630 22594
rect 24334 22530 24386 22542
rect 26910 22530 26962 22542
rect 27806 22594 27858 22606
rect 27806 22530 27858 22542
rect 29598 22594 29650 22606
rect 29598 22530 29650 22542
rect 29822 22594 29874 22606
rect 29822 22530 29874 22542
rect 30494 22594 30546 22606
rect 30494 22530 30546 22542
rect 31166 22594 31218 22606
rect 31166 22530 31218 22542
rect 32622 22594 32674 22606
rect 32622 22530 32674 22542
rect 39118 22594 39170 22606
rect 39118 22530 39170 22542
rect 40238 22594 40290 22606
rect 40238 22530 40290 22542
rect 47294 22594 47346 22606
rect 47294 22530 47346 22542
rect 48750 22594 48802 22606
rect 48750 22530 48802 22542
rect 51326 22594 51378 22606
rect 51326 22530 51378 22542
rect 51886 22594 51938 22606
rect 51886 22530 51938 22542
rect 53678 22594 53730 22606
rect 53678 22530 53730 22542
rect 54350 22594 54402 22606
rect 57262 22594 57314 22606
rect 55122 22542 55134 22594
rect 55186 22542 55198 22594
rect 54350 22530 54402 22542
rect 57262 22530 57314 22542
rect 22990 22482 23042 22494
rect 22990 22418 23042 22430
rect 27470 22482 27522 22494
rect 27470 22418 27522 22430
rect 28590 22482 28642 22494
rect 31950 22482 32002 22494
rect 30146 22430 30158 22482
rect 30210 22430 30222 22482
rect 28590 22418 28642 22430
rect 31950 22418 32002 22430
rect 32286 22482 32338 22494
rect 32286 22418 32338 22430
rect 33070 22482 33122 22494
rect 33070 22418 33122 22430
rect 33518 22482 33570 22494
rect 33518 22418 33570 22430
rect 35758 22482 35810 22494
rect 35758 22418 35810 22430
rect 49422 22482 49474 22494
rect 49422 22418 49474 22430
rect 50206 22482 50258 22494
rect 50206 22418 50258 22430
rect 50654 22482 50706 22494
rect 50654 22418 50706 22430
rect 53230 22482 53282 22494
rect 53230 22418 53282 22430
rect 54686 22482 54738 22494
rect 54686 22418 54738 22430
rect 56478 22482 56530 22494
rect 57138 22430 57150 22482
rect 57202 22430 57214 22482
rect 56478 22418 56530 22430
rect 29922 22318 29934 22370
rect 29986 22318 29998 22370
rect 1344 22202 58576 22236
rect 1344 22150 19838 22202
rect 19890 22150 19942 22202
rect 19994 22150 20046 22202
rect 20098 22150 50558 22202
rect 50610 22150 50662 22202
rect 50714 22150 50766 22202
rect 50818 22150 58576 22202
rect 1344 22116 58576 22150
rect 26114 21982 26126 22034
rect 26178 21982 26190 22034
rect 39566 21922 39618 21934
rect 23762 21870 23774 21922
rect 23826 21870 23838 21922
rect 30594 21870 30606 21922
rect 30658 21870 30670 21922
rect 39566 21858 39618 21870
rect 41022 21922 41074 21934
rect 41022 21858 41074 21870
rect 41470 21922 41522 21934
rect 41470 21858 41522 21870
rect 41918 21922 41970 21934
rect 41918 21858 41970 21870
rect 47294 21922 47346 21934
rect 47294 21858 47346 21870
rect 53006 21922 53058 21934
rect 53006 21858 53058 21870
rect 21534 21810 21586 21822
rect 25342 21810 25394 21822
rect 23202 21758 23214 21810
rect 23266 21758 23278 21810
rect 21534 21746 21586 21758
rect 25342 21746 25394 21758
rect 25678 21810 25730 21822
rect 25678 21746 25730 21758
rect 27358 21810 27410 21822
rect 27358 21746 27410 21758
rect 28702 21810 28754 21822
rect 31726 21810 31778 21822
rect 29922 21758 29934 21810
rect 29986 21758 29998 21810
rect 30930 21758 30942 21810
rect 30994 21807 31006 21810
rect 31154 21807 31166 21810
rect 30994 21761 31166 21807
rect 30994 21758 31006 21761
rect 31154 21758 31166 21761
rect 31218 21758 31230 21810
rect 28702 21746 28754 21758
rect 31726 21746 31778 21758
rect 34414 21810 34466 21822
rect 34414 21746 34466 21758
rect 34974 21810 35026 21822
rect 34974 21746 35026 21758
rect 35646 21810 35698 21822
rect 35646 21746 35698 21758
rect 35870 21810 35922 21822
rect 35870 21746 35922 21758
rect 38222 21810 38274 21822
rect 38222 21746 38274 21758
rect 42366 21810 42418 21822
rect 42366 21746 42418 21758
rect 43038 21810 43090 21822
rect 43038 21746 43090 21758
rect 43598 21810 43650 21822
rect 43598 21746 43650 21758
rect 45054 21810 45106 21822
rect 45054 21746 45106 21758
rect 49422 21810 49474 21822
rect 49422 21746 49474 21758
rect 52222 21810 52274 21822
rect 52222 21746 52274 21758
rect 55246 21810 55298 21822
rect 55246 21746 55298 21758
rect 56702 21810 56754 21822
rect 56702 21746 56754 21758
rect 19854 21698 19906 21710
rect 19854 21634 19906 21646
rect 20190 21698 20242 21710
rect 20190 21634 20242 21646
rect 22654 21698 22706 21710
rect 22654 21634 22706 21646
rect 25118 21698 25170 21710
rect 25118 21634 25170 21646
rect 26462 21698 26514 21710
rect 30270 21698 30322 21710
rect 32286 21698 32338 21710
rect 29138 21646 29150 21698
rect 29202 21646 29214 21698
rect 31938 21646 31950 21698
rect 32002 21646 32014 21698
rect 26462 21634 26514 21646
rect 30270 21634 30322 21646
rect 32286 21634 32338 21646
rect 44606 21698 44658 21710
rect 44606 21634 44658 21646
rect 45166 21698 45218 21710
rect 45166 21634 45218 21646
rect 45390 21698 45442 21710
rect 45390 21634 45442 21646
rect 48862 21698 48914 21710
rect 48862 21634 48914 21646
rect 49758 21698 49810 21710
rect 49758 21634 49810 21646
rect 50094 21698 50146 21710
rect 50094 21634 50146 21646
rect 50430 21698 50482 21710
rect 50430 21634 50482 21646
rect 50990 21698 51042 21710
rect 50990 21634 51042 21646
rect 51550 21698 51602 21710
rect 51550 21634 51602 21646
rect 54126 21698 54178 21710
rect 54126 21634 54178 21646
rect 24670 21586 24722 21598
rect 24670 21522 24722 21534
rect 25454 21586 25506 21598
rect 25454 21522 25506 21534
rect 26910 21586 26962 21598
rect 26910 21522 26962 21534
rect 34078 21586 34130 21598
rect 34078 21522 34130 21534
rect 36654 21586 36706 21598
rect 36654 21522 36706 21534
rect 37102 21586 37154 21598
rect 37102 21522 37154 21534
rect 37550 21586 37602 21598
rect 37550 21522 37602 21534
rect 38670 21586 38722 21598
rect 38670 21522 38722 21534
rect 39118 21586 39170 21598
rect 39118 21522 39170 21534
rect 40014 21586 40066 21598
rect 40014 21522 40066 21534
rect 44158 21586 44210 21598
rect 44158 21522 44210 21534
rect 47854 21586 47906 21598
rect 55470 21586 55522 21598
rect 53442 21534 53454 21586
rect 53506 21534 53518 21586
rect 47854 21522 47906 21534
rect 55470 21522 55522 21534
rect 56030 21586 56082 21598
rect 56030 21522 56082 21534
rect 57150 21586 57202 21598
rect 57150 21522 57202 21534
rect 36206 21474 36258 21486
rect 42702 21474 42754 21486
rect 36642 21422 36654 21474
rect 36706 21471 36718 21474
rect 36866 21471 36878 21474
rect 36706 21425 36878 21471
rect 36706 21422 36718 21425
rect 36866 21422 36878 21425
rect 36930 21471 36942 21474
rect 37538 21471 37550 21474
rect 36930 21425 37550 21471
rect 36930 21422 36942 21425
rect 37538 21422 37550 21425
rect 37602 21422 37614 21474
rect 38210 21422 38222 21474
rect 38274 21471 38286 21474
rect 38658 21471 38670 21474
rect 38274 21425 38670 21471
rect 38274 21422 38286 21425
rect 38658 21422 38670 21425
rect 38722 21422 38734 21474
rect 36206 21410 36258 21422
rect 42702 21410 42754 21422
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 22530 20974 22542 21026
rect 22594 20974 22606 21026
rect 22754 20974 22766 21026
rect 22818 21023 22830 21026
rect 24210 21023 24222 21026
rect 22818 20977 24222 21023
rect 22818 20974 22830 20977
rect 24210 20974 24222 20977
rect 24274 20974 24286 21026
rect 35186 20974 35198 21026
rect 35250 20974 35262 21026
rect 49186 20974 49198 21026
rect 49250 20974 49262 21026
rect 51874 20974 51886 21026
rect 51938 20974 51950 21026
rect 30258 20862 30270 20914
rect 30322 20862 30334 20914
rect 32498 20862 32510 20914
rect 32562 20862 32574 20914
rect 22878 20802 22930 20814
rect 22878 20738 22930 20750
rect 23326 20802 23378 20814
rect 23326 20738 23378 20750
rect 23774 20802 23826 20814
rect 23774 20738 23826 20750
rect 24222 20802 24274 20814
rect 24222 20738 24274 20750
rect 24670 20802 24722 20814
rect 24670 20738 24722 20750
rect 26350 20802 26402 20814
rect 26350 20738 26402 20750
rect 26798 20802 26850 20814
rect 26798 20738 26850 20750
rect 27694 20802 27746 20814
rect 27694 20738 27746 20750
rect 28142 20802 28194 20814
rect 28142 20738 28194 20750
rect 33966 20802 34018 20814
rect 33966 20738 34018 20750
rect 34974 20802 35026 20814
rect 34974 20738 35026 20750
rect 36318 20802 36370 20814
rect 36318 20738 36370 20750
rect 37214 20802 37266 20814
rect 37214 20738 37266 20750
rect 44942 20802 44994 20814
rect 44942 20738 44994 20750
rect 45502 20802 45554 20814
rect 45502 20738 45554 20750
rect 49086 20802 49138 20814
rect 49086 20738 49138 20750
rect 54910 20802 54962 20814
rect 54910 20738 54962 20750
rect 55358 20802 55410 20814
rect 55358 20738 55410 20750
rect 56254 20802 56306 20814
rect 56254 20738 56306 20750
rect 30606 20690 30658 20702
rect 18498 20638 18510 20690
rect 18562 20638 18574 20690
rect 30606 20626 30658 20638
rect 30830 20690 30882 20702
rect 30830 20626 30882 20638
rect 31166 20690 31218 20702
rect 31166 20626 31218 20638
rect 31390 20690 31442 20702
rect 31390 20626 31442 20638
rect 31614 20690 31666 20702
rect 31614 20626 31666 20638
rect 31950 20690 32002 20702
rect 31950 20626 32002 20638
rect 32846 20690 32898 20702
rect 32846 20626 32898 20638
rect 33070 20690 33122 20702
rect 33070 20626 33122 20638
rect 37550 20690 37602 20702
rect 37550 20626 37602 20638
rect 40350 20690 40402 20702
rect 40350 20626 40402 20638
rect 41470 20690 41522 20702
rect 41470 20626 41522 20638
rect 41582 20690 41634 20702
rect 41582 20626 41634 20638
rect 46398 20690 46450 20702
rect 46398 20626 46450 20638
rect 48078 20690 48130 20702
rect 48078 20626 48130 20638
rect 48638 20690 48690 20702
rect 48638 20626 48690 20638
rect 49534 20690 49586 20702
rect 50542 20690 50594 20702
rect 53566 20690 53618 20702
rect 49746 20638 49758 20690
rect 49810 20638 49822 20690
rect 50866 20638 50878 20690
rect 50930 20638 50942 20690
rect 49534 20626 49586 20638
rect 50542 20626 50594 20638
rect 53566 20626 53618 20638
rect 53790 20690 53842 20702
rect 53790 20626 53842 20638
rect 55806 20690 55858 20702
rect 55806 20626 55858 20638
rect 21422 20578 21474 20590
rect 21422 20514 21474 20526
rect 21534 20578 21586 20590
rect 21534 20514 21586 20526
rect 22094 20578 22146 20590
rect 22094 20514 22146 20526
rect 31838 20578 31890 20590
rect 31838 20514 31890 20526
rect 32062 20578 32114 20590
rect 32062 20514 32114 20526
rect 35646 20578 35698 20590
rect 35646 20514 35698 20526
rect 36206 20578 36258 20590
rect 42702 20578 42754 20590
rect 41794 20526 41806 20578
rect 41858 20526 41870 20578
rect 36206 20514 36258 20526
rect 42702 20514 42754 20526
rect 45950 20578 46002 20590
rect 45950 20514 46002 20526
rect 47630 20578 47682 20590
rect 47630 20514 47682 20526
rect 19742 20466 19794 20478
rect 19742 20402 19794 20414
rect 20302 20466 20354 20478
rect 20302 20402 20354 20414
rect 20750 20466 20802 20478
rect 20750 20402 20802 20414
rect 25454 20466 25506 20478
rect 25454 20402 25506 20414
rect 25902 20466 25954 20478
rect 27246 20466 27298 20478
rect 27122 20414 27134 20466
rect 27186 20414 27198 20466
rect 25902 20402 25954 20414
rect 25442 20302 25454 20354
rect 25506 20351 25518 20354
rect 25890 20351 25902 20354
rect 25506 20305 25902 20351
rect 25506 20302 25518 20305
rect 25890 20302 25902 20305
rect 25954 20351 25966 20354
rect 26898 20351 26910 20354
rect 25954 20305 26910 20351
rect 25954 20302 25966 20305
rect 26898 20302 26910 20305
rect 26962 20351 26974 20354
rect 27137 20351 27183 20414
rect 27246 20402 27298 20414
rect 28590 20466 28642 20478
rect 28590 20402 28642 20414
rect 29486 20466 29538 20478
rect 29486 20402 29538 20414
rect 29934 20466 29986 20478
rect 29934 20402 29986 20414
rect 33518 20466 33570 20478
rect 33518 20402 33570 20414
rect 38334 20466 38386 20478
rect 38334 20402 38386 20414
rect 40798 20466 40850 20478
rect 40798 20402 40850 20414
rect 43710 20466 43762 20478
rect 43710 20402 43762 20414
rect 46846 20466 46898 20478
rect 46846 20402 46898 20414
rect 54238 20466 54290 20478
rect 54238 20402 54290 20414
rect 26962 20305 27183 20351
rect 26962 20302 26974 20305
rect 27346 20302 27358 20354
rect 27410 20351 27422 20354
rect 27682 20351 27694 20354
rect 27410 20305 27694 20351
rect 27410 20302 27422 20305
rect 27682 20302 27694 20305
rect 27746 20302 27758 20354
rect 1344 20186 58576 20220
rect 1344 20134 19838 20186
rect 19890 20134 19942 20186
rect 19994 20134 20046 20186
rect 20098 20134 50558 20186
rect 50610 20134 50662 20186
rect 50714 20134 50766 20186
rect 50818 20134 58576 20186
rect 1344 20100 58576 20134
rect 51426 19966 51438 20018
rect 51490 19966 51502 20018
rect 20638 19906 20690 19918
rect 20638 19842 20690 19854
rect 24110 19906 24162 19918
rect 24110 19842 24162 19854
rect 25342 19906 25394 19918
rect 25342 19842 25394 19854
rect 26014 19906 26066 19918
rect 26014 19842 26066 19854
rect 28926 19906 28978 19918
rect 33070 19906 33122 19918
rect 30706 19854 30718 19906
rect 30770 19854 30782 19906
rect 28926 19842 28978 19854
rect 33070 19842 33122 19854
rect 33742 19906 33794 19918
rect 33742 19842 33794 19854
rect 34414 19906 34466 19918
rect 34414 19842 34466 19854
rect 35198 19906 35250 19918
rect 35198 19842 35250 19854
rect 46622 19906 46674 19918
rect 46622 19842 46674 19854
rect 48302 19906 48354 19918
rect 48302 19842 48354 19854
rect 52894 19906 52946 19918
rect 52894 19842 52946 19854
rect 22766 19794 22818 19806
rect 21074 19742 21086 19794
rect 21138 19742 21150 19794
rect 22766 19730 22818 19742
rect 29598 19794 29650 19806
rect 29598 19730 29650 19742
rect 30830 19794 30882 19806
rect 30830 19730 30882 19742
rect 33406 19794 33458 19806
rect 33406 19730 33458 19742
rect 34078 19794 34130 19806
rect 34078 19730 34130 19742
rect 34750 19794 34802 19806
rect 40910 19794 40962 19806
rect 38658 19742 38670 19794
rect 38722 19742 38734 19794
rect 34750 19730 34802 19742
rect 40910 19730 40962 19742
rect 41358 19794 41410 19806
rect 52222 19794 52274 19806
rect 43474 19742 43486 19794
rect 43538 19742 43550 19794
rect 49074 19742 49086 19794
rect 49138 19742 49150 19794
rect 41358 19730 41410 19742
rect 52222 19730 52274 19742
rect 54686 19794 54738 19806
rect 54686 19730 54738 19742
rect 20974 19682 21026 19694
rect 17714 19630 17726 19682
rect 17778 19630 17790 19682
rect 20974 19618 21026 19630
rect 29262 19682 29314 19694
rect 29262 19618 29314 19630
rect 29710 19682 29762 19694
rect 29710 19618 29762 19630
rect 30606 19682 30658 19694
rect 30606 19618 30658 19630
rect 31054 19682 31106 19694
rect 31054 19618 31106 19630
rect 32286 19682 32338 19694
rect 32286 19618 32338 19630
rect 35982 19682 36034 19694
rect 35982 19618 36034 19630
rect 36318 19682 36370 19694
rect 51886 19682 51938 19694
rect 39106 19630 39118 19682
rect 39170 19630 39182 19682
rect 47730 19630 47742 19682
rect 47794 19630 47806 19682
rect 49970 19630 49982 19682
rect 50034 19630 50046 19682
rect 51538 19630 51550 19682
rect 51602 19630 51614 19682
rect 36318 19618 36370 19630
rect 51886 19618 51938 19630
rect 52558 19682 52610 19694
rect 52558 19618 52610 19630
rect 53454 19682 53506 19694
rect 53454 19618 53506 19630
rect 54014 19682 54066 19694
rect 54014 19618 54066 19630
rect 24558 19570 24610 19582
rect 24558 19506 24610 19518
rect 26462 19570 26514 19582
rect 26462 19506 26514 19518
rect 26910 19570 26962 19582
rect 26910 19506 26962 19518
rect 27582 19570 27634 19582
rect 27582 19506 27634 19518
rect 28030 19570 28082 19582
rect 28030 19506 28082 19518
rect 28478 19570 28530 19582
rect 28478 19506 28530 19518
rect 45614 19570 45666 19582
rect 45614 19506 45666 19518
rect 46062 19570 46114 19582
rect 55470 19570 55522 19582
rect 47618 19518 47630 19570
rect 47682 19518 47694 19570
rect 46062 19506 46114 19518
rect 55470 19506 55522 19518
rect 19294 19458 19346 19470
rect 44270 19458 44322 19470
rect 28242 19406 28254 19458
rect 28306 19455 28318 19458
rect 28914 19455 28926 19458
rect 28306 19409 28926 19455
rect 28306 19406 28318 19409
rect 28914 19406 28926 19409
rect 28978 19406 28990 19458
rect 40226 19406 40238 19458
rect 40290 19406 40302 19458
rect 50082 19406 50094 19458
rect 50146 19406 50158 19458
rect 19294 19394 19346 19406
rect 44270 19394 44322 19406
rect 22754 19294 22766 19346
rect 22818 19294 22830 19346
rect 1344 19178 58576 19212
rect 1344 19126 4478 19178
rect 4530 19126 4582 19178
rect 4634 19126 4686 19178
rect 4738 19126 35198 19178
rect 35250 19126 35302 19178
rect 35354 19126 35406 19178
rect 35458 19126 58576 19178
rect 1344 19092 58576 19126
rect 27682 18958 27694 19010
rect 27746 19007 27758 19010
rect 28130 19007 28142 19010
rect 27746 18961 28142 19007
rect 27746 18958 27758 18961
rect 28130 18958 28142 18961
rect 28194 18958 28206 19010
rect 38882 18958 38894 19010
rect 38946 19007 38958 19010
rect 40226 19007 40238 19010
rect 38946 18961 40238 19007
rect 38946 18958 38958 18961
rect 40226 18958 40238 18961
rect 40290 18958 40302 19010
rect 54674 18958 54686 19010
rect 54738 18958 54750 19010
rect 26686 18898 26738 18910
rect 33182 18898 33234 18910
rect 26898 18846 26910 18898
rect 26962 18895 26974 18898
rect 27234 18895 27246 18898
rect 26962 18849 27246 18895
rect 26962 18846 26974 18849
rect 27234 18846 27246 18849
rect 27298 18895 27310 18898
rect 28242 18895 28254 18898
rect 27298 18849 28254 18895
rect 27298 18846 27310 18849
rect 28242 18846 28254 18849
rect 28306 18846 28318 18898
rect 35970 18846 35982 18898
rect 36034 18895 36046 18898
rect 36418 18895 36430 18898
rect 36034 18849 36430 18895
rect 36034 18846 36046 18849
rect 36418 18846 36430 18849
rect 36482 18846 36494 18898
rect 39218 18846 39230 18898
rect 39282 18895 39294 18898
rect 40002 18895 40014 18898
rect 39282 18849 40014 18895
rect 39282 18846 39294 18849
rect 40002 18846 40014 18849
rect 40066 18846 40078 18898
rect 52770 18846 52782 18898
rect 52834 18895 52846 18898
rect 53218 18895 53230 18898
rect 52834 18849 53230 18895
rect 52834 18846 52846 18849
rect 53218 18846 53230 18849
rect 53282 18846 53294 18898
rect 26686 18834 26738 18846
rect 33182 18834 33234 18846
rect 20414 18786 20466 18798
rect 20414 18722 20466 18734
rect 21870 18786 21922 18798
rect 21870 18722 21922 18734
rect 22318 18786 22370 18798
rect 22318 18722 22370 18734
rect 27246 18786 27298 18798
rect 27246 18722 27298 18734
rect 27694 18786 27746 18798
rect 27694 18722 27746 18734
rect 28142 18786 28194 18798
rect 28142 18722 28194 18734
rect 28590 18786 28642 18798
rect 28590 18722 28642 18734
rect 35534 18786 35586 18798
rect 17502 18674 17554 18686
rect 17502 18610 17554 18622
rect 18286 18674 18338 18686
rect 18286 18610 18338 18622
rect 18958 18674 19010 18686
rect 23214 18674 23266 18686
rect 19730 18622 19742 18674
rect 19794 18622 19806 18674
rect 18958 18610 19010 18622
rect 23214 18610 23266 18622
rect 23886 18674 23938 18686
rect 31378 18678 31390 18730
rect 31442 18678 31454 18730
rect 35534 18722 35586 18734
rect 36430 18786 36482 18798
rect 36430 18722 36482 18734
rect 40238 18786 40290 18798
rect 40238 18722 40290 18734
rect 46398 18786 46450 18798
rect 46398 18722 46450 18734
rect 49982 18786 50034 18798
rect 52782 18786 52834 18798
rect 51874 18734 51886 18786
rect 51938 18734 51950 18786
rect 49982 18722 50034 18734
rect 52782 18722 52834 18734
rect 53230 18786 53282 18798
rect 53230 18722 53282 18734
rect 53678 18786 53730 18798
rect 53678 18722 53730 18734
rect 23886 18610 23938 18622
rect 31726 18674 31778 18686
rect 31726 18610 31778 18622
rect 32846 18674 32898 18686
rect 32846 18610 32898 18622
rect 35982 18674 36034 18686
rect 35982 18610 36034 18622
rect 39342 18674 39394 18686
rect 39342 18610 39394 18622
rect 40574 18674 40626 18686
rect 40574 18610 40626 18622
rect 41246 18674 41298 18686
rect 41246 18610 41298 18622
rect 41582 18674 41634 18686
rect 41582 18610 41634 18622
rect 42702 18674 42754 18686
rect 42702 18610 42754 18622
rect 48862 18674 48914 18686
rect 48862 18610 48914 18622
rect 50094 18674 50146 18686
rect 57026 18622 57038 18674
rect 57090 18622 57102 18674
rect 50094 18610 50146 18622
rect 16606 18562 16658 18574
rect 16606 18498 16658 18510
rect 17726 18562 17778 18574
rect 17726 18498 17778 18510
rect 18062 18562 18114 18574
rect 18062 18498 18114 18510
rect 21422 18562 21474 18574
rect 21422 18498 21474 18510
rect 22878 18562 22930 18574
rect 22878 18498 22930 18510
rect 23550 18562 23602 18574
rect 23550 18498 23602 18510
rect 24446 18562 24498 18574
rect 24446 18498 24498 18510
rect 25006 18562 25058 18574
rect 25006 18498 25058 18510
rect 26350 18562 26402 18574
rect 26350 18498 26402 18510
rect 29598 18562 29650 18574
rect 29598 18498 29650 18510
rect 31278 18562 31330 18574
rect 31278 18498 31330 18510
rect 33854 18562 33906 18574
rect 33854 18498 33906 18510
rect 34750 18562 34802 18574
rect 34750 18498 34802 18510
rect 38558 18562 38610 18574
rect 38558 18498 38610 18510
rect 38894 18562 38946 18574
rect 38894 18498 38946 18510
rect 39790 18562 39842 18574
rect 39790 18498 39842 18510
rect 40910 18562 40962 18574
rect 40910 18498 40962 18510
rect 42142 18562 42194 18574
rect 42142 18498 42194 18510
rect 43374 18562 43426 18574
rect 43374 18498 43426 18510
rect 47070 18562 47122 18574
rect 47070 18498 47122 18510
rect 47966 18562 48018 18574
rect 49422 18562 49474 18574
rect 48738 18559 48750 18562
rect 47966 18498 48018 18510
rect 48641 18513 48750 18559
rect 17054 18450 17106 18462
rect 17054 18386 17106 18398
rect 19182 18450 19234 18462
rect 19182 18386 19234 18398
rect 19518 18450 19570 18462
rect 19518 18386 19570 18398
rect 20078 18450 20130 18462
rect 20078 18386 20130 18398
rect 25678 18450 25730 18462
rect 25678 18386 25730 18398
rect 35086 18450 35138 18462
rect 35086 18386 35138 18398
rect 45278 18450 45330 18462
rect 45278 18386 45330 18398
rect 45726 18450 45778 18462
rect 45726 18386 45778 18398
rect 47518 18450 47570 18462
rect 47518 18386 47570 18398
rect 48414 18450 48466 18462
rect 48414 18386 48466 18398
rect 18722 18286 18734 18338
rect 18786 18286 18798 18338
rect 47506 18286 47518 18338
rect 47570 18335 47582 18338
rect 48066 18335 48078 18338
rect 47570 18289 48078 18335
rect 47570 18286 47582 18289
rect 48066 18286 48078 18289
rect 48130 18335 48142 18338
rect 48641 18335 48687 18513
rect 48738 18510 48750 18513
rect 48802 18510 48814 18562
rect 49422 18498 49474 18510
rect 50654 18562 50706 18574
rect 50866 18510 50878 18562
rect 50930 18510 50942 18562
rect 50654 18498 50706 18510
rect 49086 18450 49138 18462
rect 49086 18386 49138 18398
rect 48130 18289 48687 18335
rect 48130 18286 48142 18289
rect 1344 18170 58576 18204
rect 1344 18118 19838 18170
rect 19890 18118 19942 18170
rect 19994 18118 20046 18170
rect 20098 18118 50558 18170
rect 50610 18118 50662 18170
rect 50714 18118 50766 18170
rect 50818 18118 58576 18170
rect 1344 18084 58576 18118
rect 54002 17950 54014 18002
rect 54066 17950 54078 18002
rect 20750 17890 20802 17902
rect 20750 17826 20802 17838
rect 22542 17890 22594 17902
rect 22542 17826 22594 17838
rect 25790 17890 25842 17902
rect 25790 17826 25842 17838
rect 26350 17890 26402 17902
rect 26350 17826 26402 17838
rect 27358 17890 27410 17902
rect 27358 17826 27410 17838
rect 29822 17890 29874 17902
rect 29822 17826 29874 17838
rect 35310 17890 35362 17902
rect 35310 17826 35362 17838
rect 38110 17890 38162 17902
rect 38110 17826 38162 17838
rect 43486 17890 43538 17902
rect 43486 17826 43538 17838
rect 48190 17890 48242 17902
rect 48190 17826 48242 17838
rect 50542 17890 50594 17902
rect 50542 17826 50594 17838
rect 53118 17890 53170 17902
rect 53118 17826 53170 17838
rect 19742 17778 19794 17790
rect 19742 17714 19794 17726
rect 28030 17778 28082 17790
rect 28030 17714 28082 17726
rect 30494 17778 30546 17790
rect 30494 17714 30546 17726
rect 30830 17778 30882 17790
rect 30830 17714 30882 17726
rect 38446 17778 38498 17790
rect 38446 17714 38498 17726
rect 41358 17778 41410 17790
rect 41358 17714 41410 17726
rect 42926 17778 42978 17790
rect 42926 17714 42978 17726
rect 46846 17778 46898 17790
rect 46846 17714 46898 17726
rect 47406 17778 47458 17790
rect 47406 17714 47458 17726
rect 47854 17778 47906 17790
rect 47854 17714 47906 17726
rect 48078 17778 48130 17790
rect 48078 17714 48130 17726
rect 49534 17778 49586 17790
rect 49534 17714 49586 17726
rect 51102 17778 51154 17790
rect 51102 17714 51154 17726
rect 52334 17778 52386 17790
rect 52334 17714 52386 17726
rect 17614 17666 17666 17678
rect 17614 17602 17666 17614
rect 18286 17666 18338 17678
rect 18286 17602 18338 17614
rect 20078 17666 20130 17678
rect 20078 17602 20130 17614
rect 20414 17666 20466 17678
rect 20414 17602 20466 17614
rect 21310 17666 21362 17678
rect 21310 17602 21362 17614
rect 21870 17666 21922 17678
rect 21870 17602 21922 17614
rect 28702 17666 28754 17678
rect 28702 17602 28754 17614
rect 29262 17666 29314 17678
rect 29262 17602 29314 17614
rect 30158 17666 30210 17678
rect 30158 17602 30210 17614
rect 43934 17666 43986 17678
rect 49870 17666 49922 17678
rect 45938 17614 45950 17666
rect 46002 17614 46014 17666
rect 47618 17614 47630 17666
rect 47682 17614 47694 17666
rect 43934 17602 43986 17614
rect 49870 17602 49922 17614
rect 50206 17666 50258 17678
rect 50206 17602 50258 17614
rect 51662 17666 51714 17678
rect 51662 17602 51714 17614
rect 53342 17666 53394 17678
rect 53342 17602 53394 17614
rect 16830 17554 16882 17566
rect 16830 17490 16882 17502
rect 18734 17554 18786 17566
rect 18734 17490 18786 17502
rect 24222 17554 24274 17566
rect 24222 17490 24274 17502
rect 24670 17554 24722 17566
rect 24670 17490 24722 17502
rect 25342 17554 25394 17566
rect 25342 17490 25394 17502
rect 26910 17554 26962 17566
rect 26910 17490 26962 17502
rect 37662 17554 37714 17566
rect 48862 17554 48914 17566
rect 42130 17502 42142 17554
rect 42194 17502 42206 17554
rect 37662 17490 37714 17502
rect 48862 17490 48914 17502
rect 44706 17390 44718 17442
rect 44770 17390 44782 17442
rect 40450 17278 40462 17330
rect 40514 17278 40526 17330
rect 1344 17162 58576 17196
rect 1344 17110 4478 17162
rect 4530 17110 4582 17162
rect 4634 17110 4686 17162
rect 4738 17110 35198 17162
rect 35250 17110 35302 17162
rect 35354 17110 35406 17162
rect 35458 17110 58576 17162
rect 1344 17076 58576 17110
rect 37650 16830 37662 16882
rect 37714 16879 37726 16882
rect 37714 16833 38831 16879
rect 37714 16830 37726 16833
rect 20750 16770 20802 16782
rect 20750 16706 20802 16718
rect 27246 16770 27298 16782
rect 38670 16770 38722 16782
rect 34962 16718 34974 16770
rect 35026 16718 35038 16770
rect 38785 16767 38831 16833
rect 55582 16770 55634 16782
rect 38994 16767 39006 16770
rect 38785 16721 39006 16767
rect 38994 16718 39006 16721
rect 39058 16718 39070 16770
rect 50194 16718 50206 16770
rect 50258 16718 50270 16770
rect 27246 16706 27298 16718
rect 38670 16706 38722 16718
rect 55582 16706 55634 16718
rect 21422 16658 21474 16670
rect 15026 16606 15038 16658
rect 15090 16606 15102 16658
rect 21422 16594 21474 16606
rect 21870 16658 21922 16670
rect 21870 16594 21922 16606
rect 22206 16658 22258 16670
rect 22206 16594 22258 16606
rect 23774 16658 23826 16670
rect 23774 16594 23826 16606
rect 24446 16658 24498 16670
rect 24446 16594 24498 16606
rect 25006 16658 25058 16670
rect 25006 16594 25058 16606
rect 29822 16658 29874 16670
rect 29822 16594 29874 16606
rect 30158 16658 30210 16670
rect 30158 16594 30210 16606
rect 31278 16658 31330 16670
rect 31278 16594 31330 16606
rect 37326 16658 37378 16670
rect 37326 16594 37378 16606
rect 38222 16658 38274 16670
rect 38222 16594 38274 16606
rect 40350 16658 40402 16670
rect 40350 16594 40402 16606
rect 43038 16658 43090 16670
rect 43038 16594 43090 16606
rect 46286 16658 46338 16670
rect 46286 16594 46338 16606
rect 46734 16658 46786 16670
rect 52558 16658 52610 16670
rect 48962 16606 48974 16658
rect 49026 16606 49038 16658
rect 49746 16606 49758 16658
rect 49810 16606 49822 16658
rect 50754 16606 50766 16658
rect 50818 16606 50830 16658
rect 46734 16594 46786 16606
rect 52558 16594 52610 16606
rect 23438 16546 23490 16558
rect 23438 16482 23490 16494
rect 24110 16546 24162 16558
rect 24110 16482 24162 16494
rect 25566 16546 25618 16558
rect 25566 16482 25618 16494
rect 27582 16546 27634 16558
rect 27582 16482 27634 16494
rect 28590 16546 28642 16558
rect 28590 16482 28642 16494
rect 29150 16546 29202 16558
rect 29150 16482 29202 16494
rect 29486 16546 29538 16558
rect 31950 16546 32002 16558
rect 30594 16494 30606 16546
rect 30658 16494 30670 16546
rect 29486 16482 29538 16494
rect 31950 16482 32002 16494
rect 33854 16546 33906 16558
rect 33854 16482 33906 16494
rect 37774 16546 37826 16558
rect 37774 16482 37826 16494
rect 39230 16546 39282 16558
rect 39230 16482 39282 16494
rect 39454 16546 39506 16558
rect 39454 16482 39506 16494
rect 39902 16546 39954 16558
rect 39902 16482 39954 16494
rect 43374 16546 43426 16558
rect 43374 16482 43426 16494
rect 44830 16546 44882 16558
rect 52894 16546 52946 16558
rect 47170 16494 47182 16546
rect 47234 16494 47246 16546
rect 51202 16494 51214 16546
rect 51266 16494 51278 16546
rect 44830 16482 44882 16494
rect 52894 16482 52946 16494
rect 53566 16546 53618 16558
rect 53566 16482 53618 16494
rect 54238 16546 54290 16558
rect 54238 16482 54290 16494
rect 20190 16434 20242 16446
rect 22990 16434 23042 16446
rect 21746 16382 21758 16434
rect 21810 16382 21822 16434
rect 20190 16370 20242 16382
rect 22990 16370 23042 16382
rect 26238 16434 26290 16446
rect 26238 16370 26290 16382
rect 28254 16434 28306 16446
rect 28254 16370 28306 16382
rect 33518 16434 33570 16446
rect 33518 16370 33570 16382
rect 46062 16434 46114 16446
rect 46062 16370 46114 16382
rect 52558 16434 52610 16446
rect 54562 16382 54574 16434
rect 54626 16382 54638 16434
rect 54898 16382 54910 16434
rect 54962 16382 54974 16434
rect 52558 16370 52610 16382
rect 19170 16270 19182 16322
rect 19234 16270 19246 16322
rect 44146 16270 44158 16322
rect 44210 16270 44222 16322
rect 1344 16154 58576 16188
rect 1344 16102 19838 16154
rect 19890 16102 19942 16154
rect 19994 16102 20046 16154
rect 20098 16102 50558 16154
rect 50610 16102 50662 16154
rect 50714 16102 50766 16154
rect 50818 16102 58576 16154
rect 1344 16068 58576 16102
rect 25554 15934 25566 15986
rect 25618 15934 25630 15986
rect 40786 15934 40798 15986
rect 40850 15983 40862 15986
rect 41122 15983 41134 15986
rect 40850 15937 41134 15983
rect 40850 15934 40862 15937
rect 41122 15934 41134 15937
rect 41186 15934 41198 15986
rect 51762 15934 51774 15986
rect 51826 15934 51838 15986
rect 52770 15934 52782 15986
rect 52834 15934 52846 15986
rect 19966 15874 20018 15886
rect 19966 15810 20018 15822
rect 22654 15874 22706 15886
rect 37774 15874 37826 15886
rect 24098 15822 24110 15874
rect 24162 15822 24174 15874
rect 28466 15822 28478 15874
rect 28530 15822 28542 15874
rect 22654 15810 22706 15822
rect 37774 15810 37826 15822
rect 40350 15874 40402 15886
rect 40350 15810 40402 15822
rect 41022 15874 41074 15886
rect 41022 15810 41074 15822
rect 42366 15874 42418 15886
rect 42366 15810 42418 15822
rect 44158 15874 44210 15886
rect 47518 15874 47570 15886
rect 44930 15822 44942 15874
rect 44994 15822 45006 15874
rect 44158 15810 44210 15822
rect 47518 15810 47570 15822
rect 49310 15874 49362 15886
rect 49310 15810 49362 15822
rect 50766 15874 50818 15886
rect 50766 15810 50818 15822
rect 51214 15874 51266 15886
rect 51214 15810 51266 15822
rect 19294 15762 19346 15774
rect 19294 15698 19346 15710
rect 20526 15762 20578 15774
rect 20526 15698 20578 15710
rect 21086 15762 21138 15774
rect 21086 15698 21138 15710
rect 21758 15762 21810 15774
rect 21758 15698 21810 15710
rect 25342 15762 25394 15774
rect 25342 15698 25394 15710
rect 25454 15762 25506 15774
rect 28814 15762 28866 15774
rect 25778 15710 25790 15762
rect 25842 15710 25854 15762
rect 25454 15698 25506 15710
rect 28814 15698 28866 15710
rect 30046 15762 30098 15774
rect 30046 15698 30098 15710
rect 31950 15762 32002 15774
rect 31950 15698 32002 15710
rect 33070 15762 33122 15774
rect 33070 15698 33122 15710
rect 36206 15762 36258 15774
rect 36206 15698 36258 15710
rect 36766 15762 36818 15774
rect 36766 15698 36818 15710
rect 37438 15762 37490 15774
rect 37438 15698 37490 15710
rect 39566 15762 39618 15774
rect 39566 15698 39618 15710
rect 41358 15762 41410 15774
rect 41358 15698 41410 15710
rect 42030 15762 42082 15774
rect 42030 15698 42082 15710
rect 43486 15762 43538 15774
rect 43486 15698 43538 15710
rect 46174 15762 46226 15774
rect 46174 15698 46226 15710
rect 18958 15650 19010 15662
rect 18958 15586 19010 15598
rect 19630 15650 19682 15662
rect 19630 15586 19682 15598
rect 22990 15650 23042 15662
rect 22990 15586 23042 15598
rect 23438 15650 23490 15662
rect 23438 15586 23490 15598
rect 23886 15650 23938 15662
rect 28254 15650 28306 15662
rect 24322 15598 24334 15650
rect 24386 15598 24398 15650
rect 26002 15598 26014 15650
rect 26066 15598 26078 15650
rect 23886 15586 23938 15598
rect 28254 15586 28306 15598
rect 31278 15650 31330 15662
rect 31278 15586 31330 15598
rect 37102 15650 37154 15662
rect 37102 15586 37154 15598
rect 38334 15650 38386 15662
rect 38334 15586 38386 15598
rect 38894 15650 38946 15662
rect 38894 15586 38946 15598
rect 41694 15650 41746 15662
rect 41694 15586 41746 15598
rect 42926 15650 42978 15662
rect 42926 15586 42978 15598
rect 47070 15650 47122 15662
rect 47070 15586 47122 15598
rect 47966 15650 48018 15662
rect 47966 15586 48018 15598
rect 49758 15650 49810 15662
rect 49758 15586 49810 15598
rect 52558 15650 52610 15662
rect 54238 15650 54290 15662
rect 53330 15598 53342 15650
rect 53394 15598 53406 15650
rect 52558 15586 52610 15598
rect 54238 15586 54290 15598
rect 18174 15538 18226 15550
rect 18174 15474 18226 15486
rect 18622 15538 18674 15550
rect 18622 15474 18674 15486
rect 26798 15538 26850 15550
rect 26798 15474 26850 15486
rect 29038 15538 29090 15550
rect 29038 15474 29090 15486
rect 48862 15538 48914 15550
rect 48862 15474 48914 15486
rect 50206 15538 50258 15550
rect 50206 15474 50258 15486
rect 18162 15374 18174 15426
rect 18226 15423 18238 15426
rect 18610 15423 18622 15426
rect 18226 15377 18622 15423
rect 18226 15374 18238 15377
rect 18610 15374 18622 15377
rect 18674 15374 18686 15426
rect 1344 15146 58576 15180
rect 1344 15094 4478 15146
rect 4530 15094 4582 15146
rect 4634 15094 4686 15146
rect 4738 15094 35198 15146
rect 35250 15094 35302 15146
rect 35354 15094 35406 15146
rect 35458 15094 58576 15146
rect 1344 15060 58576 15094
rect 19058 14926 19070 14978
rect 19122 14926 19134 14978
rect 30482 14926 30494 14978
rect 30546 14926 30558 14978
rect 45378 14814 45390 14866
rect 45442 14863 45454 14866
rect 46274 14863 46286 14866
rect 45442 14817 46286 14863
rect 45442 14814 45454 14817
rect 46274 14814 46286 14817
rect 46338 14863 46350 14866
rect 46946 14863 46958 14866
rect 46338 14817 46958 14863
rect 46338 14814 46350 14817
rect 46946 14814 46958 14817
rect 47010 14814 47022 14866
rect 20302 14754 20354 14766
rect 29374 14754 29426 14766
rect 22642 14702 22654 14754
rect 22706 14702 22718 14754
rect 20302 14690 20354 14702
rect 29374 14690 29426 14702
rect 29710 14754 29762 14766
rect 29710 14690 29762 14702
rect 32734 14754 32786 14766
rect 38222 14754 38274 14766
rect 36418 14702 36430 14754
rect 36482 14702 36494 14754
rect 32734 14690 32786 14702
rect 38222 14690 38274 14702
rect 40238 14754 40290 14766
rect 40238 14690 40290 14702
rect 41694 14754 41746 14766
rect 41694 14690 41746 14702
rect 42366 14754 42418 14766
rect 42366 14690 42418 14702
rect 43822 14754 43874 14766
rect 43822 14690 43874 14702
rect 45838 14754 45890 14766
rect 45838 14690 45890 14702
rect 46286 14754 46338 14766
rect 46286 14690 46338 14702
rect 47182 14754 47234 14766
rect 47182 14690 47234 14702
rect 47630 14754 47682 14766
rect 47630 14690 47682 14702
rect 49310 14754 49362 14766
rect 49310 14690 49362 14702
rect 50542 14754 50594 14766
rect 50542 14690 50594 14702
rect 50990 14754 51042 14766
rect 50990 14690 51042 14702
rect 51662 14754 51714 14766
rect 51662 14690 51714 14702
rect 52110 14754 52162 14766
rect 52110 14690 52162 14702
rect 52782 14754 52834 14766
rect 52782 14690 52834 14702
rect 22430 14642 22482 14654
rect 18610 14590 18622 14642
rect 18674 14590 18686 14642
rect 22430 14578 22482 14590
rect 26014 14642 26066 14654
rect 26014 14578 26066 14590
rect 26910 14642 26962 14654
rect 26910 14578 26962 14590
rect 30158 14642 30210 14654
rect 30158 14578 30210 14590
rect 30382 14642 30434 14654
rect 30382 14578 30434 14590
rect 30606 14642 30658 14654
rect 30606 14578 30658 14590
rect 30830 14642 30882 14654
rect 30830 14578 30882 14590
rect 33182 14642 33234 14654
rect 37886 14642 37938 14654
rect 45390 14642 45442 14654
rect 34738 14590 34750 14642
rect 34802 14590 34814 14642
rect 37090 14590 37102 14642
rect 37154 14590 37166 14642
rect 39666 14590 39678 14642
rect 39730 14590 39742 14642
rect 33182 14578 33234 14590
rect 37886 14578 37938 14590
rect 45390 14578 45442 14590
rect 53230 14642 53282 14654
rect 53230 14578 53282 14590
rect 24446 14530 24498 14542
rect 22082 14478 22094 14530
rect 22146 14478 22158 14530
rect 23986 14478 23998 14530
rect 24050 14478 24062 14530
rect 24446 14466 24498 14478
rect 26238 14530 26290 14542
rect 26238 14466 26290 14478
rect 34078 14530 34130 14542
rect 34078 14466 34130 14478
rect 35646 14530 35698 14542
rect 35646 14466 35698 14478
rect 39006 14530 39058 14542
rect 39006 14466 39058 14478
rect 40574 14530 40626 14542
rect 40574 14466 40626 14478
rect 44942 14530 44994 14542
rect 44942 14466 44994 14478
rect 19854 14418 19906 14430
rect 19854 14354 19906 14366
rect 20750 14418 20802 14430
rect 20750 14354 20802 14366
rect 27694 14418 27746 14430
rect 27694 14354 27746 14366
rect 28142 14418 28194 14430
rect 28142 14354 28194 14366
rect 28590 14418 28642 14430
rect 28590 14354 28642 14366
rect 32286 14418 32338 14430
rect 32286 14354 32338 14366
rect 38558 14418 38610 14430
rect 38558 14354 38610 14366
rect 44270 14418 44322 14430
rect 44270 14354 44322 14366
rect 46734 14418 46786 14430
rect 46734 14354 46786 14366
rect 50094 14418 50146 14430
rect 50094 14354 50146 14366
rect 26562 14254 26574 14306
rect 26626 14254 26638 14306
rect 27682 14254 27694 14306
rect 27746 14303 27758 14306
rect 28242 14303 28254 14306
rect 27746 14257 28254 14303
rect 27746 14254 27758 14257
rect 28242 14254 28254 14257
rect 28306 14254 28318 14306
rect 33506 14254 33518 14306
rect 33570 14254 33582 14306
rect 46722 14254 46734 14306
rect 46786 14303 46798 14306
rect 47170 14303 47182 14306
rect 46786 14257 47182 14303
rect 46786 14254 46798 14257
rect 47170 14254 47182 14257
rect 47234 14254 47246 14306
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 21970 13918 21982 13970
rect 22034 13918 22046 13970
rect 26114 13918 26126 13970
rect 26178 13967 26190 13970
rect 27682 13967 27694 13970
rect 26178 13921 27694 13967
rect 26178 13918 26190 13921
rect 27682 13918 27694 13921
rect 27746 13918 27758 13970
rect 37986 13918 37998 13970
rect 38050 13918 38062 13970
rect 20974 13858 21026 13870
rect 20974 13794 21026 13806
rect 21422 13858 21474 13870
rect 21422 13794 21474 13806
rect 22766 13858 22818 13870
rect 22766 13794 22818 13806
rect 23214 13858 23266 13870
rect 23214 13794 23266 13806
rect 24222 13858 24274 13870
rect 24222 13794 24274 13806
rect 24670 13858 24722 13870
rect 24670 13794 24722 13806
rect 25454 13858 25506 13870
rect 25454 13794 25506 13806
rect 25902 13858 25954 13870
rect 25902 13794 25954 13806
rect 26350 13858 26402 13870
rect 26350 13794 26402 13806
rect 26798 13858 26850 13870
rect 26798 13794 26850 13806
rect 27694 13858 27746 13870
rect 27694 13794 27746 13806
rect 29262 13858 29314 13870
rect 29262 13794 29314 13806
rect 29710 13858 29762 13870
rect 29710 13794 29762 13806
rect 32062 13858 32114 13870
rect 32062 13794 32114 13806
rect 39006 13858 39058 13870
rect 39006 13794 39058 13806
rect 40350 13858 40402 13870
rect 40350 13794 40402 13806
rect 41358 13858 41410 13870
rect 41358 13794 41410 13806
rect 42702 13858 42754 13870
rect 42702 13794 42754 13806
rect 45614 13858 45666 13870
rect 45614 13794 45666 13806
rect 51214 13858 51266 13870
rect 51214 13794 51266 13806
rect 22318 13746 22370 13758
rect 22318 13682 22370 13694
rect 41022 13746 41074 13758
rect 41022 13682 41074 13694
rect 41694 13746 41746 13758
rect 41694 13682 41746 13694
rect 42030 13746 42082 13758
rect 42030 13682 42082 13694
rect 42366 13746 42418 13758
rect 44494 13746 44546 13758
rect 43138 13694 43150 13746
rect 43202 13694 43214 13746
rect 42366 13682 42418 13694
rect 44494 13682 44546 13694
rect 47182 13746 47234 13758
rect 47182 13682 47234 13694
rect 27246 13634 27298 13646
rect 27246 13570 27298 13582
rect 28142 13634 28194 13646
rect 28142 13570 28194 13582
rect 32510 13634 32562 13646
rect 32510 13570 32562 13582
rect 33742 13634 33794 13646
rect 34862 13634 34914 13646
rect 33954 13582 33966 13634
rect 34018 13582 34030 13634
rect 33742 13570 33794 13582
rect 34862 13570 34914 13582
rect 43822 13634 43874 13646
rect 43822 13570 43874 13582
rect 46398 13634 46450 13646
rect 46398 13570 46450 13582
rect 19406 13522 19458 13534
rect 19406 13458 19458 13470
rect 20526 13522 20578 13534
rect 20526 13458 20578 13470
rect 28814 13522 28866 13534
rect 28814 13458 28866 13470
rect 30158 13522 30210 13534
rect 30158 13458 30210 13470
rect 33182 13522 33234 13534
rect 33182 13458 33234 13470
rect 34302 13522 34354 13534
rect 34302 13458 34354 13470
rect 37326 13522 37378 13534
rect 37326 13458 37378 13470
rect 38558 13522 38610 13534
rect 47842 13470 47854 13522
rect 47906 13470 47918 13522
rect 38558 13458 38610 13470
rect 1344 13130 58576 13164
rect 1344 13078 4478 13130
rect 4530 13078 4582 13130
rect 4634 13078 4686 13130
rect 4738 13078 35198 13130
rect 35250 13078 35302 13130
rect 35354 13078 35406 13130
rect 35458 13078 58576 13130
rect 1344 13044 58576 13078
rect 26898 12910 26910 12962
rect 26962 12959 26974 12962
rect 27346 12959 27358 12962
rect 26962 12913 27358 12959
rect 26962 12910 26974 12913
rect 27346 12910 27358 12913
rect 27410 12959 27422 12962
rect 27794 12959 27806 12962
rect 27410 12913 27806 12959
rect 27410 12910 27422 12913
rect 27794 12910 27806 12913
rect 27858 12910 27870 12962
rect 31938 12910 31950 12962
rect 32002 12910 32014 12962
rect 33618 12910 33630 12962
rect 33682 12959 33694 12962
rect 34290 12959 34302 12962
rect 33682 12913 34302 12959
rect 33682 12910 33694 12913
rect 34290 12910 34302 12913
rect 34354 12910 34366 12962
rect 44034 12910 44046 12962
rect 44098 12910 44110 12962
rect 26574 12850 26626 12862
rect 37874 12798 37886 12850
rect 37938 12847 37950 12850
rect 38546 12847 38558 12850
rect 37938 12801 38558 12847
rect 37938 12798 37950 12801
rect 38546 12798 38558 12801
rect 38610 12847 38622 12850
rect 39106 12847 39118 12850
rect 38610 12801 39118 12847
rect 38610 12798 38622 12801
rect 39106 12798 39118 12801
rect 39170 12798 39182 12850
rect 47730 12798 47742 12850
rect 47794 12798 47806 12850
rect 26574 12786 26626 12798
rect 21422 12738 21474 12750
rect 21422 12674 21474 12686
rect 21870 12738 21922 12750
rect 21870 12674 21922 12686
rect 23326 12738 23378 12750
rect 27358 12738 27410 12750
rect 24210 12686 24222 12738
rect 24274 12686 24286 12738
rect 23326 12674 23378 12686
rect 27358 12674 27410 12686
rect 27806 12738 27858 12750
rect 27806 12674 27858 12686
rect 33630 12738 33682 12750
rect 33630 12674 33682 12686
rect 34078 12738 34130 12750
rect 34078 12674 34130 12686
rect 34526 12738 34578 12750
rect 34526 12674 34578 12686
rect 36430 12738 36482 12750
rect 36430 12674 36482 12686
rect 38110 12738 38162 12750
rect 38110 12674 38162 12686
rect 38558 12738 38610 12750
rect 38558 12674 38610 12686
rect 17614 12626 17666 12638
rect 37102 12626 37154 12638
rect 25778 12574 25790 12626
rect 25842 12574 25854 12626
rect 32722 12574 32734 12626
rect 32786 12574 32798 12626
rect 17614 12562 17666 12574
rect 37102 12562 37154 12574
rect 39006 12626 39058 12638
rect 39006 12562 39058 12574
rect 39342 12626 39394 12638
rect 39342 12562 39394 12574
rect 39678 12626 39730 12638
rect 39678 12562 39730 12574
rect 39902 12626 39954 12638
rect 39902 12562 39954 12574
rect 40574 12626 40626 12638
rect 40574 12562 40626 12574
rect 49982 12626 50034 12638
rect 49982 12562 50034 12574
rect 18286 12514 18338 12526
rect 18286 12450 18338 12462
rect 20638 12514 20690 12526
rect 20638 12450 20690 12462
rect 24334 12514 24386 12526
rect 24334 12450 24386 12462
rect 32398 12514 32450 12526
rect 32398 12450 32450 12462
rect 32846 12514 32898 12526
rect 32846 12450 32898 12462
rect 42926 12514 42978 12526
rect 42926 12450 42978 12462
rect 44942 12514 44994 12526
rect 48178 12462 48190 12514
rect 48242 12462 48254 12514
rect 44942 12450 44994 12462
rect 23774 12402 23826 12414
rect 23774 12338 23826 12350
rect 1344 12122 58576 12156
rect 1344 12070 19838 12122
rect 19890 12070 19942 12122
rect 19994 12070 20046 12122
rect 20098 12070 50558 12122
rect 50610 12070 50662 12122
rect 50714 12070 50766 12122
rect 50818 12070 58576 12122
rect 1344 12036 58576 12070
rect 22082 11902 22094 11954
rect 22146 11951 22158 11954
rect 22866 11951 22878 11954
rect 22146 11905 22878 11951
rect 22146 11902 22158 11905
rect 22866 11902 22878 11905
rect 22930 11902 22942 11954
rect 22878 11842 22930 11854
rect 22878 11778 22930 11790
rect 43598 11842 43650 11854
rect 46274 11790 46286 11842
rect 46338 11790 46350 11842
rect 43598 11778 43650 11790
rect 22430 11730 22482 11742
rect 17938 11678 17950 11730
rect 18002 11678 18014 11730
rect 19842 11678 19854 11730
rect 19906 11678 19918 11730
rect 22430 11666 22482 11678
rect 23102 11730 23154 11742
rect 23102 11666 23154 11678
rect 23998 11730 24050 11742
rect 23998 11666 24050 11678
rect 25342 11730 25394 11742
rect 25342 11666 25394 11678
rect 27806 11730 27858 11742
rect 27806 11666 27858 11678
rect 33406 11730 33458 11742
rect 33406 11666 33458 11678
rect 34638 11730 34690 11742
rect 34638 11666 34690 11678
rect 35870 11730 35922 11742
rect 35870 11666 35922 11678
rect 44046 11730 44098 11742
rect 44046 11666 44098 11678
rect 44494 11730 44546 11742
rect 44494 11666 44546 11678
rect 46622 11730 46674 11742
rect 46622 11666 46674 11678
rect 17502 11618 17554 11630
rect 17502 11554 17554 11566
rect 23550 11618 23602 11630
rect 23550 11554 23602 11566
rect 24222 11618 24274 11630
rect 24222 11554 24274 11566
rect 30942 11618 30994 11630
rect 30942 11554 30994 11566
rect 32286 11618 32338 11630
rect 32286 11554 32338 11566
rect 33070 11618 33122 11630
rect 33070 11554 33122 11566
rect 33742 11618 33794 11630
rect 33742 11554 33794 11566
rect 34078 11618 34130 11630
rect 34078 11554 34130 11566
rect 35198 11618 35250 11630
rect 35198 11554 35250 11566
rect 48078 11618 48130 11630
rect 48078 11554 48130 11566
rect 21982 11506 22034 11518
rect 21074 11454 21086 11506
rect 21138 11454 21150 11506
rect 21982 11442 22034 11454
rect 26350 11506 26402 11518
rect 28254 11506 28306 11518
rect 27234 11454 27246 11506
rect 27298 11503 27310 11506
rect 27298 11457 27743 11503
rect 27298 11454 27310 11457
rect 26350 11442 26402 11454
rect 27697 11391 27743 11457
rect 28254 11442 28306 11454
rect 28702 11506 28754 11518
rect 28702 11442 28754 11454
rect 29150 11506 29202 11518
rect 29150 11442 29202 11454
rect 30606 11506 30658 11518
rect 30606 11442 30658 11454
rect 38782 11506 38834 11518
rect 38782 11442 38834 11454
rect 39230 11506 39282 11518
rect 39230 11442 39282 11454
rect 28130 11391 28142 11394
rect 27697 11345 28142 11391
rect 28130 11342 28142 11345
rect 28194 11342 28206 11394
rect 28690 11230 28702 11282
rect 28754 11279 28766 11282
rect 29250 11279 29262 11282
rect 28754 11233 29262 11279
rect 28754 11230 28766 11233
rect 29250 11230 29262 11233
rect 29314 11230 29326 11282
rect 1344 11114 58576 11148
rect 1344 11062 4478 11114
rect 4530 11062 4582 11114
rect 4634 11062 4686 11114
rect 4738 11062 35198 11114
rect 35250 11062 35302 11114
rect 35354 11062 35406 11114
rect 35458 11062 58576 11114
rect 1344 11028 58576 11062
rect 27794 10894 27806 10946
rect 27858 10894 27870 10946
rect 42590 10834 42642 10846
rect 42590 10770 42642 10782
rect 20638 10722 20690 10734
rect 28142 10722 28194 10734
rect 25890 10670 25902 10722
rect 25954 10670 25966 10722
rect 20638 10658 20690 10670
rect 28142 10658 28194 10670
rect 38782 10722 38834 10734
rect 38782 10658 38834 10670
rect 19070 10610 19122 10622
rect 16930 10558 16942 10610
rect 16994 10558 17006 10610
rect 19070 10546 19122 10558
rect 21646 10610 21698 10622
rect 21646 10546 21698 10558
rect 21982 10610 22034 10622
rect 21982 10546 22034 10558
rect 22318 10610 22370 10622
rect 22318 10546 22370 10558
rect 23438 10610 23490 10622
rect 23438 10546 23490 10558
rect 25006 10610 25058 10622
rect 38334 10610 38386 10622
rect 27122 10558 27134 10610
rect 27186 10558 27198 10610
rect 30594 10558 30606 10610
rect 30658 10558 30670 10610
rect 25006 10546 25058 10558
rect 38334 10546 38386 10558
rect 39678 10610 39730 10622
rect 39678 10546 39730 10558
rect 40126 10610 40178 10622
rect 40126 10546 40178 10558
rect 16382 10498 16434 10510
rect 16382 10434 16434 10446
rect 21310 10498 21362 10510
rect 21310 10434 21362 10446
rect 22878 10498 22930 10510
rect 22878 10434 22930 10446
rect 26910 10498 26962 10510
rect 26910 10434 26962 10446
rect 27358 10498 27410 10510
rect 27358 10434 27410 10446
rect 29374 10498 29426 10510
rect 29374 10434 29426 10446
rect 29710 10498 29762 10510
rect 29710 10434 29762 10446
rect 30046 10498 30098 10510
rect 30046 10434 30098 10446
rect 33070 10498 33122 10510
rect 33070 10434 33122 10446
rect 19742 10386 19794 10398
rect 19742 10322 19794 10334
rect 24110 10386 24162 10398
rect 24110 10322 24162 10334
rect 28590 10386 28642 10398
rect 28590 10322 28642 10334
rect 34526 10386 34578 10398
rect 34526 10322 34578 10334
rect 39230 10386 39282 10398
rect 39230 10322 39282 10334
rect 42142 10386 42194 10398
rect 42142 10322 42194 10334
rect 1344 10106 58576 10140
rect 1344 10054 19838 10106
rect 19890 10054 19942 10106
rect 19994 10054 20046 10106
rect 20098 10054 50558 10106
rect 50610 10054 50662 10106
rect 50714 10054 50766 10106
rect 50818 10054 58576 10106
rect 1344 10020 58576 10054
rect 22418 9886 22430 9938
rect 22482 9886 22494 9938
rect 23202 9886 23214 9938
rect 23266 9935 23278 9938
rect 24658 9935 24670 9938
rect 23266 9889 24670 9935
rect 23266 9886 23278 9889
rect 24658 9886 24670 9889
rect 24722 9886 24734 9938
rect 23214 9826 23266 9838
rect 23214 9762 23266 9774
rect 24222 9826 24274 9838
rect 24222 9762 24274 9774
rect 24670 9826 24722 9838
rect 24670 9762 24722 9774
rect 25342 9826 25394 9838
rect 25342 9762 25394 9774
rect 26910 9826 26962 9838
rect 26910 9762 26962 9774
rect 41918 9826 41970 9838
rect 41918 9762 41970 9774
rect 20190 9714 20242 9726
rect 20190 9650 20242 9662
rect 25902 9714 25954 9726
rect 25902 9650 25954 9662
rect 26238 9714 26290 9726
rect 26238 9650 26290 9662
rect 27470 9714 27522 9726
rect 27470 9650 27522 9662
rect 28702 9714 28754 9726
rect 28702 9650 28754 9662
rect 29598 9714 29650 9726
rect 29598 9650 29650 9662
rect 42478 9714 42530 9726
rect 42478 9650 42530 9662
rect 43038 9714 43090 9726
rect 43038 9650 43090 9662
rect 43710 9714 43762 9726
rect 43710 9650 43762 9662
rect 19630 9602 19682 9614
rect 19630 9538 19682 9550
rect 19854 9602 19906 9614
rect 19854 9538 19906 9550
rect 26574 9602 26626 9614
rect 26574 9538 26626 9550
rect 28030 9602 28082 9614
rect 28030 9538 28082 9550
rect 34750 9602 34802 9614
rect 34750 9538 34802 9550
rect 36094 9602 36146 9614
rect 36094 9538 36146 9550
rect 36542 9602 36594 9614
rect 36542 9538 36594 9550
rect 38782 9602 38834 9614
rect 38782 9538 38834 9550
rect 40238 9602 40290 9614
rect 40238 9538 40290 9550
rect 40910 9602 40962 9614
rect 40910 9538 40962 9550
rect 41246 9602 41298 9614
rect 41246 9538 41298 9550
rect 41582 9602 41634 9614
rect 41582 9538 41634 9550
rect 18510 9490 18562 9502
rect 18510 9426 18562 9438
rect 18958 9490 19010 9502
rect 18958 9426 19010 9438
rect 23662 9490 23714 9502
rect 35198 9490 35250 9502
rect 32498 9438 32510 9490
rect 32562 9438 32574 9490
rect 23662 9426 23714 9438
rect 35198 9426 35250 9438
rect 35646 9490 35698 9502
rect 35646 9426 35698 9438
rect 23650 9326 23662 9378
rect 23714 9375 23726 9378
rect 24210 9375 24222 9378
rect 23714 9329 24222 9375
rect 23714 9326 23726 9329
rect 24210 9326 24222 9329
rect 24274 9326 24286 9378
rect 1344 9098 58576 9132
rect 1344 9046 4478 9098
rect 4530 9046 4582 9098
rect 4634 9046 4686 9098
rect 4738 9046 35198 9098
rect 35250 9046 35302 9098
rect 35354 9046 35406 9098
rect 35458 9046 58576 9098
rect 1344 9012 58576 9046
rect 21298 8878 21310 8930
rect 21362 8878 21374 8930
rect 35522 8878 35534 8930
rect 35586 8878 35598 8930
rect 44034 8878 44046 8930
rect 44098 8878 44110 8930
rect 28254 8818 28306 8830
rect 41122 8766 41134 8818
rect 41186 8766 41198 8818
rect 28254 8754 28306 8766
rect 19854 8706 19906 8718
rect 19854 8642 19906 8654
rect 20302 8706 20354 8718
rect 20302 8642 20354 8654
rect 22766 8706 22818 8718
rect 22766 8642 22818 8654
rect 23326 8706 23378 8718
rect 23326 8642 23378 8654
rect 30270 8706 30322 8718
rect 30270 8642 30322 8654
rect 30718 8706 30770 8718
rect 30718 8642 30770 8654
rect 36206 8706 36258 8718
rect 36206 8642 36258 8654
rect 42030 8706 42082 8718
rect 42030 8642 42082 8654
rect 19406 8594 19458 8606
rect 19406 8530 19458 8542
rect 23662 8594 23714 8606
rect 23662 8530 23714 8542
rect 23886 8594 23938 8606
rect 23886 8530 23938 8542
rect 25006 8594 25058 8606
rect 25006 8530 25058 8542
rect 29262 8594 29314 8606
rect 29262 8530 29314 8542
rect 29822 8594 29874 8606
rect 29822 8530 29874 8542
rect 31390 8594 31442 8606
rect 31390 8530 31442 8542
rect 31614 8594 31666 8606
rect 31614 8530 31666 8542
rect 32062 8594 32114 8606
rect 32062 8530 32114 8542
rect 32734 8594 32786 8606
rect 32734 8530 32786 8542
rect 37326 8594 37378 8606
rect 37326 8530 37378 8542
rect 37662 8594 37714 8606
rect 41806 8594 41858 8606
rect 40338 8542 40350 8594
rect 40402 8542 40414 8594
rect 37662 8530 37714 8542
rect 41806 8530 41858 8542
rect 43262 8594 43314 8606
rect 43262 8530 43314 8542
rect 18958 8482 19010 8494
rect 18958 8418 19010 8430
rect 20750 8482 20802 8494
rect 20750 8418 20802 8430
rect 22206 8482 22258 8494
rect 22206 8418 22258 8430
rect 24222 8482 24274 8494
rect 24222 8418 24274 8430
rect 27246 8482 27298 8494
rect 27246 8418 27298 8430
rect 31166 8482 31218 8494
rect 31166 8418 31218 8430
rect 35086 8482 35138 8494
rect 42254 8482 42306 8494
rect 40002 8430 40014 8482
rect 40066 8430 40078 8482
rect 35086 8418 35138 8430
rect 42254 8418 42306 8430
rect 1344 8090 58576 8124
rect 1344 8038 19838 8090
rect 19890 8038 19942 8090
rect 19994 8038 20046 8090
rect 20098 8038 50558 8090
rect 50610 8038 50662 8090
rect 50714 8038 50766 8090
rect 50818 8038 58576 8090
rect 1344 8004 58576 8038
rect 30258 7870 30270 7922
rect 30322 7919 30334 7922
rect 31266 7919 31278 7922
rect 30322 7873 31278 7919
rect 30322 7870 30334 7873
rect 31266 7870 31278 7873
rect 31330 7870 31342 7922
rect 37090 7870 37102 7922
rect 37154 7919 37166 7922
rect 37650 7919 37662 7922
rect 37154 7873 37662 7919
rect 37154 7870 37166 7873
rect 37650 7870 37662 7873
rect 37714 7870 37726 7922
rect 24670 7810 24722 7822
rect 24670 7746 24722 7758
rect 30270 7810 30322 7822
rect 30270 7746 30322 7758
rect 30718 7810 30770 7822
rect 30718 7746 30770 7758
rect 31166 7810 31218 7822
rect 31166 7746 31218 7758
rect 34078 7810 34130 7822
rect 34078 7746 34130 7758
rect 36654 7810 36706 7822
rect 36654 7746 36706 7758
rect 37102 7810 37154 7822
rect 37102 7746 37154 7758
rect 37550 7810 37602 7822
rect 37550 7746 37602 7758
rect 40350 7810 40402 7822
rect 40350 7746 40402 7758
rect 41022 7810 41074 7822
rect 41022 7746 41074 7758
rect 41470 7810 41522 7822
rect 41470 7746 41522 7758
rect 41918 7810 41970 7822
rect 41918 7746 41970 7758
rect 25230 7698 25282 7710
rect 25230 7634 25282 7646
rect 29262 7698 29314 7710
rect 29262 7634 29314 7646
rect 33406 7698 33458 7710
rect 35870 7698 35922 7710
rect 34514 7646 34526 7698
rect 34578 7646 34590 7698
rect 33406 7634 33458 7646
rect 35870 7634 35922 7646
rect 19406 7586 19458 7598
rect 19406 7522 19458 7534
rect 19518 7586 19570 7598
rect 19518 7522 19570 7534
rect 19966 7586 20018 7598
rect 19966 7522 20018 7534
rect 20638 7586 20690 7598
rect 20638 7522 20690 7534
rect 22990 7586 23042 7598
rect 22990 7522 23042 7534
rect 25118 7586 25170 7598
rect 25118 7522 25170 7534
rect 25902 7586 25954 7598
rect 25902 7522 25954 7534
rect 26126 7586 26178 7598
rect 26126 7522 26178 7534
rect 33070 7586 33122 7598
rect 33070 7522 33122 7534
rect 33742 7586 33794 7598
rect 33742 7522 33794 7534
rect 35198 7586 35250 7598
rect 35198 7522 35250 7534
rect 31950 7474 32002 7486
rect 31950 7410 32002 7422
rect 32398 7474 32450 7486
rect 32398 7410 32450 7422
rect 23998 7362 24050 7374
rect 23998 7298 24050 7310
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 35746 6862 35758 6914
rect 35810 6862 35822 6914
rect 32834 6750 32846 6802
rect 32898 6750 32910 6802
rect 25678 6690 25730 6702
rect 25678 6626 25730 6638
rect 21198 6578 21250 6590
rect 21198 6514 21250 6526
rect 21534 6578 21586 6590
rect 21534 6514 21586 6526
rect 21982 6578 22034 6590
rect 21982 6514 22034 6526
rect 22654 6578 22706 6590
rect 22654 6514 22706 6526
rect 29262 6578 29314 6590
rect 33630 6578 33682 6590
rect 31826 6526 31838 6578
rect 31890 6526 31902 6578
rect 29262 6514 29314 6526
rect 33630 6514 33682 6526
rect 33854 6578 33906 6590
rect 33854 6514 33906 6526
rect 28478 6466 28530 6478
rect 28478 6402 28530 6414
rect 29934 6466 29986 6478
rect 29934 6402 29986 6414
rect 34974 6466 35026 6478
rect 34974 6402 35026 6414
rect 4174 6354 4226 6366
rect 4174 6290 4226 6302
rect 4622 6354 4674 6366
rect 4622 6290 4674 6302
rect 18174 6354 18226 6366
rect 18174 6290 18226 6302
rect 20526 6354 20578 6366
rect 20526 6290 20578 6302
rect 25342 6354 25394 6366
rect 33618 6302 33630 6354
rect 33682 6302 33694 6354
rect 25342 6290 25394 6302
rect 1344 6074 58576 6108
rect 1344 6022 19838 6074
rect 19890 6022 19942 6074
rect 19994 6022 20046 6074
rect 20098 6022 50558 6074
rect 50610 6022 50662 6074
rect 50714 6022 50766 6074
rect 50818 6022 58576 6074
rect 1344 5988 58576 6022
rect 27010 5854 27022 5906
rect 27074 5903 27086 5906
rect 27906 5903 27918 5906
rect 27074 5857 27918 5903
rect 27074 5854 27086 5857
rect 27906 5854 27918 5857
rect 27970 5854 27982 5906
rect 20078 5794 20130 5806
rect 20078 5730 20130 5742
rect 20526 5794 20578 5806
rect 20526 5730 20578 5742
rect 20974 5794 21026 5806
rect 20974 5730 21026 5742
rect 22542 5794 22594 5806
rect 22542 5730 22594 5742
rect 24334 5794 24386 5806
rect 24334 5730 24386 5742
rect 25342 5794 25394 5806
rect 25342 5730 25394 5742
rect 27022 5794 27074 5806
rect 27022 5730 27074 5742
rect 27470 5794 27522 5806
rect 27470 5730 27522 5742
rect 27918 5794 27970 5806
rect 27918 5730 27970 5742
rect 28366 5794 28418 5806
rect 28366 5730 28418 5742
rect 32398 5794 32450 5806
rect 32398 5730 32450 5742
rect 21534 5682 21586 5694
rect 21534 5618 21586 5630
rect 21870 5682 21922 5694
rect 21870 5618 21922 5630
rect 22206 5682 22258 5694
rect 23662 5682 23714 5694
rect 22978 5630 22990 5682
rect 23042 5630 23054 5682
rect 22206 5618 22258 5630
rect 23662 5618 23714 5630
rect 29262 5570 29314 5582
rect 33070 5570 33122 5582
rect 28802 5518 28814 5570
rect 28866 5518 28878 5570
rect 31826 5518 31838 5570
rect 31890 5518 31902 5570
rect 33618 5518 33630 5570
rect 33682 5518 33694 5570
rect 29262 5506 29314 5518
rect 33070 5506 33122 5518
rect 25902 5458 25954 5470
rect 25902 5394 25954 5406
rect 26350 5458 26402 5470
rect 26350 5394 26402 5406
rect 31502 5458 31554 5470
rect 36082 5406 36094 5458
rect 36146 5406 36158 5458
rect 31502 5394 31554 5406
rect 25442 5294 25454 5346
rect 25506 5343 25518 5346
rect 26114 5343 26126 5346
rect 25506 5297 26126 5343
rect 25506 5294 25518 5297
rect 26114 5294 26126 5297
rect 26178 5343 26190 5346
rect 26338 5343 26350 5346
rect 26178 5297 26350 5343
rect 26178 5294 26190 5297
rect 26338 5294 26350 5297
rect 26402 5294 26414 5346
rect 1344 5066 58576 5100
rect 1344 5014 4478 5066
rect 4530 5014 4582 5066
rect 4634 5014 4686 5066
rect 4738 5014 35198 5066
rect 35250 5014 35302 5066
rect 35354 5014 35406 5066
rect 35458 5014 58576 5066
rect 1344 4980 58576 5014
rect 32386 4846 32398 4898
rect 32450 4895 32462 4898
rect 32834 4895 32846 4898
rect 32450 4849 32846 4895
rect 32450 4846 32462 4849
rect 32834 4846 32846 4849
rect 32898 4895 32910 4898
rect 33506 4895 33518 4898
rect 32898 4849 33518 4895
rect 32898 4846 32910 4849
rect 33506 4846 33518 4849
rect 33570 4846 33582 4898
rect 23998 4674 24050 4686
rect 23998 4610 24050 4622
rect 24670 4674 24722 4686
rect 24670 4610 24722 4622
rect 25454 4674 25506 4686
rect 25454 4610 25506 4622
rect 27694 4674 27746 4686
rect 27694 4610 27746 4622
rect 28478 4674 28530 4686
rect 28478 4610 28530 4622
rect 28926 4674 28978 4686
rect 28926 4610 28978 4622
rect 32398 4674 32450 4686
rect 32398 4610 32450 4622
rect 32846 4674 32898 4686
rect 32846 4610 32898 4622
rect 33294 4674 33346 4686
rect 33294 4610 33346 4622
rect 33742 4674 33794 4686
rect 33742 4610 33794 4622
rect 1344 4058 58576 4092
rect 1344 4006 19838 4058
rect 19890 4006 19942 4058
rect 19994 4006 20046 4058
rect 20098 4006 50558 4058
rect 50610 4006 50662 4058
rect 50714 4006 50766 4058
rect 50818 4006 58576 4058
rect 1344 3972 58576 4006
<< via1 >>
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4478 55414 4530 55466
rect 4582 55414 4634 55466
rect 4686 55414 4738 55466
rect 35198 55414 35250 55466
rect 35302 55414 35354 55466
rect 35406 55414 35458 55466
rect 19838 54406 19890 54458
rect 19942 54406 19994 54458
rect 20046 54406 20098 54458
rect 50558 54406 50610 54458
rect 50662 54406 50714 54458
rect 50766 54406 50818 54458
rect 55246 54126 55298 54178
rect 4478 53398 4530 53450
rect 4582 53398 4634 53450
rect 4686 53398 4738 53450
rect 35198 53398 35250 53450
rect 35302 53398 35354 53450
rect 35406 53398 35458 53450
rect 19838 52390 19890 52442
rect 19942 52390 19994 52442
rect 20046 52390 20098 52442
rect 50558 52390 50610 52442
rect 50662 52390 50714 52442
rect 50766 52390 50818 52442
rect 5854 52110 5906 52162
rect 4478 51382 4530 51434
rect 4582 51382 4634 51434
rect 4686 51382 4738 51434
rect 35198 51382 35250 51434
rect 35302 51382 35354 51434
rect 35406 51382 35458 51434
rect 19838 50374 19890 50426
rect 19942 50374 19994 50426
rect 20046 50374 20098 50426
rect 50558 50374 50610 50426
rect 50662 50374 50714 50426
rect 50766 50374 50818 50426
rect 36990 49758 37042 49810
rect 41358 49758 41410 49810
rect 41806 49758 41858 49810
rect 42254 49758 42306 49810
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 41694 48974 41746 49026
rect 31278 48862 31330 48914
rect 32734 48862 32786 48914
rect 30830 48750 30882 48802
rect 31950 48750 32002 48802
rect 37438 48750 37490 48802
rect 40798 48750 40850 48802
rect 41246 48750 41298 48802
rect 42142 48750 42194 48802
rect 42366 48750 42418 48802
rect 34862 48638 34914 48690
rect 36430 48638 36482 48690
rect 38110 48638 38162 48690
rect 40126 48638 40178 48690
rect 43374 48638 43426 48690
rect 44158 48638 44210 48690
rect 19838 48358 19890 48410
rect 19942 48358 19994 48410
rect 20046 48358 20098 48410
rect 50558 48358 50610 48410
rect 50662 48358 50714 48410
rect 50766 48358 50818 48410
rect 6190 48078 6242 48130
rect 41806 48078 41858 48130
rect 43710 48078 43762 48130
rect 37102 47966 37154 48018
rect 39342 47966 39394 48018
rect 42814 47966 42866 48018
rect 3390 47854 3442 47906
rect 3950 47854 4002 47906
rect 26014 47854 26066 47906
rect 26574 47854 26626 47906
rect 36766 47854 36818 47906
rect 40350 47854 40402 47906
rect 40798 47854 40850 47906
rect 41470 47854 41522 47906
rect 43486 47854 43538 47906
rect 3054 47742 3106 47794
rect 24670 47742 24722 47794
rect 25566 47742 25618 47794
rect 28702 47742 28754 47794
rect 35422 47742 35474 47794
rect 35870 47742 35922 47794
rect 36318 47742 36370 47794
rect 6526 47630 6578 47682
rect 35422 47518 35474 47570
rect 35870 47518 35922 47570
rect 36654 47518 36706 47570
rect 4478 47350 4530 47402
rect 4582 47350 4634 47402
rect 4686 47350 4738 47402
rect 35198 47350 35250 47402
rect 35302 47350 35354 47402
rect 35406 47350 35458 47402
rect 34862 47182 34914 47234
rect 5630 46958 5682 47010
rect 5742 46958 5794 47010
rect 6302 47070 6354 47122
rect 38670 47070 38722 47122
rect 39454 47070 39506 47122
rect 40014 47070 40066 47122
rect 39454 46958 39506 47010
rect 5742 46846 5794 46898
rect 22542 46846 22594 46898
rect 22990 46846 23042 46898
rect 25006 46846 25058 46898
rect 39006 46846 39058 46898
rect 40238 46846 40290 46898
rect 40686 46846 40738 46898
rect 30494 46734 30546 46786
rect 31502 46734 31554 46786
rect 6190 46622 6242 46674
rect 21646 46622 21698 46674
rect 22094 46622 22146 46674
rect 25790 46622 25842 46674
rect 26350 46622 26402 46674
rect 27582 46622 27634 46674
rect 29262 46622 29314 46674
rect 29710 46622 29762 46674
rect 30158 46622 30210 46674
rect 39902 46622 39954 46674
rect 42926 46622 42978 46674
rect 29262 46510 29314 46562
rect 30158 46510 30210 46562
rect 38894 46510 38946 46562
rect 39902 46510 39954 46562
rect 44046 46510 44098 46562
rect 19838 46342 19890 46394
rect 19942 46342 19994 46394
rect 20046 46342 20098 46394
rect 50558 46342 50610 46394
rect 50662 46342 50714 46394
rect 50766 46342 50818 46394
rect 7198 46062 7250 46114
rect 27806 46062 27858 46114
rect 30942 46062 30994 46114
rect 41134 46062 41186 46114
rect 41582 46062 41634 46114
rect 28590 45950 28642 46002
rect 4510 45838 4562 45890
rect 5070 45838 5122 45890
rect 8430 45838 8482 45890
rect 11678 45838 11730 45890
rect 28142 45838 28194 45890
rect 35086 45838 35138 45890
rect 35870 45838 35922 45890
rect 36430 45838 36482 45890
rect 38558 45838 38610 45890
rect 46062 45838 46114 45890
rect 48190 45838 48242 45890
rect 1822 45726 1874 45778
rect 4174 45726 4226 45778
rect 9662 45726 9714 45778
rect 26462 45726 26514 45778
rect 26910 45726 26962 45778
rect 27358 45726 27410 45778
rect 33182 45726 33234 45778
rect 34638 45726 34690 45778
rect 35534 45726 35586 45778
rect 7646 45614 7698 45666
rect 26574 45614 26626 45666
rect 26910 45614 26962 45666
rect 27358 45614 27410 45666
rect 28142 45614 28194 45666
rect 31838 45614 31890 45666
rect 40014 45614 40066 45666
rect 43150 45614 43202 45666
rect 8318 45502 8370 45554
rect 11566 45502 11618 45554
rect 4478 45334 4530 45386
rect 4582 45334 4634 45386
rect 4686 45334 4738 45386
rect 35198 45334 35250 45386
rect 35302 45334 35354 45386
rect 35406 45334 35458 45386
rect 5630 45166 5682 45218
rect 22094 45166 22146 45218
rect 22990 45166 23042 45218
rect 12798 45054 12850 45106
rect 22206 44942 22258 44994
rect 28590 44942 28642 44994
rect 37662 44942 37714 44994
rect 1822 44830 1874 44882
rect 2382 44830 2434 44882
rect 5742 44830 5794 44882
rect 6078 44830 6130 44882
rect 6638 44830 6690 44882
rect 9662 44830 9714 44882
rect 10222 44830 10274 44882
rect 23438 44830 23490 44882
rect 23998 44830 24050 44882
rect 26350 44830 26402 44882
rect 26686 44830 26738 44882
rect 29486 44830 29538 44882
rect 29934 44830 29986 44882
rect 30270 44830 30322 44882
rect 32622 44830 32674 44882
rect 33182 44830 33234 44882
rect 41470 44830 41522 44882
rect 45614 44830 45666 44882
rect 38334 44718 38386 44770
rect 46510 44718 46562 44770
rect 47294 44718 47346 44770
rect 4510 44606 4562 44658
rect 4958 44606 5010 44658
rect 8766 44606 8818 44658
rect 9214 44606 9266 44658
rect 12350 44606 12402 44658
rect 22654 44606 22706 44658
rect 23102 44606 23154 44658
rect 33630 44606 33682 44658
rect 35646 44606 35698 44658
rect 36430 44606 36482 44658
rect 37214 44606 37266 44658
rect 38894 44606 38946 44658
rect 41134 44606 41186 44658
rect 42254 44606 42306 44658
rect 45166 44606 45218 44658
rect 27806 44494 27858 44546
rect 19838 44326 19890 44378
rect 19942 44326 19994 44378
rect 20046 44326 20098 44378
rect 50558 44326 50610 44378
rect 50662 44326 50714 44378
rect 50766 44326 50818 44378
rect 10222 44158 10274 44210
rect 1822 44046 1874 44098
rect 4846 44046 4898 44098
rect 8542 44046 8594 44098
rect 8878 44046 8930 44098
rect 9886 44046 9938 44098
rect 10334 44046 10386 44098
rect 13582 44046 13634 44098
rect 27246 44046 27298 44098
rect 33294 44046 33346 44098
rect 35646 44046 35698 44098
rect 38894 44046 38946 44098
rect 43710 44046 43762 44098
rect 45390 44046 45442 44098
rect 48190 44046 48242 44098
rect 14478 43934 14530 43986
rect 18174 43934 18226 43986
rect 27694 43934 27746 43986
rect 28814 43934 28866 43986
rect 34302 43934 34354 43986
rect 35086 43934 35138 43986
rect 40910 43934 40962 43986
rect 41582 43934 41634 43986
rect 43038 43934 43090 43986
rect 2158 43822 2210 43874
rect 2718 43822 2770 43874
rect 5742 43822 5794 43874
rect 6302 43822 6354 43874
rect 10894 43822 10946 43874
rect 11454 43822 11506 43874
rect 14590 43822 14642 43874
rect 17390 43822 17442 43874
rect 28142 43822 28194 43874
rect 33518 43822 33570 43874
rect 36206 43822 36258 43874
rect 36766 43822 36818 43874
rect 41246 43822 41298 43874
rect 41918 43822 41970 43874
rect 42478 43822 42530 43874
rect 54126 43822 54178 43874
rect 16830 43710 16882 43762
rect 20190 43710 20242 43762
rect 32286 43710 32338 43762
rect 45726 43710 45778 43762
rect 46958 43710 47010 43762
rect 47406 43710 47458 43762
rect 51774 43710 51826 43762
rect 5294 43598 5346 43650
rect 14030 43598 14082 43650
rect 31390 43598 31442 43650
rect 39342 43598 39394 43650
rect 4478 43318 4530 43370
rect 4582 43318 4634 43370
rect 4686 43318 4738 43370
rect 35198 43318 35250 43370
rect 35302 43318 35354 43370
rect 35406 43318 35458 43370
rect 5630 43150 5682 43202
rect 6078 43150 6130 43202
rect 13470 43150 13522 43202
rect 12798 43038 12850 43090
rect 35870 42926 35922 42978
rect 37102 42926 37154 42978
rect 37886 42926 37938 42978
rect 46734 42926 46786 42978
rect 48078 42926 48130 42978
rect 1822 42814 1874 42866
rect 2382 42814 2434 42866
rect 5742 42814 5794 42866
rect 6190 42814 6242 42866
rect 9662 42814 9714 42866
rect 10222 42814 10274 42866
rect 13582 42814 13634 42866
rect 17054 42814 17106 42866
rect 19854 42814 19906 42866
rect 23774 42814 23826 42866
rect 31726 42814 31778 42866
rect 32398 42814 32450 42866
rect 33854 42814 33906 42866
rect 39678 42814 39730 42866
rect 40350 42814 40402 42866
rect 41806 42814 41858 42866
rect 47966 42814 48018 42866
rect 48190 42814 48242 42866
rect 22318 42702 22370 42754
rect 22542 42702 22594 42754
rect 22766 42702 22818 42754
rect 23438 42702 23490 42754
rect 32062 42702 32114 42754
rect 33294 42702 33346 42754
rect 34526 42702 34578 42754
rect 35310 42702 35362 42754
rect 40014 42702 40066 42754
rect 41134 42702 41186 42754
rect 42478 42702 42530 42754
rect 47518 42702 47570 42754
rect 47742 42702 47794 42754
rect 4622 42590 4674 42642
rect 4958 42590 5010 42642
rect 6638 42590 6690 42642
rect 9326 42590 9378 42642
rect 12350 42590 12402 42642
rect 16718 42590 16770 42642
rect 17838 42590 17890 42642
rect 21422 42590 21474 42642
rect 21870 42590 21922 42642
rect 26350 42590 26402 42642
rect 27358 42590 27410 42642
rect 27806 42590 27858 42642
rect 29374 42590 29426 42642
rect 29822 42590 29874 42642
rect 32734 42590 32786 42642
rect 40686 42590 40738 42642
rect 43934 42590 43986 42642
rect 44942 42590 44994 42642
rect 45390 42590 45442 42642
rect 45838 42590 45890 42642
rect 46286 42590 46338 42642
rect 47182 42590 47234 42642
rect 48638 42590 48690 42642
rect 49086 42590 49138 42642
rect 49534 42590 49586 42642
rect 50878 42590 50930 42642
rect 51214 42590 51266 42642
rect 51662 42590 51714 42642
rect 52110 42590 52162 42642
rect 52782 42590 52834 42642
rect 53342 42590 53394 42642
rect 53790 42590 53842 42642
rect 54238 42590 54290 42642
rect 21870 42478 21922 42530
rect 22430 42478 22482 42530
rect 44942 42478 44994 42530
rect 46286 42478 46338 42530
rect 47294 42478 47346 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 3502 42030 3554 42082
rect 6638 42030 6690 42082
rect 13470 42030 13522 42082
rect 29262 42030 29314 42082
rect 47182 42030 47234 42082
rect 52334 42030 52386 42082
rect 3390 41918 3442 41970
rect 20526 41918 20578 41970
rect 21870 41918 21922 41970
rect 26126 41918 26178 41970
rect 26462 41918 26514 41970
rect 27134 41918 27186 41970
rect 28030 41918 28082 41970
rect 28590 41918 28642 41970
rect 33406 41918 33458 41970
rect 34638 41918 34690 41970
rect 35198 41918 35250 41970
rect 35870 41918 35922 41970
rect 37998 41918 38050 41970
rect 43934 41918 43986 41970
rect 46734 41918 46786 41970
rect 47518 41918 47570 41970
rect 48862 41918 48914 41970
rect 53118 41918 53170 41970
rect 55582 41918 55634 41970
rect 3838 41806 3890 41858
rect 4398 41806 4450 41858
rect 10782 41806 10834 41858
rect 11342 41806 11394 41858
rect 13918 41806 13970 41858
rect 14478 41806 14530 41858
rect 18510 41806 18562 41858
rect 21310 41806 21362 41858
rect 26798 41806 26850 41858
rect 27470 41806 27522 41858
rect 30046 41806 30098 41858
rect 33070 41806 33122 41858
rect 33742 41806 33794 41858
rect 34078 41806 34130 41858
rect 40910 41806 40962 41858
rect 44270 41806 44322 41858
rect 44494 41806 44546 41858
rect 44718 41806 44770 41858
rect 45614 41806 45666 41858
rect 49198 41806 49250 41858
rect 49422 41806 49474 41858
rect 49758 41806 49810 41858
rect 49870 41806 49922 41858
rect 52782 41806 52834 41858
rect 53454 41806 53506 41858
rect 53790 41806 53842 41858
rect 54350 41806 54402 41858
rect 54910 41806 54962 41858
rect 1822 41694 1874 41746
rect 3054 41694 3106 41746
rect 10446 41694 10498 41746
rect 18174 41694 18226 41746
rect 30494 41694 30546 41746
rect 32510 41694 32562 41746
rect 36766 41694 36818 41746
rect 37102 41694 37154 41746
rect 37550 41694 37602 41746
rect 39902 41694 39954 41746
rect 40462 41694 40514 41746
rect 43038 41694 43090 41746
rect 43486 41694 43538 41746
rect 50878 41694 50930 41746
rect 51550 41694 51602 41746
rect 51998 41694 52050 41746
rect 6974 41582 7026 41634
rect 14366 41582 14418 41634
rect 50318 41582 50370 41634
rect 41358 41470 41410 41522
rect 45054 41470 45106 41522
rect 4478 41302 4530 41354
rect 4582 41302 4634 41354
rect 4686 41302 4738 41354
rect 35198 41302 35250 41354
rect 35302 41302 35354 41354
rect 35406 41302 35458 41354
rect 5630 41134 5682 41186
rect 17054 41134 17106 41186
rect 17614 41134 17666 41186
rect 53342 41134 53394 41186
rect 21310 41022 21362 41074
rect 22318 41022 22370 41074
rect 42590 41022 42642 41074
rect 6078 40910 6130 40962
rect 17166 40910 17218 40962
rect 17614 40910 17666 40962
rect 23550 40910 23602 40962
rect 31614 40910 31666 40962
rect 34414 40910 34466 40962
rect 34750 40910 34802 40962
rect 35870 40910 35922 40962
rect 1822 40798 1874 40850
rect 2382 40798 2434 40850
rect 5742 40798 5794 40850
rect 9662 40798 9714 40850
rect 10222 40798 10274 40850
rect 17950 40798 18002 40850
rect 20750 40798 20802 40850
rect 24222 40798 24274 40850
rect 26014 40798 26066 40850
rect 27470 40798 27522 40850
rect 30494 40798 30546 40850
rect 30718 40798 30770 40850
rect 37326 40798 37378 40850
rect 37886 40798 37938 40850
rect 38670 40798 38722 40850
rect 41582 40798 41634 40850
rect 42926 40798 42978 40850
rect 44046 40798 44098 40850
rect 45390 40798 45442 40850
rect 46174 40798 46226 40850
rect 46734 40798 46786 40850
rect 47518 40798 47570 40850
rect 53230 40798 53282 40850
rect 54462 40798 54514 40850
rect 13470 40686 13522 40738
rect 23886 40686 23938 40738
rect 29822 40686 29874 40738
rect 31166 40686 31218 40738
rect 37662 40686 37714 40738
rect 41246 40686 41298 40738
rect 43038 40686 43090 40738
rect 4510 40574 4562 40626
rect 4958 40574 5010 40626
rect 6190 40574 6242 40626
rect 9326 40574 9378 40626
rect 12350 40574 12402 40626
rect 12798 40574 12850 40626
rect 13582 40574 13634 40626
rect 18734 40574 18786 40626
rect 21422 40574 21474 40626
rect 21870 40574 21922 40626
rect 22318 40574 22370 40626
rect 23102 40574 23154 40626
rect 27582 40574 27634 40626
rect 29374 40574 29426 40626
rect 30270 40574 30322 40626
rect 37102 40574 37154 40626
rect 42366 40574 42418 40626
rect 21870 40462 21922 40514
rect 22430 40462 22482 40514
rect 27022 40462 27074 40514
rect 54574 40686 54626 40738
rect 56142 40686 56194 40738
rect 43486 40574 43538 40626
rect 44942 40574 44994 40626
rect 43486 40462 43538 40514
rect 49422 40462 49474 40514
rect 19838 40294 19890 40346
rect 19942 40294 19994 40346
rect 20046 40294 20098 40346
rect 50558 40294 50610 40346
rect 50662 40294 50714 40346
rect 50766 40294 50818 40346
rect 17390 40126 17442 40178
rect 21982 40126 22034 40178
rect 37550 40126 37602 40178
rect 1822 40014 1874 40066
rect 6862 40014 6914 40066
rect 13470 40014 13522 40066
rect 24222 40014 24274 40066
rect 24670 40014 24722 40066
rect 32286 40014 32338 40066
rect 34078 40014 34130 40066
rect 39902 40014 39954 40066
rect 43710 40014 43762 40066
rect 47854 40014 47906 40066
rect 52334 40014 52386 40066
rect 53118 40014 53170 40066
rect 54910 40014 54962 40066
rect 16830 39902 16882 39954
rect 17838 39902 17890 39954
rect 18398 39902 18450 39954
rect 19742 39902 19794 39954
rect 22430 39902 22482 39954
rect 22878 39902 22930 39954
rect 25118 39902 25170 39954
rect 25454 39902 25506 39954
rect 27134 39902 27186 39954
rect 29262 39902 29314 39954
rect 29822 39902 29874 39954
rect 30382 39902 30434 39954
rect 33070 39902 33122 39954
rect 34974 39902 35026 39954
rect 35534 39902 35586 39954
rect 38334 39902 38386 39954
rect 40910 39902 40962 39954
rect 41582 39902 41634 39954
rect 42478 39902 42530 39954
rect 43038 39902 43090 39954
rect 45054 39902 45106 39954
rect 45726 39902 45778 39954
rect 46510 39902 46562 39954
rect 47182 39902 47234 39954
rect 49198 39902 49250 39954
rect 49534 39902 49586 39954
rect 49870 39902 49922 39954
rect 50206 39902 50258 39954
rect 51102 39902 51154 39954
rect 51662 39902 51714 39954
rect 53230 39902 53282 39954
rect 54574 39902 54626 39954
rect 55582 39902 55634 39954
rect 4174 39790 4226 39842
rect 4734 39790 4786 39842
rect 10782 39790 10834 39842
rect 11342 39790 11394 39842
rect 18958 39790 19010 39842
rect 22654 39790 22706 39842
rect 28478 39790 28530 39842
rect 36430 39790 36482 39842
rect 37886 39790 37938 39842
rect 41246 39790 41298 39842
rect 41918 39790 41970 39842
rect 44494 39790 44546 39842
rect 45390 39790 45442 39842
rect 46062 39790 46114 39842
rect 50542 39790 50594 39842
rect 53006 39790 53058 39842
rect 53454 39796 53506 39848
rect 54014 39790 54066 39842
rect 54350 39790 54402 39842
rect 55358 39790 55410 39842
rect 3838 39678 3890 39730
rect 10446 39678 10498 39730
rect 16494 39678 16546 39730
rect 18510 39678 18562 39730
rect 29934 39678 29986 39730
rect 35646 39678 35698 39730
rect 36990 39678 37042 39730
rect 56702 39678 56754 39730
rect 57150 39678 57202 39730
rect 7310 39566 7362 39618
rect 13918 39566 13970 39618
rect 21758 39566 21810 39618
rect 27918 39566 27970 39618
rect 28366 39566 28418 39618
rect 36094 39566 36146 39618
rect 28814 39454 28866 39506
rect 34526 39454 34578 39506
rect 4478 39286 4530 39338
rect 4582 39286 4634 39338
rect 4686 39286 4738 39338
rect 35198 39286 35250 39338
rect 35302 39286 35354 39338
rect 35406 39286 35458 39338
rect 4958 39118 5010 39170
rect 12686 39118 12738 39170
rect 18062 39118 18114 39170
rect 19518 39118 19570 39170
rect 37214 39118 37266 39170
rect 38334 39118 38386 39170
rect 21646 39006 21698 39058
rect 25454 39006 25506 39058
rect 36990 39006 37042 39058
rect 37774 39006 37826 39058
rect 39230 39006 39282 39058
rect 17390 38894 17442 38946
rect 28030 38894 28082 38946
rect 29374 38894 29426 38946
rect 30046 38894 30098 38946
rect 32510 38894 32562 38946
rect 34414 38894 34466 38946
rect 37214 38894 37266 38946
rect 37662 38894 37714 38946
rect 38110 38894 38162 38946
rect 38558 38894 38610 38946
rect 43038 38894 43090 38946
rect 50878 38894 50930 38946
rect 51774 38894 51826 38946
rect 52782 38894 52834 38946
rect 54686 38894 54738 38946
rect 8318 38782 8370 38834
rect 8878 38782 8930 38834
rect 12798 38782 12850 38834
rect 18734 38782 18786 38834
rect 19966 38782 20018 38834
rect 22654 38782 22706 38834
rect 26574 38782 26626 38834
rect 27582 38782 27634 38834
rect 28478 38782 28530 38834
rect 33630 38782 33682 38834
rect 42254 38782 42306 38834
rect 46734 38782 46786 38834
rect 55358 38782 55410 38834
rect 56478 38782 56530 38834
rect 4622 38670 4674 38722
rect 5070 38670 5122 38722
rect 5742 38670 5794 38722
rect 13470 38670 13522 38722
rect 16606 38670 16658 38722
rect 17838 38670 17890 38722
rect 18510 38670 18562 38722
rect 18958 38670 19010 38722
rect 20414 38670 20466 38722
rect 20638 38670 20690 38722
rect 21310 38670 21362 38722
rect 27134 38670 27186 38722
rect 27246 38670 27298 38722
rect 33182 38670 33234 38722
rect 33742 38670 33794 38722
rect 38894 38670 38946 38722
rect 40462 38670 40514 38722
rect 41134 38670 41186 38722
rect 42702 38670 42754 38722
rect 47182 38670 47234 38722
rect 47406 38670 47458 38722
rect 6078 38558 6130 38610
rect 13582 38558 13634 38610
rect 17054 38558 17106 38610
rect 22206 38558 22258 38610
rect 23438 38558 23490 38610
rect 27806 38558 27858 38610
rect 28254 38558 28306 38610
rect 39790 38558 39842 38610
rect 41918 38558 41970 38610
rect 44942 38558 44994 38610
rect 49982 38558 50034 38610
rect 50430 38558 50482 38610
rect 51326 38558 51378 38610
rect 53230 38558 53282 38610
rect 53678 38558 53730 38610
rect 57038 38558 57090 38610
rect 26126 38446 26178 38498
rect 32734 38446 32786 38498
rect 46286 38446 46338 38498
rect 49982 38446 50034 38498
rect 51326 38446 51378 38498
rect 52558 38446 52610 38498
rect 53230 38446 53282 38498
rect 53678 38446 53730 38498
rect 19838 38278 19890 38330
rect 19942 38278 19994 38330
rect 20046 38278 20098 38330
rect 50558 38278 50610 38330
rect 50662 38278 50714 38330
rect 50766 38278 50818 38330
rect 7086 38110 7138 38162
rect 7534 38110 7586 38162
rect 18846 38110 18898 38162
rect 19406 38110 19458 38162
rect 27470 38110 27522 38162
rect 33742 38110 33794 38162
rect 36318 38110 36370 38162
rect 39230 38110 39282 38162
rect 39790 38110 39842 38162
rect 49310 38110 49362 38162
rect 49646 38110 49698 38162
rect 50654 38110 50706 38162
rect 51662 38110 51714 38162
rect 6190 37998 6242 38050
rect 7198 37998 7250 38050
rect 14366 37998 14418 38050
rect 17502 37998 17554 38050
rect 17950 37998 18002 38050
rect 19518 37998 19570 38050
rect 25454 37998 25506 38050
rect 28142 37998 28194 38050
rect 28590 37998 28642 38050
rect 38782 37998 38834 38050
rect 41918 37998 41970 38050
rect 48190 37998 48242 38050
rect 49310 37998 49362 38050
rect 50206 37998 50258 38050
rect 50654 37998 50706 38050
rect 56030 37998 56082 38050
rect 20414 37886 20466 37938
rect 21534 37886 21586 37938
rect 21758 37886 21810 37938
rect 22094 37886 22146 37938
rect 23550 37886 23602 37938
rect 25790 37886 25842 37938
rect 26462 37886 26514 37938
rect 27022 37886 27074 37938
rect 41246 37886 41298 37938
rect 41582 37886 41634 37938
rect 43710 37886 43762 37938
rect 46846 37886 46898 37938
rect 47294 37886 47346 37938
rect 52558 37886 52610 37938
rect 3502 37774 3554 37826
rect 4062 37774 4114 37826
rect 7646 37774 7698 37826
rect 11678 37774 11730 37826
rect 12238 37774 12290 37826
rect 18398 37774 18450 37826
rect 19406 37774 19458 37826
rect 19966 37774 20018 37826
rect 20302 37774 20354 37826
rect 21086 37774 21138 37826
rect 21310 37774 21362 37826
rect 22654 37774 22706 37826
rect 25118 37774 25170 37826
rect 26014 37774 26066 37826
rect 35310 37774 35362 37826
rect 36654 37774 36706 37826
rect 40910 37774 40962 37826
rect 42478 37774 42530 37826
rect 43038 37774 43090 37826
rect 45278 37774 45330 37826
rect 51550 37774 51602 37826
rect 52726 37774 52778 37826
rect 53790 37774 53842 37826
rect 3166 37662 3218 37714
rect 11342 37662 11394 37714
rect 16830 37662 16882 37714
rect 18846 37662 18898 37714
rect 23214 37662 23266 37714
rect 25566 37662 25618 37714
rect 26350 37662 26402 37714
rect 32510 37662 32562 37714
rect 39230 37662 39282 37714
rect 39678 37662 39730 37714
rect 40350 37662 40402 37714
rect 44942 37662 44994 37714
rect 47518 37662 47570 37714
rect 48862 37662 48914 37714
rect 49758 37662 49810 37714
rect 51102 37662 51154 37714
rect 55582 37662 55634 37714
rect 56702 37662 56754 37714
rect 57150 37662 57202 37714
rect 57598 37662 57650 37714
rect 6638 37550 6690 37602
rect 14814 37550 14866 37602
rect 51102 37550 51154 37602
rect 51326 37550 51378 37602
rect 21198 37438 21250 37490
rect 22206 37438 22258 37490
rect 22542 37438 22594 37490
rect 46398 37438 46450 37490
rect 49758 37438 49810 37490
rect 50206 37438 50258 37490
rect 54350 37438 54402 37490
rect 4478 37270 4530 37322
rect 4582 37270 4634 37322
rect 4686 37270 4738 37322
rect 35198 37270 35250 37322
rect 35302 37270 35354 37322
rect 35406 37270 35458 37322
rect 4398 37102 4450 37154
rect 23102 37102 23154 37154
rect 33070 37102 33122 37154
rect 43822 37102 43874 37154
rect 8766 36878 8818 36930
rect 14702 36878 14754 36930
rect 19182 36878 19234 36930
rect 20750 36878 20802 36930
rect 24782 36878 24834 36930
rect 37326 36878 37378 36930
rect 37998 36878 38050 36930
rect 50430 36878 50482 36930
rect 4510 36766 4562 36818
rect 5630 36766 5682 36818
rect 6190 36766 6242 36818
rect 15038 36766 15090 36818
rect 17838 36766 17890 36818
rect 20414 36766 20466 36818
rect 21310 36766 21362 36818
rect 23550 36766 23602 36818
rect 30718 36766 30770 36818
rect 32510 36766 32562 36818
rect 42926 36766 42978 36818
rect 43038 36766 43090 36818
rect 43934 36766 43986 36818
rect 44046 36766 44098 36818
rect 46174 36766 46226 36818
rect 49646 36766 49698 36818
rect 49870 36766 49922 36818
rect 50094 36766 50146 36818
rect 50318 36766 50370 36818
rect 50654 36766 50706 36818
rect 51550 36878 51602 36930
rect 51438 36766 51490 36818
rect 53678 36766 53730 36818
rect 56926 36766 56978 36818
rect 57486 36766 57538 36818
rect 18510 36654 18562 36706
rect 19070 36654 19122 36706
rect 20078 36654 20130 36706
rect 21982 36654 22034 36706
rect 22206 36654 22258 36706
rect 22430 36654 22482 36706
rect 22654 36654 22706 36706
rect 23998 36654 24050 36706
rect 24222 36654 24274 36706
rect 29262 36654 29314 36706
rect 29374 36654 29426 36706
rect 29934 36654 29986 36706
rect 37662 36654 37714 36706
rect 38334 36654 38386 36706
rect 38670 36654 38722 36706
rect 39006 36654 39058 36706
rect 39902 36654 39954 36706
rect 40462 36654 40514 36706
rect 45502 36654 45554 36706
rect 46062 36654 46114 36706
rect 46734 36654 46786 36706
rect 47070 36654 47122 36706
rect 47742 36654 47794 36706
rect 50542 36654 50594 36706
rect 50878 36654 50930 36706
rect 51214 36654 51266 36706
rect 52110 36654 52162 36706
rect 53006 36654 53058 36706
rect 53342 36654 53394 36706
rect 54462 36654 54514 36706
rect 55134 36654 55186 36706
rect 57150 36654 57202 36706
rect 57934 36654 57986 36706
rect 4062 36542 4114 36594
rect 4958 36542 5010 36594
rect 8318 36542 8370 36594
rect 11006 36542 11058 36594
rect 13582 36542 13634 36594
rect 15822 36542 15874 36594
rect 18062 36542 18114 36594
rect 21646 36542 21698 36594
rect 28590 36542 28642 36594
rect 32174 36542 32226 36594
rect 35982 36542 36034 36594
rect 36430 36542 36482 36594
rect 39342 36542 39394 36594
rect 41134 36542 41186 36594
rect 41918 36542 41970 36594
rect 51662 36542 51714 36594
rect 54014 36542 54066 36594
rect 55806 36542 55858 36594
rect 56590 36542 56642 36594
rect 4846 36430 4898 36482
rect 13470 36430 13522 36482
rect 22766 36430 22818 36482
rect 30382 36430 30434 36482
rect 45054 36430 45106 36482
rect 48862 36430 48914 36482
rect 19838 36262 19890 36314
rect 19942 36262 19994 36314
rect 20046 36262 20098 36314
rect 50558 36262 50610 36314
rect 50662 36262 50714 36314
rect 50766 36262 50818 36314
rect 3726 36094 3778 36146
rect 4510 36094 4562 36146
rect 37998 36094 38050 36146
rect 39790 36094 39842 36146
rect 2718 35982 2770 36034
rect 5854 35982 5906 36034
rect 6190 35982 6242 36034
rect 21310 35982 21362 36034
rect 21758 35982 21810 36034
rect 21982 35982 22034 36034
rect 24782 35982 24834 36034
rect 25342 35982 25394 36034
rect 30158 35982 30210 36034
rect 36318 35982 36370 36034
rect 40798 35982 40850 36034
rect 44382 35982 44434 36034
rect 44830 35982 44882 36034
rect 45614 35982 45666 36034
rect 46734 35982 46786 36034
rect 48302 35982 48354 36034
rect 51550 35982 51602 36034
rect 52334 35982 52386 36034
rect 56702 35982 56754 36034
rect 12126 35870 12178 35922
rect 14478 35870 14530 35922
rect 18958 35870 19010 35922
rect 19070 35870 19122 35922
rect 19742 35870 19794 35922
rect 22878 35870 22930 35922
rect 23774 35870 23826 35922
rect 25566 35870 25618 35922
rect 25790 35870 25842 35922
rect 27022 35870 27074 35922
rect 43150 35870 43202 35922
rect 49086 35870 49138 35922
rect 49422 35870 49474 35922
rect 50318 35870 50370 35922
rect 54238 35870 54290 35922
rect 3054 35758 3106 35810
rect 3614 35758 3666 35810
rect 10782 35758 10834 35810
rect 11342 35758 11394 35810
rect 14590 35758 14642 35810
rect 18398 35758 18450 35810
rect 19518 35758 19570 35810
rect 19630 35758 19682 35810
rect 19966 35758 20018 35810
rect 24110 35758 24162 35810
rect 24334 35758 24386 35810
rect 25118 35758 25170 35810
rect 25902 35758 25954 35810
rect 26238 35758 26290 35810
rect 29374 35758 29426 35810
rect 32174 35758 32226 35810
rect 34974 35758 35026 35810
rect 36766 35758 36818 35810
rect 37326 35758 37378 35810
rect 38894 35758 38946 35810
rect 39230 35758 39282 35810
rect 41246 35758 41298 35810
rect 43486 35758 43538 35810
rect 48750 35758 48802 35810
rect 49758 35758 49810 35810
rect 50878 35758 50930 35810
rect 53454 35758 53506 35810
rect 53678 35758 53730 35810
rect 54014 35758 54066 35810
rect 54574 35758 54626 35810
rect 55918 35758 55970 35810
rect 10894 35646 10946 35698
rect 20526 35646 20578 35698
rect 22542 35646 22594 35698
rect 23214 35646 23266 35698
rect 40350 35646 40402 35698
rect 43934 35646 43986 35698
rect 57150 35646 57202 35698
rect 57598 35646 57650 35698
rect 10110 35534 10162 35586
rect 14142 35534 14194 35586
rect 29038 35534 29090 35586
rect 34638 35534 34690 35586
rect 53566 35534 53618 35586
rect 17950 35422 18002 35474
rect 22094 35422 22146 35474
rect 22318 35422 22370 35474
rect 22654 35422 22706 35474
rect 22878 35422 22930 35474
rect 55582 35422 55634 35474
rect 56702 35422 56754 35474
rect 57374 35422 57426 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 55470 35086 55522 35138
rect 13582 34974 13634 35026
rect 5630 34862 5682 34914
rect 15486 34862 15538 34914
rect 19182 34862 19234 34914
rect 22878 34862 22930 34914
rect 34750 34862 34802 34914
rect 35646 34862 35698 34914
rect 38782 34862 38834 34914
rect 44270 34862 44322 34914
rect 46398 34862 46450 34914
rect 53902 34862 53954 34914
rect 1822 34750 1874 34802
rect 2382 34750 2434 34802
rect 9774 34750 9826 34802
rect 10446 34750 10498 34802
rect 13470 34750 13522 34802
rect 13694 34750 13746 34802
rect 15822 34750 15874 34802
rect 18622 34750 18674 34802
rect 20190 34750 20242 34802
rect 22542 34750 22594 34802
rect 23326 34750 23378 34802
rect 23550 34750 23602 34802
rect 24446 34750 24498 34802
rect 27358 34750 27410 34802
rect 29262 34750 29314 34802
rect 32062 34750 32114 34802
rect 33070 34750 33122 34802
rect 36094 34750 36146 34802
rect 37102 34750 37154 34802
rect 37886 34750 37938 34802
rect 40126 34750 40178 34802
rect 41582 34750 41634 34802
rect 47742 34750 47794 34802
rect 49646 34750 49698 34802
rect 51550 34750 51602 34802
rect 52782 34750 52834 34802
rect 53006 34750 53058 34802
rect 53454 34750 53506 34802
rect 55470 34750 55522 34802
rect 57598 34750 57650 34802
rect 58046 34750 58098 34802
rect 8542 34638 8594 34690
rect 9886 34638 9938 34690
rect 12126 34638 12178 34690
rect 16606 34638 16658 34690
rect 19854 34638 19906 34690
rect 20302 34638 20354 34690
rect 22878 34638 22930 34690
rect 23774 34638 23826 34690
rect 27134 34638 27186 34690
rect 27582 34638 27634 34690
rect 30046 34638 30098 34690
rect 33406 34638 33458 34690
rect 34078 34638 34130 34690
rect 35198 34638 35250 34690
rect 37662 34638 37714 34690
rect 39454 34638 39506 34690
rect 42254 34638 42306 34690
rect 45054 34638 45106 34690
rect 48526 34638 48578 34690
rect 49758 34638 49810 34690
rect 50318 34638 50370 34690
rect 51326 34638 51378 34690
rect 51886 34638 51938 34690
rect 55806 34638 55858 34690
rect 57374 34638 57426 34690
rect 4622 34526 4674 34578
rect 4958 34526 5010 34578
rect 5742 34526 5794 34578
rect 8990 34526 9042 34578
rect 9326 34526 9378 34578
rect 10110 34526 10162 34578
rect 23102 34526 23154 34578
rect 23998 34526 24050 34578
rect 24222 34526 24274 34578
rect 25902 34526 25954 34578
rect 28590 34526 28642 34578
rect 32734 34526 32786 34578
rect 33182 34526 33234 34578
rect 40798 34526 40850 34578
rect 43486 34526 43538 34578
rect 50766 34526 50818 34578
rect 52894 34526 52946 34578
rect 9438 34414 9490 34466
rect 12910 34414 12962 34466
rect 19406 34414 19458 34466
rect 28030 34414 28082 34466
rect 50878 34414 50930 34466
rect 19838 34246 19890 34298
rect 19942 34246 19994 34298
rect 20046 34246 20098 34298
rect 50558 34246 50610 34298
rect 50662 34246 50714 34298
rect 50766 34246 50818 34298
rect 1822 34078 1874 34130
rect 2718 34078 2770 34130
rect 12126 34078 12178 34130
rect 12574 34078 12626 34130
rect 46622 34078 46674 34130
rect 50542 34078 50594 34130
rect 5518 33966 5570 34018
rect 15038 33966 15090 34018
rect 22654 33966 22706 34018
rect 25566 33966 25618 34018
rect 26798 33966 26850 34018
rect 28142 33966 28194 34018
rect 29486 33966 29538 34018
rect 36542 33966 36594 34018
rect 36990 33966 37042 34018
rect 37550 33966 37602 34018
rect 38782 33966 38834 34018
rect 39230 33966 39282 34018
rect 39678 33966 39730 34018
rect 40350 33966 40402 34018
rect 41022 33966 41074 34018
rect 41470 33966 41522 34018
rect 42366 33966 42418 34018
rect 53230 33966 53282 34018
rect 55022 33966 55074 34018
rect 55806 33966 55858 34018
rect 58158 33966 58210 34018
rect 10334 33854 10386 33906
rect 11006 33854 11058 33906
rect 13022 33854 13074 33906
rect 13582 33854 13634 33906
rect 13694 33854 13746 33906
rect 14142 33854 14194 33906
rect 14702 33854 14754 33906
rect 16158 33854 16210 33906
rect 18958 33854 19010 33906
rect 19070 33854 19122 33906
rect 25230 33854 25282 33906
rect 27134 33854 27186 33906
rect 34078 33854 34130 33906
rect 35870 33854 35922 33906
rect 36206 33854 36258 33906
rect 42814 33854 42866 33906
rect 43486 33854 43538 33906
rect 44270 33854 44322 33906
rect 45614 33854 45666 33906
rect 46286 33854 46338 33906
rect 47070 33854 47122 33906
rect 47518 33854 47570 33906
rect 49086 33854 49138 33906
rect 49646 33854 49698 33906
rect 52558 33854 52610 33906
rect 52894 33854 52946 33906
rect 54350 33854 54402 33906
rect 56926 33854 56978 33906
rect 57710 33854 57762 33906
rect 2718 33742 2770 33794
rect 3278 33742 3330 33794
rect 14478 33742 14530 33794
rect 15934 33742 15986 33794
rect 16382 33742 16434 33794
rect 18398 33742 18450 33794
rect 21982 33742 22034 33794
rect 27694 33742 27746 33794
rect 28702 33742 28754 33794
rect 32398 33742 32450 33794
rect 33518 33742 33570 33794
rect 34862 33742 34914 33794
rect 35198 33742 35250 33794
rect 43150 33742 43202 33794
rect 43822 33742 43874 33794
rect 44942 33742 44994 33794
rect 49422 33742 49474 33794
rect 50206 33742 50258 33794
rect 51102 33742 51154 33794
rect 51326 33742 51378 33794
rect 51774 33742 51826 33794
rect 52222 33742 52274 33794
rect 53790 33742 53842 33794
rect 56030 33742 56082 33794
rect 56702 33742 56754 33794
rect 1822 33630 1874 33682
rect 2382 33630 2434 33682
rect 5854 33630 5906 33682
rect 14366 33630 14418 33682
rect 21534 33630 21586 33682
rect 24670 33630 24722 33682
rect 26462 33630 26514 33682
rect 32062 33630 32114 33682
rect 34190 33630 34242 33682
rect 35534 33630 35586 33682
rect 41918 33630 41970 33682
rect 48190 33630 48242 33682
rect 57374 33630 57426 33682
rect 27918 33518 27970 33570
rect 31502 33518 31554 33570
rect 16046 33406 16098 33458
rect 17950 33406 18002 33458
rect 27246 33406 27298 33458
rect 32510 33406 32562 33458
rect 33070 33406 33122 33458
rect 48638 33406 48690 33458
rect 4478 33238 4530 33290
rect 4582 33238 4634 33290
rect 4686 33238 4738 33290
rect 35198 33238 35250 33290
rect 35302 33238 35354 33290
rect 35406 33238 35458 33290
rect 4846 33070 4898 33122
rect 34750 33070 34802 33122
rect 35198 33070 35250 33122
rect 40798 33070 40850 33122
rect 12462 32958 12514 33010
rect 14702 32958 14754 33010
rect 20414 32958 20466 33010
rect 46062 32958 46114 33010
rect 50654 32958 50706 33010
rect 51214 32958 51266 33010
rect 22430 32846 22482 32898
rect 28366 32846 28418 32898
rect 31950 32846 32002 32898
rect 34190 32846 34242 32898
rect 34750 32846 34802 32898
rect 35198 32846 35250 32898
rect 35758 32846 35810 32898
rect 37326 32846 37378 32898
rect 39118 32846 39170 32898
rect 43262 32846 43314 32898
rect 45614 32846 45666 32898
rect 50654 32846 50706 32898
rect 51102 32846 51154 32898
rect 56366 32846 56418 32898
rect 57710 32846 57762 32898
rect 58158 32846 58210 32898
rect 4510 32734 4562 32786
rect 11902 32734 11954 32786
rect 15150 32734 15202 32786
rect 15374 32734 15426 32786
rect 17278 32734 17330 32786
rect 17614 32734 17666 32786
rect 18510 32734 18562 32786
rect 23214 32734 23266 32786
rect 26014 32734 26066 32786
rect 27022 32734 27074 32786
rect 27246 32734 27298 32786
rect 27806 32734 27858 32786
rect 32174 32734 32226 32786
rect 33518 32734 33570 32786
rect 37886 32734 37938 32786
rect 38110 32734 38162 32786
rect 40238 32734 40290 32786
rect 42814 32734 42866 32786
rect 46622 32734 46674 32786
rect 48974 32734 49026 32786
rect 49310 32734 49362 32786
rect 53230 32734 53282 32786
rect 53566 32734 53618 32786
rect 53902 32734 53954 32786
rect 56702 32734 56754 32786
rect 57262 32734 57314 32786
rect 4398 32622 4450 32674
rect 12798 32622 12850 32674
rect 14142 32622 14194 32674
rect 15710 32622 15762 32674
rect 16942 32622 16994 32674
rect 19070 32622 19122 32674
rect 20750 32622 20802 32674
rect 23998 32622 24050 32674
rect 26350 32622 26402 32674
rect 26686 32622 26738 32674
rect 27582 32622 27634 32674
rect 32510 32622 32562 32674
rect 34078 32622 34130 32674
rect 40126 32622 40178 32674
rect 41918 32622 41970 32674
rect 46958 32622 47010 32674
rect 52894 32622 52946 32674
rect 54350 32622 54402 32674
rect 55022 32622 55074 32674
rect 55694 32622 55746 32674
rect 56814 32622 56866 32674
rect 57150 32622 57202 32674
rect 4958 32510 5010 32562
rect 14478 32510 14530 32562
rect 17950 32510 18002 32562
rect 19742 32510 19794 32562
rect 22766 32510 22818 32562
rect 22878 32510 22930 32562
rect 26798 32510 26850 32562
rect 31950 32510 32002 32562
rect 32846 32510 32898 32562
rect 43710 32510 43762 32562
rect 44158 32510 44210 32562
rect 45166 32510 45218 32562
rect 52110 32510 52162 32562
rect 56254 32510 56306 32562
rect 11790 32398 11842 32450
rect 27694 32398 27746 32450
rect 33070 32398 33122 32450
rect 38446 32398 38498 32450
rect 19838 32230 19890 32282
rect 19942 32230 19994 32282
rect 20046 32230 20098 32282
rect 50558 32230 50610 32282
rect 50662 32230 50714 32282
rect 50766 32230 50818 32282
rect 41246 32062 41298 32114
rect 5518 31950 5570 32002
rect 13470 31950 13522 32002
rect 19742 31950 19794 32002
rect 22878 31950 22930 32002
rect 23662 31950 23714 32002
rect 27918 31950 27970 32002
rect 28366 31950 28418 32002
rect 32174 31950 32226 32002
rect 44382 31950 44434 32002
rect 51550 31950 51602 32002
rect 52894 31950 52946 32002
rect 2382 31838 2434 31890
rect 5854 31838 5906 31890
rect 14366 31838 14418 31890
rect 15934 31838 15986 31890
rect 16046 31838 16098 31890
rect 20974 31838 21026 31890
rect 21086 31838 21138 31890
rect 21870 31838 21922 31890
rect 22542 31838 22594 31890
rect 23886 31838 23938 31890
rect 24110 31838 24162 31890
rect 25342 31838 25394 31890
rect 25566 31838 25618 31890
rect 25902 31838 25954 31890
rect 26238 31838 26290 31890
rect 26350 31838 26402 31890
rect 2718 31726 2770 31778
rect 3278 31726 3330 31778
rect 10782 31726 10834 31778
rect 11342 31726 11394 31778
rect 13918 31726 13970 31778
rect 14478 31726 14530 31778
rect 15374 31726 15426 31778
rect 20414 31726 20466 31778
rect 20862 31726 20914 31778
rect 21310 31732 21362 31784
rect 27022 31782 27074 31834
rect 27582 31838 27634 31890
rect 31278 31838 31330 31890
rect 31838 31838 31890 31890
rect 32510 31838 32562 31890
rect 33294 31838 33346 31890
rect 35758 31838 35810 31890
rect 37774 31838 37826 31890
rect 38446 31838 38498 31890
rect 39118 31838 39170 31890
rect 41694 31838 41746 31890
rect 42814 31838 42866 31890
rect 43374 31838 43426 31890
rect 44046 31838 44098 31890
rect 45390 31838 45442 31890
rect 46622 31838 46674 31890
rect 47182 31838 47234 31890
rect 51998 31838 52050 31890
rect 53342 31838 53394 31890
rect 21758 31726 21810 31778
rect 23214 31726 23266 31778
rect 24334 31726 24386 31778
rect 25230 31726 25282 31778
rect 27246 31726 27298 31778
rect 31614 31726 31666 31778
rect 33070 31726 33122 31778
rect 33518 31738 33570 31790
rect 34414 31726 34466 31778
rect 34750 31726 34802 31778
rect 36318 31726 36370 31778
rect 36654 31726 36706 31778
rect 36990 31726 37042 31778
rect 37326 31726 37378 31778
rect 40910 31726 40962 31778
rect 43486 31726 43538 31778
rect 46398 31726 46450 31778
rect 47966 31726 48018 31778
rect 49870 31726 49922 31778
rect 53454 31726 53506 31778
rect 55022 31753 55074 31805
rect 10446 31614 10498 31666
rect 14926 31614 14978 31666
rect 16830 31614 16882 31666
rect 23662 31614 23714 31666
rect 24558 31614 24610 31666
rect 30830 31614 30882 31666
rect 39902 31614 39954 31666
rect 40350 31614 40402 31666
rect 45390 31614 45442 31666
rect 46846 31614 46898 31666
rect 47518 31614 47570 31666
rect 49534 31614 49586 31666
rect 50206 31614 50258 31666
rect 51102 31614 51154 31666
rect 52446 31614 52498 31666
rect 55806 31614 55858 31666
rect 56702 31614 56754 31666
rect 57150 31614 57202 31666
rect 17726 31502 17778 31554
rect 25790 31502 25842 31554
rect 31502 31502 31554 31554
rect 45726 31502 45778 31554
rect 26910 31390 26962 31442
rect 33406 31390 33458 31442
rect 42478 31390 42530 31442
rect 4478 31222 4530 31274
rect 4582 31222 4634 31274
rect 4686 31222 4738 31274
rect 35198 31222 35250 31274
rect 35302 31222 35354 31274
rect 35406 31222 35458 31274
rect 17278 31054 17330 31106
rect 18734 31054 18786 31106
rect 23886 31054 23938 31106
rect 25118 31054 25170 31106
rect 27582 31054 27634 31106
rect 32958 31054 33010 31106
rect 15038 30942 15090 30994
rect 26126 30942 26178 30994
rect 5630 30830 5682 30882
rect 16158 30830 16210 30882
rect 28254 30830 28306 30882
rect 31166 30830 31218 30882
rect 32286 30830 32338 30882
rect 32734 30830 32786 30882
rect 32846 30830 32898 30882
rect 36318 30942 36370 30994
rect 33518 30830 33570 30882
rect 33854 30830 33906 30882
rect 35534 30830 35586 30882
rect 40574 30830 40626 30882
rect 43598 30830 43650 30882
rect 44046 30830 44098 30882
rect 45614 30830 45666 30882
rect 46398 30830 46450 30882
rect 53678 30830 53730 30882
rect 55582 30830 55634 30882
rect 1822 30718 1874 30770
rect 2382 30718 2434 30770
rect 9662 30718 9714 30770
rect 10222 30718 10274 30770
rect 14590 30718 14642 30770
rect 17950 30718 18002 30770
rect 19182 30718 19234 30770
rect 19406 30718 19458 30770
rect 23550 30718 23602 30770
rect 23774 30718 23826 30770
rect 23998 30718 24050 30770
rect 24222 30718 24274 30770
rect 24558 30718 24610 30770
rect 24782 30718 24834 30770
rect 26462 30718 26514 30770
rect 27358 30718 27410 30770
rect 27918 30718 27970 30770
rect 28590 30718 28642 30770
rect 30718 30718 30770 30770
rect 32734 30718 32786 30770
rect 33182 30718 33234 30770
rect 33518 30718 33570 30770
rect 33966 30718 34018 30770
rect 35646 30718 35698 30770
rect 37662 30718 37714 30770
rect 39678 30718 39730 30770
rect 41134 30718 41186 30770
rect 41358 30718 41410 30770
rect 41806 30718 41858 30770
rect 44942 30718 44994 30770
rect 45166 30718 45218 30770
rect 45390 30718 45442 30770
rect 45950 30718 46002 30770
rect 46174 30718 46226 30770
rect 14030 30606 14082 30658
rect 14478 30606 14530 30658
rect 15486 30606 15538 30658
rect 16046 30606 16098 30658
rect 17726 30606 17778 30658
rect 18286 30606 18338 30658
rect 19630 30606 19682 30658
rect 22766 30606 22818 30658
rect 25006 30606 25058 30658
rect 25566 30606 25618 30658
rect 25678 30606 25730 30658
rect 26350 30606 26402 30658
rect 26910 30606 26962 30658
rect 27022 30606 27074 30658
rect 27694 30606 27746 30658
rect 28366 30606 28418 30658
rect 30830 30606 30882 30658
rect 31390 30606 31442 30658
rect 32062 30606 32114 30658
rect 32958 30606 33010 30658
rect 33742 30606 33794 30658
rect 34414 30606 34466 30658
rect 36990 30606 37042 30658
rect 39230 30606 39282 30658
rect 45614 30606 45666 30658
rect 46622 30606 46674 30658
rect 49310 30606 49362 30658
rect 53006 30606 53058 30658
rect 53566 30606 53618 30658
rect 54238 30606 54290 30658
rect 54686 30606 54738 30658
rect 4622 30494 4674 30546
rect 4958 30494 5010 30546
rect 5742 30494 5794 30546
rect 6078 30494 6130 30546
rect 9326 30494 9378 30546
rect 12462 30494 12514 30546
rect 12798 30494 12850 30546
rect 23102 30494 23154 30546
rect 26014 30494 26066 30546
rect 26686 30494 26738 30546
rect 29262 30494 29314 30546
rect 29710 30494 29762 30546
rect 31726 30494 31778 30546
rect 34750 30494 34802 30546
rect 37326 30494 37378 30546
rect 39118 30494 39170 30546
rect 43150 30494 43202 30546
rect 45054 30494 45106 30546
rect 47070 30494 47122 30546
rect 48302 30494 48354 30546
rect 48750 30494 48802 30546
rect 49982 30494 50034 30546
rect 55134 30494 55186 30546
rect 56030 30494 56082 30546
rect 6190 30382 6242 30434
rect 13582 30382 13634 30434
rect 31054 30382 31106 30434
rect 37998 30382 38050 30434
rect 51886 30382 51938 30434
rect 52558 30382 52610 30434
rect 54910 30382 54962 30434
rect 55806 30382 55858 30434
rect 19838 30214 19890 30266
rect 19942 30214 19994 30266
rect 20046 30214 20098 30266
rect 50558 30214 50610 30266
rect 50662 30214 50714 30266
rect 50766 30214 50818 30266
rect 3838 30046 3890 30098
rect 10334 30046 10386 30098
rect 14254 30046 14306 30098
rect 24446 30046 24498 30098
rect 25566 30046 25618 30098
rect 26462 30046 26514 30098
rect 28142 30046 28194 30098
rect 48638 30046 48690 30098
rect 50542 30046 50594 30098
rect 51102 30046 51154 30098
rect 4734 29934 4786 29986
rect 5182 29934 5234 29986
rect 8542 29934 8594 29986
rect 13470 29934 13522 29986
rect 13918 29934 13970 29986
rect 24334 29934 24386 29986
rect 27806 29934 27858 29986
rect 30158 29934 30210 29986
rect 31726 29934 31778 29986
rect 32174 29934 32226 29986
rect 34190 29934 34242 29986
rect 36654 29934 36706 29986
rect 37998 29934 38050 29986
rect 38446 29934 38498 29986
rect 38894 29934 38946 29986
rect 39902 29934 39954 29986
rect 40350 29934 40402 29986
rect 43374 29934 43426 29986
rect 45166 29934 45218 29986
rect 46398 29934 46450 29986
rect 15262 29822 15314 29874
rect 23886 29822 23938 29874
rect 24222 29822 24274 29874
rect 24782 29822 24834 29874
rect 25230 29822 25282 29874
rect 25566 29822 25618 29874
rect 25678 29822 25730 29874
rect 26574 29822 26626 29874
rect 26910 29822 26962 29874
rect 27022 29822 27074 29874
rect 27470 29822 27522 29874
rect 29598 29822 29650 29874
rect 30494 29822 30546 29874
rect 31054 29822 31106 29874
rect 31390 29822 31442 29874
rect 32510 29822 32562 29874
rect 34526 29822 34578 29874
rect 35758 29822 35810 29874
rect 36206 29822 36258 29874
rect 41246 29822 41298 29874
rect 41694 29822 41746 29874
rect 42366 29822 42418 29874
rect 42702 29822 42754 29874
rect 43038 29822 43090 29874
rect 43822 29822 43874 29874
rect 49646 29822 49698 29874
rect 51326 29822 51378 29874
rect 51662 29822 51714 29874
rect 51998 29822 52050 29874
rect 52782 29822 52834 29874
rect 54126 29822 54178 29874
rect 3390 29710 3442 29762
rect 3726 29710 3778 29762
rect 4174 29710 4226 29762
rect 7310 29710 7362 29762
rect 7870 29710 7922 29762
rect 8990 29710 9042 29762
rect 9998 29710 10050 29762
rect 10446 29710 10498 29762
rect 10782 29710 10834 29762
rect 11342 29710 11394 29762
rect 14702 29710 14754 29762
rect 14926 29710 14978 29762
rect 26126 29710 26178 29762
rect 26238 29710 26290 29762
rect 28478 29710 28530 29762
rect 29262 29710 29314 29762
rect 29934 29710 29986 29762
rect 33070 29710 33122 29762
rect 33182 29710 33234 29762
rect 33294 29710 33346 29762
rect 33518 29710 33570 29762
rect 33742 29710 33794 29762
rect 34862 29710 34914 29762
rect 35422 29710 35474 29762
rect 35534 29710 35586 29762
rect 41470 29710 41522 29762
rect 44494 29710 44546 29762
rect 49086 29710 49138 29762
rect 49310 29710 49362 29762
rect 52334 29710 52386 29762
rect 53454 29710 53506 29762
rect 1822 29598 1874 29650
rect 2942 29598 2994 29650
rect 28926 29598 28978 29650
rect 29598 29598 29650 29650
rect 37102 29598 37154 29650
rect 37550 29598 37602 29650
rect 39454 29598 39506 29650
rect 45950 29598 46002 29650
rect 48190 29598 48242 29650
rect 50542 29598 50594 29650
rect 50990 29598 51042 29650
rect 54910 29598 54962 29650
rect 55806 29598 55858 29650
rect 35198 29486 35250 29538
rect 3278 29374 3330 29426
rect 4286 29374 4338 29426
rect 8878 29374 8930 29426
rect 9886 29374 9938 29426
rect 40798 29374 40850 29426
rect 4478 29206 4530 29258
rect 4582 29206 4634 29258
rect 4686 29206 4738 29258
rect 35198 29206 35250 29258
rect 35302 29206 35354 29258
rect 35406 29206 35458 29258
rect 13470 29038 13522 29090
rect 27134 29038 27186 29090
rect 27694 29038 27746 29090
rect 40126 29038 40178 29090
rect 50878 29038 50930 29090
rect 54014 29038 54066 29090
rect 1934 28926 1986 28978
rect 8766 28926 8818 28978
rect 12798 28926 12850 28978
rect 35646 28926 35698 28978
rect 36430 28926 36482 28978
rect 9326 28814 9378 28866
rect 15150 28814 15202 28866
rect 24782 28814 24834 28866
rect 25230 28814 25282 28866
rect 26014 28814 26066 28866
rect 27582 28814 27634 28866
rect 31502 28814 31554 28866
rect 35198 28814 35250 28866
rect 35646 28814 35698 28866
rect 36094 28814 36146 28866
rect 37102 28814 37154 28866
rect 39118 28814 39170 28866
rect 39902 28814 39954 28866
rect 41246 28814 41298 28866
rect 43374 28814 43426 28866
rect 43822 28814 43874 28866
rect 44270 28814 44322 28866
rect 46174 28814 46226 28866
rect 49870 28814 49922 28866
rect 54014 28814 54066 28866
rect 4510 28702 4562 28754
rect 5070 28702 5122 28754
rect 5630 28702 5682 28754
rect 6190 28702 6242 28754
rect 9662 28702 9714 28754
rect 10222 28702 10274 28754
rect 13582 28702 13634 28754
rect 14030 28702 14082 28754
rect 14478 28702 14530 28754
rect 20302 28702 20354 28754
rect 21310 28702 21362 28754
rect 22318 28702 22370 28754
rect 24446 28702 24498 28754
rect 25118 28702 25170 28754
rect 26350 28702 26402 28754
rect 29486 28702 29538 28754
rect 29710 28702 29762 28754
rect 30158 28702 30210 28754
rect 30382 28702 30434 28754
rect 30606 28702 30658 28754
rect 31054 28702 31106 28754
rect 32062 28702 32114 28754
rect 32510 28702 32562 28754
rect 32846 28702 32898 28754
rect 32958 28702 33010 28754
rect 33070 28702 33122 28754
rect 33294 28702 33346 28754
rect 33518 28702 33570 28754
rect 33966 28702 34018 28754
rect 34190 28702 34242 28754
rect 34414 28702 34466 28754
rect 34638 28702 34690 28754
rect 40574 28702 40626 28754
rect 46846 28702 46898 28754
rect 49086 28702 49138 28754
rect 51550 28702 51602 28754
rect 55134 28702 55186 28754
rect 56926 28702 56978 28754
rect 15038 28590 15090 28642
rect 20750 28590 20802 28642
rect 25454 28590 25506 28642
rect 25678 28590 25730 28642
rect 27134 28590 27186 28642
rect 29822 28590 29874 28642
rect 30718 28590 30770 28642
rect 31278 28590 31330 28642
rect 34078 28590 34130 28642
rect 38782 28590 38834 28642
rect 41022 28590 41074 28642
rect 44830 28590 44882 28642
rect 48190 28590 48242 28642
rect 51326 28590 51378 28642
rect 51886 28590 51938 28642
rect 52782 28590 52834 28642
rect 54238 28590 54290 28642
rect 57038 28590 57090 28642
rect 2382 28478 2434 28530
rect 8430 28478 8482 28530
rect 12462 28478 12514 28530
rect 21646 28478 21698 28530
rect 22766 28478 22818 28530
rect 24558 28478 24610 28530
rect 25006 28478 25058 28530
rect 25902 28478 25954 28530
rect 26798 28478 26850 28530
rect 31502 28478 31554 28530
rect 32398 28478 32450 28530
rect 45166 28478 45218 28530
rect 50654 28478 50706 28530
rect 25790 28366 25842 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 5630 28030 5682 28082
rect 6302 28030 6354 28082
rect 22654 28030 22706 28082
rect 33406 28030 33458 28082
rect 35534 28030 35586 28082
rect 38446 28030 38498 28082
rect 39454 28030 39506 28082
rect 49758 28030 49810 28082
rect 3838 27918 3890 27970
rect 4286 27918 4338 27970
rect 8990 27918 9042 27970
rect 12462 27918 12514 27970
rect 12798 27918 12850 27970
rect 22990 27918 23042 27970
rect 23438 27918 23490 27970
rect 25230 27918 25282 27970
rect 26686 27918 26738 27970
rect 27470 27918 27522 27970
rect 29710 27918 29762 27970
rect 30830 27918 30882 27970
rect 31838 27918 31890 27970
rect 34526 27918 34578 27970
rect 35198 27918 35250 27970
rect 38558 27918 38610 27970
rect 39454 27918 39506 27970
rect 45166 27918 45218 27970
rect 45614 27918 45666 27970
rect 51550 27918 51602 27970
rect 53118 27918 53170 27970
rect 57710 27918 57762 27970
rect 1822 27806 1874 27858
rect 3390 27806 3442 27858
rect 21646 27806 21698 27858
rect 25566 27806 25618 27858
rect 26126 27806 26178 27858
rect 27022 27806 27074 27858
rect 32174 27806 32226 27858
rect 33406 27806 33458 27858
rect 33518 27806 33570 27858
rect 33854 27806 33906 27858
rect 34190 27806 34242 27858
rect 46622 27806 46674 27858
rect 48302 27806 48354 27858
rect 48750 27806 48802 27858
rect 49422 27806 49474 27858
rect 52110 27806 52162 27858
rect 53566 27806 53618 27858
rect 54910 27806 54962 27858
rect 56702 27806 56754 27858
rect 56926 27806 56978 27858
rect 57150 27806 57202 27858
rect 6414 27694 6466 27746
rect 6974 27694 7026 27746
rect 9662 27694 9714 27746
rect 10222 27694 10274 27746
rect 17390 27694 17442 27746
rect 19518 27694 19570 27746
rect 20862 27694 20914 27746
rect 21758 27694 21810 27746
rect 22206 27694 22258 27746
rect 23998 27694 24050 27746
rect 24222 27694 24274 27746
rect 24446 27694 24498 27746
rect 24670 27694 24722 27746
rect 26350 27694 26402 27746
rect 29598 27694 29650 27746
rect 29822 27694 29874 27746
rect 30046 27694 30098 27746
rect 30270 27694 30322 27746
rect 30718 27694 30770 27746
rect 30942 27694 30994 27746
rect 31166 27694 31218 27746
rect 31390 27694 31442 27746
rect 33070 27694 33122 27746
rect 35086 27694 35138 27746
rect 35310 27694 35362 27746
rect 35646 27694 35698 27746
rect 35870 27694 35922 27746
rect 41806 27694 41858 27746
rect 42142 27694 42194 27746
rect 50318 27694 50370 27746
rect 50542 27694 50594 27746
rect 51214 27694 51266 27746
rect 51550 27694 51602 27746
rect 52446 27694 52498 27746
rect 52782 27694 52834 27746
rect 54238 27694 54290 27746
rect 55694 27694 55746 27746
rect 56590 27694 56642 27746
rect 57262 27694 57314 27746
rect 58158 27694 58210 27746
rect 17726 27582 17778 27634
rect 26014 27582 26066 27634
rect 39006 27582 39058 27634
rect 40350 27582 40402 27634
rect 41022 27582 41074 27634
rect 46062 27582 46114 27634
rect 47742 27582 47794 27634
rect 23886 27470 23938 27522
rect 46958 27470 47010 27522
rect 49086 27470 49138 27522
rect 22878 27358 22930 27410
rect 34526 27358 34578 27410
rect 34750 27358 34802 27410
rect 42702 27358 42754 27410
rect 4478 27190 4530 27242
rect 4582 27190 4634 27242
rect 4686 27190 4738 27242
rect 35198 27190 35250 27242
rect 35302 27190 35354 27242
rect 35406 27190 35458 27242
rect 30718 27022 30770 27074
rect 48862 27022 48914 27074
rect 49422 27022 49474 27074
rect 50094 27022 50146 27074
rect 23886 26910 23938 26962
rect 33182 26910 33234 26962
rect 5742 26798 5794 26850
rect 22542 26798 22594 26850
rect 25118 26798 25170 26850
rect 26126 26798 26178 26850
rect 27022 26798 27074 26850
rect 33742 26798 33794 26850
rect 34078 26798 34130 26850
rect 34862 26798 34914 26850
rect 37102 26798 37154 26850
rect 42030 26798 42082 26850
rect 15934 26686 15986 26738
rect 21870 26686 21922 26738
rect 23774 26686 23826 26738
rect 24446 26686 24498 26738
rect 24670 26686 24722 26738
rect 25566 26686 25618 26738
rect 25678 26686 25730 26738
rect 26574 26686 26626 26738
rect 29934 26686 29986 26738
rect 30158 26686 30210 26738
rect 30382 26686 30434 26738
rect 30606 26686 30658 26738
rect 31166 26686 31218 26738
rect 31502 26686 31554 26738
rect 31726 26686 31778 26738
rect 32286 26686 32338 26738
rect 32510 26686 32562 26738
rect 32846 26686 32898 26738
rect 33966 26686 34018 26738
rect 34974 26686 35026 26738
rect 39454 26686 39506 26738
rect 42702 26686 42754 26738
rect 42926 26686 42978 26738
rect 48862 26686 48914 26738
rect 50094 26686 50146 26738
rect 50766 26686 50818 26738
rect 50990 26686 51042 26738
rect 51214 26686 51266 26738
rect 51662 26686 51714 26738
rect 51886 26686 51938 26738
rect 53566 26686 53618 26738
rect 54126 26686 54178 26738
rect 55806 26686 55858 26738
rect 57262 26686 57314 26738
rect 16382 26574 16434 26626
rect 16942 26574 16994 26626
rect 17054 26574 17106 26626
rect 17726 26574 17778 26626
rect 17838 26574 17890 26626
rect 19854 26574 19906 26626
rect 21646 26574 21698 26626
rect 22094 26574 22146 26626
rect 23550 26574 23602 26626
rect 24222 26574 24274 26626
rect 25006 26574 25058 26626
rect 25230 26574 25282 26626
rect 26350 26574 26402 26626
rect 33518 26574 33570 26626
rect 34190 26574 34242 26626
rect 34302 26574 34354 26626
rect 34750 26574 34802 26626
rect 34974 26574 35026 26626
rect 35534 26574 35586 26626
rect 38446 26574 38498 26626
rect 38782 26574 38834 26626
rect 39118 26574 39170 26626
rect 39902 26574 39954 26626
rect 40574 26574 40626 26626
rect 43150 26574 43202 26626
rect 51438 26574 51490 26626
rect 56926 26574 56978 26626
rect 20750 26462 20802 26514
rect 23326 26462 23378 26514
rect 25902 26462 25954 26514
rect 27358 26462 27410 26514
rect 28590 26462 28642 26514
rect 29598 26462 29650 26514
rect 32062 26462 32114 26514
rect 33854 26462 33906 26514
rect 35198 26462 35250 26514
rect 35870 26462 35922 26514
rect 35982 26462 36034 26514
rect 36430 26462 36482 26514
rect 37550 26462 37602 26514
rect 37998 26462 38050 26514
rect 41246 26462 41298 26514
rect 43934 26462 43986 26514
rect 45502 26462 45554 26514
rect 49310 26462 49362 26514
rect 49758 26462 49810 26514
rect 51998 26462 52050 26514
rect 52782 26462 52834 26514
rect 54350 26462 54402 26514
rect 24334 26350 24386 26402
rect 35086 26350 35138 26402
rect 36990 26350 37042 26402
rect 38110 26350 38162 26402
rect 42254 26350 42306 26402
rect 48526 26350 48578 26402
rect 50430 26350 50482 26402
rect 19838 26182 19890 26234
rect 19942 26182 19994 26234
rect 20046 26182 20098 26234
rect 50558 26182 50610 26234
rect 50662 26182 50714 26234
rect 50766 26182 50818 26234
rect 22766 26014 22818 26066
rect 41134 26014 41186 26066
rect 43150 26014 43202 26066
rect 45838 26014 45890 26066
rect 49758 26014 49810 26066
rect 50990 26014 51042 26066
rect 52110 26014 52162 26066
rect 52670 26014 52722 26066
rect 16718 25902 16770 25954
rect 20526 25902 20578 25954
rect 25230 25902 25282 25954
rect 26014 25902 26066 25954
rect 26910 25902 26962 25954
rect 28478 25902 28530 25954
rect 29374 25902 29426 25954
rect 32510 25902 32562 25954
rect 33182 25902 33234 25954
rect 34414 25902 34466 25954
rect 36542 25902 36594 25954
rect 36990 25902 37042 25954
rect 49310 25902 49362 25954
rect 49758 25902 49810 25954
rect 51550 25902 51602 25954
rect 52110 25902 52162 25954
rect 53342 25902 53394 25954
rect 55022 25902 55074 25954
rect 55358 25902 55410 25954
rect 17614 25790 17666 25842
rect 18174 25790 18226 25842
rect 21870 25790 21922 25842
rect 23438 25790 23490 25842
rect 24446 25790 24498 25842
rect 25566 25790 25618 25842
rect 26126 25790 26178 25842
rect 27022 25790 27074 25842
rect 29710 25790 29762 25842
rect 30830 25790 30882 25842
rect 31390 25790 31442 25842
rect 31614 25790 31666 25842
rect 35422 25790 35474 25842
rect 41246 25790 41298 25842
rect 46846 25790 46898 25842
rect 54014 25790 54066 25842
rect 13470 25678 13522 25730
rect 17950 25678 18002 25730
rect 22430 25678 22482 25730
rect 23102 25678 23154 25730
rect 23886 25678 23938 25730
rect 25902 25678 25954 25730
rect 26350 25678 26402 25730
rect 26798 25678 26850 25730
rect 27246 25678 27298 25730
rect 30270 25678 30322 25730
rect 30494 25678 30546 25730
rect 30606 25678 30658 25730
rect 31726 25678 31778 25730
rect 31950 25678 32002 25730
rect 32174 25678 32226 25730
rect 33630 25678 33682 25730
rect 35870 25678 35922 25730
rect 36206 25678 36258 25730
rect 37550 25678 37602 25730
rect 37774 25678 37826 25730
rect 37886 25678 37938 25730
rect 38110 25678 38162 25730
rect 39118 25678 39170 25730
rect 39342 25678 39394 25730
rect 39678 25678 39730 25730
rect 41022 25678 41074 25730
rect 44830 25678 44882 25730
rect 46286 25678 46338 25730
rect 46510 25678 46562 25730
rect 54462 25678 54514 25730
rect 18958 25566 19010 25618
rect 20974 25566 21026 25618
rect 21422 25566 21474 25618
rect 24558 25566 24610 25618
rect 28030 25566 28082 25618
rect 28926 25566 28978 25618
rect 29934 25566 29986 25618
rect 31166 25566 31218 25618
rect 34974 25566 35026 25618
rect 35646 25566 35698 25618
rect 38558 25566 38610 25618
rect 50206 25566 50258 25618
rect 50654 25566 50706 25618
rect 51102 25566 51154 25618
rect 52558 25566 52610 25618
rect 55582 25566 55634 25618
rect 56030 25566 56082 25618
rect 56702 25566 56754 25618
rect 57150 25566 57202 25618
rect 57598 25566 57650 25618
rect 30158 25454 30210 25506
rect 49870 25454 49922 25506
rect 50654 25454 50706 25506
rect 56702 25454 56754 25506
rect 57598 25454 57650 25506
rect 18622 25342 18674 25394
rect 50430 25342 50482 25394
rect 51102 25342 51154 25394
rect 51326 25342 51378 25394
rect 51662 25342 51714 25394
rect 52558 25342 52610 25394
rect 4478 25174 4530 25226
rect 4582 25174 4634 25226
rect 4686 25174 4738 25226
rect 35198 25174 35250 25226
rect 35302 25174 35354 25226
rect 35406 25174 35458 25226
rect 24894 25006 24946 25058
rect 26798 25006 26850 25058
rect 47406 25006 47458 25058
rect 49198 25006 49250 25058
rect 50094 25006 50146 25058
rect 29934 24894 29986 24946
rect 30830 24894 30882 24946
rect 31390 24894 31442 24946
rect 34974 24894 35026 24946
rect 50206 24894 50258 24946
rect 16942 24782 16994 24834
rect 19182 24782 19234 24834
rect 20302 24782 20354 24834
rect 21646 24782 21698 24834
rect 22094 24782 22146 24834
rect 22878 24782 22930 24834
rect 27918 24782 27970 24834
rect 28590 24782 28642 24834
rect 36430 24782 36482 24834
rect 45726 24782 45778 24834
rect 13470 24670 13522 24722
rect 22430 24670 22482 24722
rect 23214 24670 23266 24722
rect 23326 24670 23378 24722
rect 24110 24670 24162 24722
rect 24670 24670 24722 24722
rect 25566 24670 25618 24722
rect 26462 24670 26514 24722
rect 26910 24670 26962 24722
rect 29374 24670 29426 24722
rect 32734 24670 32786 24722
rect 37998 24670 38050 24722
rect 38670 24670 38722 24722
rect 39790 24670 39842 24722
rect 40350 24670 40402 24722
rect 48414 24670 48466 24722
rect 50990 24670 51042 24722
rect 53454 24670 53506 24722
rect 53790 24670 53842 24722
rect 55246 24670 55298 24722
rect 57150 24670 57202 24722
rect 23886 24558 23938 24610
rect 24334 24558 24386 24610
rect 24558 24558 24610 24610
rect 25342 24558 25394 24610
rect 25790 24558 25842 24610
rect 26686 24558 26738 24610
rect 27470 24558 27522 24610
rect 29598 24558 29650 24610
rect 30270 24558 30322 24610
rect 30494 24558 30546 24610
rect 31054 24558 31106 24610
rect 31278 24558 31330 24610
rect 31838 24558 31890 24610
rect 31950 24558 32002 24610
rect 32846 24558 32898 24610
rect 33182 24558 33234 24610
rect 33518 24558 33570 24610
rect 38894 24558 38946 24610
rect 42366 24558 42418 24610
rect 43598 24558 43650 24610
rect 47854 24558 47906 24610
rect 48302 24558 48354 24610
rect 50654 24558 50706 24610
rect 51214 24558 51266 24610
rect 53118 24558 53170 24610
rect 54574 24558 54626 24610
rect 56814 24558 56866 24610
rect 19854 24446 19906 24498
rect 20750 24446 20802 24498
rect 22542 24446 22594 24498
rect 22878 24446 22930 24498
rect 23550 24446 23602 24498
rect 29822 24446 29874 24498
rect 30606 24446 30658 24498
rect 31502 24446 31554 24498
rect 35534 24446 35586 24498
rect 35982 24446 36034 24498
rect 37326 24446 37378 24498
rect 49086 24446 49138 24498
rect 49534 24446 49586 24498
rect 49982 24446 50034 24498
rect 52110 24446 52162 24498
rect 52782 24446 52834 24498
rect 54126 24446 54178 24498
rect 55918 24446 55970 24498
rect 56702 24446 56754 24498
rect 57822 24446 57874 24498
rect 19854 24334 19906 24386
rect 20750 24334 20802 24386
rect 41470 24334 41522 24386
rect 49086 24334 49138 24386
rect 49982 24334 50034 24386
rect 19838 24166 19890 24218
rect 19942 24166 19994 24218
rect 20046 24166 20098 24218
rect 50558 24166 50610 24218
rect 50662 24166 50714 24218
rect 50766 24166 50818 24218
rect 26350 23998 26402 24050
rect 30606 23998 30658 24050
rect 49982 23998 50034 24050
rect 50654 23998 50706 24050
rect 56702 23998 56754 24050
rect 57486 23998 57538 24050
rect 21086 23886 21138 23938
rect 21758 23886 21810 23938
rect 24110 23886 24162 23938
rect 24558 23886 24610 23938
rect 26462 23886 26514 23938
rect 27246 23886 27298 23938
rect 31390 23886 31442 23938
rect 33742 23886 33794 23938
rect 38222 23886 38274 23938
rect 44830 23886 44882 23938
rect 45278 23886 45330 23938
rect 47518 23886 47570 23938
rect 49982 23886 50034 23938
rect 55694 23886 55746 23938
rect 56702 23886 56754 23938
rect 14590 23774 14642 23826
rect 19182 23774 19234 23826
rect 19406 23774 19458 23826
rect 23102 23774 23154 23826
rect 25454 23774 25506 23826
rect 25790 23774 25842 23826
rect 27470 23774 27522 23826
rect 27582 23774 27634 23826
rect 34190 23774 34242 23826
rect 37214 23774 37266 23826
rect 37550 23774 37602 23826
rect 38782 23774 38834 23826
rect 40014 23774 40066 23826
rect 42814 23774 42866 23826
rect 45726 23774 45778 23826
rect 47070 23774 47122 23826
rect 47742 23774 47794 23826
rect 48750 23774 48802 23826
rect 52334 23774 52386 23826
rect 53230 23774 53282 23826
rect 11678 23662 11730 23714
rect 17502 23662 17554 23714
rect 18846 23662 18898 23714
rect 22654 23662 22706 23714
rect 23550 23662 23602 23714
rect 26686 23662 26738 23714
rect 29486 23662 29538 23714
rect 31726 23662 31778 23714
rect 31950 23662 32002 23714
rect 32398 23662 32450 23714
rect 33070 23662 33122 23714
rect 33406 23662 33458 23714
rect 37886 23662 37938 23714
rect 39342 23662 39394 23714
rect 41134 23662 41186 23714
rect 41358 23662 41410 23714
rect 41470 23662 41522 23714
rect 51662 23662 51714 23714
rect 51774 23662 51826 23714
rect 54574 23662 54626 23714
rect 54686 23662 54738 23714
rect 34638 23550 34690 23602
rect 36430 23550 36482 23602
rect 36878 23550 36930 23602
rect 41918 23550 41970 23602
rect 48638 23550 48690 23602
rect 48974 23550 49026 23602
rect 50430 23550 50482 23602
rect 51214 23550 51266 23602
rect 57150 23550 57202 23602
rect 57598 23550 57650 23602
rect 24670 23438 24722 23490
rect 40798 23438 40850 23490
rect 49534 23438 49586 23490
rect 57150 23438 57202 23490
rect 57598 23438 57650 23490
rect 46622 23326 46674 23378
rect 4478 23158 4530 23210
rect 4582 23158 4634 23210
rect 4686 23158 4738 23210
rect 35198 23158 35250 23210
rect 35302 23158 35354 23210
rect 35406 23158 35458 23210
rect 16606 22990 16658 23042
rect 25902 22990 25954 23042
rect 37326 22990 37378 23042
rect 40126 22990 40178 23042
rect 41358 22990 41410 23042
rect 41806 22990 41858 23042
rect 50878 22990 50930 23042
rect 17614 22766 17666 22818
rect 19406 22766 19458 22818
rect 19854 22766 19906 22818
rect 20302 22766 20354 22818
rect 20750 22766 20802 22818
rect 21646 22766 21698 22818
rect 22094 22766 22146 22818
rect 22542 22766 22594 22818
rect 33966 22766 34018 22818
rect 36206 22766 36258 22818
rect 38894 22766 38946 22818
rect 40910 22766 40962 22818
rect 41918 22878 41970 22930
rect 41358 22766 41410 22818
rect 41806 22766 41858 22818
rect 42254 22766 42306 22818
rect 42702 22766 42754 22818
rect 52782 22766 52834 22818
rect 58158 22766 58210 22818
rect 15150 22654 15202 22706
rect 24670 22654 24722 22706
rect 25678 22654 25730 22706
rect 26350 22654 26402 22706
rect 26798 22654 26850 22706
rect 29262 22654 29314 22706
rect 29486 22654 29538 22706
rect 30046 22654 30098 22706
rect 30718 22654 30770 22706
rect 30942 22654 30994 22706
rect 31278 22654 31330 22706
rect 31390 22654 31442 22706
rect 37886 22654 37938 22706
rect 40462 22654 40514 22706
rect 40686 22654 40738 22706
rect 40910 22654 40962 22706
rect 46622 22654 46674 22706
rect 46958 22654 47010 22706
rect 47630 22654 47682 22706
rect 48190 22654 48242 22706
rect 51550 22654 51602 22706
rect 54014 22654 54066 22706
rect 55806 22654 55858 22706
rect 57486 22654 57538 22706
rect 57710 22654 57762 22706
rect 24334 22542 24386 22594
rect 25566 22542 25618 22594
rect 26910 22542 26962 22594
rect 27806 22542 27858 22594
rect 29598 22542 29650 22594
rect 29822 22542 29874 22594
rect 30494 22542 30546 22594
rect 31166 22542 31218 22594
rect 32622 22542 32674 22594
rect 39118 22542 39170 22594
rect 40238 22542 40290 22594
rect 47294 22542 47346 22594
rect 48750 22542 48802 22594
rect 51326 22542 51378 22594
rect 51886 22542 51938 22594
rect 53678 22542 53730 22594
rect 54350 22542 54402 22594
rect 55134 22542 55186 22594
rect 57262 22542 57314 22594
rect 22990 22430 23042 22482
rect 27470 22430 27522 22482
rect 28590 22430 28642 22482
rect 30158 22430 30210 22482
rect 31950 22430 32002 22482
rect 32286 22430 32338 22482
rect 33070 22430 33122 22482
rect 33518 22430 33570 22482
rect 35758 22430 35810 22482
rect 49422 22430 49474 22482
rect 50206 22430 50258 22482
rect 50654 22430 50706 22482
rect 53230 22430 53282 22482
rect 54686 22430 54738 22482
rect 56478 22430 56530 22482
rect 57150 22430 57202 22482
rect 29934 22318 29986 22370
rect 19838 22150 19890 22202
rect 19942 22150 19994 22202
rect 20046 22150 20098 22202
rect 50558 22150 50610 22202
rect 50662 22150 50714 22202
rect 50766 22150 50818 22202
rect 26126 21982 26178 22034
rect 23774 21870 23826 21922
rect 30606 21870 30658 21922
rect 39566 21870 39618 21922
rect 41022 21870 41074 21922
rect 41470 21870 41522 21922
rect 41918 21870 41970 21922
rect 47294 21870 47346 21922
rect 53006 21870 53058 21922
rect 21534 21758 21586 21810
rect 23214 21758 23266 21810
rect 25342 21758 25394 21810
rect 25678 21758 25730 21810
rect 27358 21758 27410 21810
rect 28702 21758 28754 21810
rect 29934 21758 29986 21810
rect 30942 21758 30994 21810
rect 31166 21758 31218 21810
rect 31726 21758 31778 21810
rect 34414 21758 34466 21810
rect 34974 21758 35026 21810
rect 35646 21758 35698 21810
rect 35870 21758 35922 21810
rect 38222 21758 38274 21810
rect 42366 21758 42418 21810
rect 43038 21758 43090 21810
rect 43598 21758 43650 21810
rect 45054 21758 45106 21810
rect 49422 21758 49474 21810
rect 52222 21758 52274 21810
rect 55246 21758 55298 21810
rect 56702 21758 56754 21810
rect 19854 21646 19906 21698
rect 20190 21646 20242 21698
rect 22654 21646 22706 21698
rect 25118 21646 25170 21698
rect 26462 21646 26514 21698
rect 29150 21646 29202 21698
rect 30270 21646 30322 21698
rect 31950 21646 32002 21698
rect 32286 21646 32338 21698
rect 44606 21646 44658 21698
rect 45166 21646 45218 21698
rect 45390 21646 45442 21698
rect 48862 21646 48914 21698
rect 49758 21646 49810 21698
rect 50094 21646 50146 21698
rect 50430 21646 50482 21698
rect 50990 21646 51042 21698
rect 51550 21646 51602 21698
rect 54126 21646 54178 21698
rect 24670 21534 24722 21586
rect 25454 21534 25506 21586
rect 26910 21534 26962 21586
rect 34078 21534 34130 21586
rect 36654 21534 36706 21586
rect 37102 21534 37154 21586
rect 37550 21534 37602 21586
rect 38670 21534 38722 21586
rect 39118 21534 39170 21586
rect 40014 21534 40066 21586
rect 44158 21534 44210 21586
rect 47854 21534 47906 21586
rect 53454 21534 53506 21586
rect 55470 21534 55522 21586
rect 56030 21534 56082 21586
rect 57150 21534 57202 21586
rect 36206 21422 36258 21474
rect 36654 21422 36706 21474
rect 36878 21422 36930 21474
rect 37550 21422 37602 21474
rect 38222 21422 38274 21474
rect 38670 21422 38722 21474
rect 42702 21422 42754 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 22542 20974 22594 21026
rect 22766 20974 22818 21026
rect 24222 20974 24274 21026
rect 35198 20974 35250 21026
rect 49198 20974 49250 21026
rect 51886 20974 51938 21026
rect 30270 20862 30322 20914
rect 32510 20862 32562 20914
rect 22878 20750 22930 20802
rect 23326 20750 23378 20802
rect 23774 20750 23826 20802
rect 24222 20750 24274 20802
rect 24670 20750 24722 20802
rect 26350 20750 26402 20802
rect 26798 20750 26850 20802
rect 27694 20750 27746 20802
rect 28142 20750 28194 20802
rect 33966 20750 34018 20802
rect 34974 20750 35026 20802
rect 36318 20750 36370 20802
rect 37214 20750 37266 20802
rect 44942 20750 44994 20802
rect 45502 20750 45554 20802
rect 49086 20750 49138 20802
rect 54910 20750 54962 20802
rect 55358 20750 55410 20802
rect 56254 20750 56306 20802
rect 18510 20638 18562 20690
rect 30606 20638 30658 20690
rect 30830 20638 30882 20690
rect 31166 20638 31218 20690
rect 31390 20638 31442 20690
rect 31614 20638 31666 20690
rect 31950 20638 32002 20690
rect 32846 20638 32898 20690
rect 33070 20638 33122 20690
rect 37550 20638 37602 20690
rect 40350 20638 40402 20690
rect 41470 20638 41522 20690
rect 41582 20638 41634 20690
rect 46398 20638 46450 20690
rect 48078 20638 48130 20690
rect 48638 20638 48690 20690
rect 49534 20638 49586 20690
rect 49758 20638 49810 20690
rect 50542 20638 50594 20690
rect 50878 20638 50930 20690
rect 53566 20638 53618 20690
rect 53790 20638 53842 20690
rect 55806 20638 55858 20690
rect 21422 20526 21474 20578
rect 21534 20526 21586 20578
rect 22094 20526 22146 20578
rect 31838 20526 31890 20578
rect 32062 20526 32114 20578
rect 35646 20526 35698 20578
rect 36206 20526 36258 20578
rect 41806 20526 41858 20578
rect 42702 20526 42754 20578
rect 45950 20526 46002 20578
rect 47630 20526 47682 20578
rect 19742 20414 19794 20466
rect 20302 20414 20354 20466
rect 20750 20414 20802 20466
rect 25454 20414 25506 20466
rect 25902 20414 25954 20466
rect 27134 20414 27186 20466
rect 27246 20414 27298 20466
rect 25454 20302 25506 20354
rect 25902 20302 25954 20354
rect 26910 20302 26962 20354
rect 28590 20414 28642 20466
rect 29486 20414 29538 20466
rect 29934 20414 29986 20466
rect 33518 20414 33570 20466
rect 38334 20414 38386 20466
rect 40798 20414 40850 20466
rect 43710 20414 43762 20466
rect 46846 20414 46898 20466
rect 54238 20414 54290 20466
rect 27358 20302 27410 20354
rect 27694 20302 27746 20354
rect 19838 20134 19890 20186
rect 19942 20134 19994 20186
rect 20046 20134 20098 20186
rect 50558 20134 50610 20186
rect 50662 20134 50714 20186
rect 50766 20134 50818 20186
rect 51438 19966 51490 20018
rect 20638 19854 20690 19906
rect 24110 19854 24162 19906
rect 25342 19854 25394 19906
rect 26014 19854 26066 19906
rect 28926 19854 28978 19906
rect 30718 19854 30770 19906
rect 33070 19854 33122 19906
rect 33742 19854 33794 19906
rect 34414 19854 34466 19906
rect 35198 19854 35250 19906
rect 46622 19854 46674 19906
rect 48302 19854 48354 19906
rect 52894 19854 52946 19906
rect 21086 19742 21138 19794
rect 22766 19742 22818 19794
rect 29598 19742 29650 19794
rect 30830 19742 30882 19794
rect 33406 19742 33458 19794
rect 34078 19742 34130 19794
rect 34750 19742 34802 19794
rect 38670 19742 38722 19794
rect 40910 19742 40962 19794
rect 41358 19742 41410 19794
rect 43486 19742 43538 19794
rect 49086 19742 49138 19794
rect 52222 19742 52274 19794
rect 54686 19742 54738 19794
rect 17726 19630 17778 19682
rect 20974 19630 21026 19682
rect 29262 19630 29314 19682
rect 29710 19630 29762 19682
rect 30606 19630 30658 19682
rect 31054 19630 31106 19682
rect 32286 19630 32338 19682
rect 35982 19630 36034 19682
rect 36318 19630 36370 19682
rect 39118 19630 39170 19682
rect 47742 19630 47794 19682
rect 49982 19630 50034 19682
rect 51550 19630 51602 19682
rect 51886 19630 51938 19682
rect 52558 19630 52610 19682
rect 53454 19630 53506 19682
rect 54014 19630 54066 19682
rect 24558 19518 24610 19570
rect 26462 19518 26514 19570
rect 26910 19518 26962 19570
rect 27582 19518 27634 19570
rect 28030 19518 28082 19570
rect 28478 19518 28530 19570
rect 45614 19518 45666 19570
rect 46062 19518 46114 19570
rect 47630 19518 47682 19570
rect 55470 19518 55522 19570
rect 19294 19406 19346 19458
rect 28254 19406 28306 19458
rect 28926 19406 28978 19458
rect 40238 19406 40290 19458
rect 44270 19406 44322 19458
rect 50094 19406 50146 19458
rect 22766 19294 22818 19346
rect 4478 19126 4530 19178
rect 4582 19126 4634 19178
rect 4686 19126 4738 19178
rect 35198 19126 35250 19178
rect 35302 19126 35354 19178
rect 35406 19126 35458 19178
rect 27694 18958 27746 19010
rect 28142 18958 28194 19010
rect 38894 18958 38946 19010
rect 40238 18958 40290 19010
rect 54686 18958 54738 19010
rect 26686 18846 26738 18898
rect 26910 18846 26962 18898
rect 27246 18846 27298 18898
rect 28254 18846 28306 18898
rect 33182 18846 33234 18898
rect 35982 18846 36034 18898
rect 36430 18846 36482 18898
rect 39230 18846 39282 18898
rect 40014 18846 40066 18898
rect 52782 18846 52834 18898
rect 53230 18846 53282 18898
rect 20414 18734 20466 18786
rect 21870 18734 21922 18786
rect 22318 18734 22370 18786
rect 27246 18734 27298 18786
rect 27694 18734 27746 18786
rect 28142 18734 28194 18786
rect 28590 18734 28642 18786
rect 35534 18734 35586 18786
rect 17502 18622 17554 18674
rect 18286 18622 18338 18674
rect 18958 18622 19010 18674
rect 19742 18622 19794 18674
rect 23214 18622 23266 18674
rect 31390 18678 31442 18730
rect 36430 18734 36482 18786
rect 40238 18734 40290 18786
rect 46398 18734 46450 18786
rect 49982 18734 50034 18786
rect 51886 18734 51938 18786
rect 52782 18734 52834 18786
rect 53230 18734 53282 18786
rect 53678 18734 53730 18786
rect 23886 18622 23938 18674
rect 31726 18622 31778 18674
rect 32846 18622 32898 18674
rect 35982 18622 36034 18674
rect 39342 18622 39394 18674
rect 40574 18622 40626 18674
rect 41246 18622 41298 18674
rect 41582 18622 41634 18674
rect 42702 18622 42754 18674
rect 48862 18622 48914 18674
rect 50094 18622 50146 18674
rect 57038 18622 57090 18674
rect 16606 18510 16658 18562
rect 17726 18510 17778 18562
rect 18062 18510 18114 18562
rect 21422 18510 21474 18562
rect 22878 18510 22930 18562
rect 23550 18510 23602 18562
rect 24446 18510 24498 18562
rect 25006 18510 25058 18562
rect 26350 18510 26402 18562
rect 29598 18510 29650 18562
rect 31278 18510 31330 18562
rect 33854 18510 33906 18562
rect 34750 18510 34802 18562
rect 38558 18510 38610 18562
rect 38894 18510 38946 18562
rect 39790 18510 39842 18562
rect 40910 18510 40962 18562
rect 42142 18510 42194 18562
rect 43374 18510 43426 18562
rect 47070 18510 47122 18562
rect 47966 18510 48018 18562
rect 17054 18398 17106 18450
rect 19182 18398 19234 18450
rect 19518 18398 19570 18450
rect 20078 18398 20130 18450
rect 25678 18398 25730 18450
rect 35086 18398 35138 18450
rect 45278 18398 45330 18450
rect 45726 18398 45778 18450
rect 47518 18398 47570 18450
rect 48414 18398 48466 18450
rect 18734 18286 18786 18338
rect 47518 18286 47570 18338
rect 48078 18286 48130 18338
rect 48750 18510 48802 18562
rect 49422 18510 49474 18562
rect 50654 18510 50706 18562
rect 50878 18510 50930 18562
rect 49086 18398 49138 18450
rect 19838 18118 19890 18170
rect 19942 18118 19994 18170
rect 20046 18118 20098 18170
rect 50558 18118 50610 18170
rect 50662 18118 50714 18170
rect 50766 18118 50818 18170
rect 54014 17950 54066 18002
rect 20750 17838 20802 17890
rect 22542 17838 22594 17890
rect 25790 17838 25842 17890
rect 26350 17838 26402 17890
rect 27358 17838 27410 17890
rect 29822 17838 29874 17890
rect 35310 17838 35362 17890
rect 38110 17838 38162 17890
rect 43486 17838 43538 17890
rect 48190 17838 48242 17890
rect 50542 17838 50594 17890
rect 53118 17838 53170 17890
rect 19742 17726 19794 17778
rect 28030 17726 28082 17778
rect 30494 17726 30546 17778
rect 30830 17726 30882 17778
rect 38446 17726 38498 17778
rect 41358 17726 41410 17778
rect 42926 17726 42978 17778
rect 46846 17726 46898 17778
rect 47406 17726 47458 17778
rect 47854 17726 47906 17778
rect 48078 17726 48130 17778
rect 49534 17726 49586 17778
rect 51102 17726 51154 17778
rect 52334 17726 52386 17778
rect 17614 17614 17666 17666
rect 18286 17614 18338 17666
rect 20078 17614 20130 17666
rect 20414 17614 20466 17666
rect 21310 17614 21362 17666
rect 21870 17614 21922 17666
rect 28702 17614 28754 17666
rect 29262 17614 29314 17666
rect 30158 17614 30210 17666
rect 43934 17614 43986 17666
rect 45950 17614 46002 17666
rect 47630 17614 47682 17666
rect 49870 17614 49922 17666
rect 50206 17614 50258 17666
rect 51662 17614 51714 17666
rect 53342 17614 53394 17666
rect 16830 17502 16882 17554
rect 18734 17502 18786 17554
rect 24222 17502 24274 17554
rect 24670 17502 24722 17554
rect 25342 17502 25394 17554
rect 26910 17502 26962 17554
rect 37662 17502 37714 17554
rect 42142 17502 42194 17554
rect 48862 17502 48914 17554
rect 44718 17390 44770 17442
rect 40462 17278 40514 17330
rect 4478 17110 4530 17162
rect 4582 17110 4634 17162
rect 4686 17110 4738 17162
rect 35198 17110 35250 17162
rect 35302 17110 35354 17162
rect 35406 17110 35458 17162
rect 37662 16830 37714 16882
rect 20750 16718 20802 16770
rect 27246 16718 27298 16770
rect 34974 16718 35026 16770
rect 38670 16718 38722 16770
rect 39006 16718 39058 16770
rect 50206 16718 50258 16770
rect 55582 16718 55634 16770
rect 15038 16606 15090 16658
rect 21422 16606 21474 16658
rect 21870 16606 21922 16658
rect 22206 16606 22258 16658
rect 23774 16606 23826 16658
rect 24446 16606 24498 16658
rect 25006 16606 25058 16658
rect 29822 16606 29874 16658
rect 30158 16606 30210 16658
rect 31278 16606 31330 16658
rect 37326 16606 37378 16658
rect 38222 16606 38274 16658
rect 40350 16606 40402 16658
rect 43038 16606 43090 16658
rect 46286 16606 46338 16658
rect 46734 16606 46786 16658
rect 48974 16606 49026 16658
rect 49758 16606 49810 16658
rect 50766 16606 50818 16658
rect 52558 16606 52610 16658
rect 23438 16494 23490 16546
rect 24110 16494 24162 16546
rect 25566 16494 25618 16546
rect 27582 16494 27634 16546
rect 28590 16494 28642 16546
rect 29150 16494 29202 16546
rect 29486 16494 29538 16546
rect 30606 16494 30658 16546
rect 31950 16494 32002 16546
rect 33854 16494 33906 16546
rect 37774 16494 37826 16546
rect 39230 16494 39282 16546
rect 39454 16494 39506 16546
rect 39902 16494 39954 16546
rect 43374 16494 43426 16546
rect 44830 16494 44882 16546
rect 47182 16494 47234 16546
rect 51214 16494 51266 16546
rect 52894 16494 52946 16546
rect 53566 16494 53618 16546
rect 54238 16494 54290 16546
rect 20190 16382 20242 16434
rect 21758 16382 21810 16434
rect 22990 16382 23042 16434
rect 26238 16382 26290 16434
rect 28254 16382 28306 16434
rect 33518 16382 33570 16434
rect 46062 16382 46114 16434
rect 52558 16382 52610 16434
rect 54574 16382 54626 16434
rect 54910 16382 54962 16434
rect 19182 16270 19234 16322
rect 44158 16270 44210 16322
rect 19838 16102 19890 16154
rect 19942 16102 19994 16154
rect 20046 16102 20098 16154
rect 50558 16102 50610 16154
rect 50662 16102 50714 16154
rect 50766 16102 50818 16154
rect 25566 15934 25618 15986
rect 40798 15934 40850 15986
rect 41134 15934 41186 15986
rect 51774 15934 51826 15986
rect 52782 15934 52834 15986
rect 19966 15822 20018 15874
rect 22654 15822 22706 15874
rect 24110 15822 24162 15874
rect 28478 15822 28530 15874
rect 37774 15822 37826 15874
rect 40350 15822 40402 15874
rect 41022 15822 41074 15874
rect 42366 15822 42418 15874
rect 44158 15822 44210 15874
rect 44942 15822 44994 15874
rect 47518 15822 47570 15874
rect 49310 15822 49362 15874
rect 50766 15822 50818 15874
rect 51214 15822 51266 15874
rect 19294 15710 19346 15762
rect 20526 15710 20578 15762
rect 21086 15710 21138 15762
rect 21758 15710 21810 15762
rect 25342 15710 25394 15762
rect 25454 15710 25506 15762
rect 25790 15710 25842 15762
rect 28814 15710 28866 15762
rect 30046 15710 30098 15762
rect 31950 15710 32002 15762
rect 33070 15710 33122 15762
rect 36206 15710 36258 15762
rect 36766 15710 36818 15762
rect 37438 15710 37490 15762
rect 39566 15710 39618 15762
rect 41358 15710 41410 15762
rect 42030 15710 42082 15762
rect 43486 15710 43538 15762
rect 46174 15710 46226 15762
rect 18958 15598 19010 15650
rect 19630 15598 19682 15650
rect 22990 15598 23042 15650
rect 23438 15598 23490 15650
rect 23886 15598 23938 15650
rect 24334 15598 24386 15650
rect 26014 15598 26066 15650
rect 28254 15598 28306 15650
rect 31278 15598 31330 15650
rect 37102 15598 37154 15650
rect 38334 15598 38386 15650
rect 38894 15598 38946 15650
rect 41694 15598 41746 15650
rect 42926 15598 42978 15650
rect 47070 15598 47122 15650
rect 47966 15598 48018 15650
rect 49758 15598 49810 15650
rect 52558 15598 52610 15650
rect 53342 15598 53394 15650
rect 54238 15598 54290 15650
rect 18174 15486 18226 15538
rect 18622 15486 18674 15538
rect 26798 15486 26850 15538
rect 29038 15486 29090 15538
rect 48862 15486 48914 15538
rect 50206 15486 50258 15538
rect 18174 15374 18226 15426
rect 18622 15374 18674 15426
rect 4478 15094 4530 15146
rect 4582 15094 4634 15146
rect 4686 15094 4738 15146
rect 35198 15094 35250 15146
rect 35302 15094 35354 15146
rect 35406 15094 35458 15146
rect 19070 14926 19122 14978
rect 30494 14926 30546 14978
rect 45390 14814 45442 14866
rect 46286 14814 46338 14866
rect 46958 14814 47010 14866
rect 20302 14702 20354 14754
rect 22654 14702 22706 14754
rect 29374 14702 29426 14754
rect 29710 14702 29762 14754
rect 32734 14702 32786 14754
rect 36430 14702 36482 14754
rect 38222 14702 38274 14754
rect 40238 14702 40290 14754
rect 41694 14702 41746 14754
rect 42366 14702 42418 14754
rect 43822 14702 43874 14754
rect 45838 14702 45890 14754
rect 46286 14702 46338 14754
rect 47182 14702 47234 14754
rect 47630 14702 47682 14754
rect 49310 14702 49362 14754
rect 50542 14702 50594 14754
rect 50990 14702 51042 14754
rect 51662 14702 51714 14754
rect 52110 14702 52162 14754
rect 52782 14702 52834 14754
rect 18622 14590 18674 14642
rect 22430 14590 22482 14642
rect 26014 14590 26066 14642
rect 26910 14590 26962 14642
rect 30158 14590 30210 14642
rect 30382 14590 30434 14642
rect 30606 14590 30658 14642
rect 30830 14590 30882 14642
rect 33182 14590 33234 14642
rect 34750 14590 34802 14642
rect 37102 14590 37154 14642
rect 37886 14590 37938 14642
rect 39678 14590 39730 14642
rect 45390 14590 45442 14642
rect 53230 14590 53282 14642
rect 22094 14478 22146 14530
rect 23998 14478 24050 14530
rect 24446 14478 24498 14530
rect 26238 14478 26290 14530
rect 34078 14478 34130 14530
rect 35646 14478 35698 14530
rect 39006 14478 39058 14530
rect 40574 14478 40626 14530
rect 44942 14478 44994 14530
rect 19854 14366 19906 14418
rect 20750 14366 20802 14418
rect 27694 14366 27746 14418
rect 28142 14366 28194 14418
rect 28590 14366 28642 14418
rect 32286 14366 32338 14418
rect 38558 14366 38610 14418
rect 44270 14366 44322 14418
rect 46734 14366 46786 14418
rect 50094 14366 50146 14418
rect 26574 14254 26626 14306
rect 27694 14254 27746 14306
rect 28254 14254 28306 14306
rect 33518 14254 33570 14306
rect 46734 14254 46786 14306
rect 47182 14254 47234 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 21982 13918 22034 13970
rect 26126 13918 26178 13970
rect 27694 13918 27746 13970
rect 37998 13918 38050 13970
rect 20974 13806 21026 13858
rect 21422 13806 21474 13858
rect 22766 13806 22818 13858
rect 23214 13806 23266 13858
rect 24222 13806 24274 13858
rect 24670 13806 24722 13858
rect 25454 13806 25506 13858
rect 25902 13806 25954 13858
rect 26350 13806 26402 13858
rect 26798 13806 26850 13858
rect 27694 13806 27746 13858
rect 29262 13806 29314 13858
rect 29710 13806 29762 13858
rect 32062 13806 32114 13858
rect 39006 13806 39058 13858
rect 40350 13806 40402 13858
rect 41358 13806 41410 13858
rect 42702 13806 42754 13858
rect 45614 13806 45666 13858
rect 51214 13806 51266 13858
rect 22318 13694 22370 13746
rect 41022 13694 41074 13746
rect 41694 13694 41746 13746
rect 42030 13694 42082 13746
rect 42366 13694 42418 13746
rect 43150 13694 43202 13746
rect 44494 13694 44546 13746
rect 47182 13694 47234 13746
rect 27246 13582 27298 13634
rect 28142 13582 28194 13634
rect 32510 13582 32562 13634
rect 33742 13582 33794 13634
rect 33966 13582 34018 13634
rect 34862 13582 34914 13634
rect 43822 13582 43874 13634
rect 46398 13582 46450 13634
rect 19406 13470 19458 13522
rect 20526 13470 20578 13522
rect 28814 13470 28866 13522
rect 30158 13470 30210 13522
rect 33182 13470 33234 13522
rect 34302 13470 34354 13522
rect 37326 13470 37378 13522
rect 38558 13470 38610 13522
rect 47854 13470 47906 13522
rect 4478 13078 4530 13130
rect 4582 13078 4634 13130
rect 4686 13078 4738 13130
rect 35198 13078 35250 13130
rect 35302 13078 35354 13130
rect 35406 13078 35458 13130
rect 26910 12910 26962 12962
rect 27358 12910 27410 12962
rect 27806 12910 27858 12962
rect 31950 12910 32002 12962
rect 33630 12910 33682 12962
rect 34302 12910 34354 12962
rect 44046 12910 44098 12962
rect 26574 12798 26626 12850
rect 37886 12798 37938 12850
rect 38558 12798 38610 12850
rect 39118 12798 39170 12850
rect 47742 12798 47794 12850
rect 21422 12686 21474 12738
rect 21870 12686 21922 12738
rect 23326 12686 23378 12738
rect 24222 12686 24274 12738
rect 27358 12686 27410 12738
rect 27806 12686 27858 12738
rect 33630 12686 33682 12738
rect 34078 12686 34130 12738
rect 34526 12686 34578 12738
rect 36430 12686 36482 12738
rect 38110 12686 38162 12738
rect 38558 12686 38610 12738
rect 17614 12574 17666 12626
rect 25790 12574 25842 12626
rect 32734 12574 32786 12626
rect 37102 12574 37154 12626
rect 39006 12574 39058 12626
rect 39342 12574 39394 12626
rect 39678 12574 39730 12626
rect 39902 12574 39954 12626
rect 40574 12574 40626 12626
rect 49982 12574 50034 12626
rect 18286 12462 18338 12514
rect 20638 12462 20690 12514
rect 24334 12462 24386 12514
rect 32398 12462 32450 12514
rect 32846 12462 32898 12514
rect 42926 12462 42978 12514
rect 44942 12462 44994 12514
rect 48190 12462 48242 12514
rect 23774 12350 23826 12402
rect 19838 12070 19890 12122
rect 19942 12070 19994 12122
rect 20046 12070 20098 12122
rect 50558 12070 50610 12122
rect 50662 12070 50714 12122
rect 50766 12070 50818 12122
rect 22094 11902 22146 11954
rect 22878 11902 22930 11954
rect 22878 11790 22930 11842
rect 43598 11790 43650 11842
rect 46286 11790 46338 11842
rect 17950 11678 18002 11730
rect 19854 11678 19906 11730
rect 22430 11678 22482 11730
rect 23102 11678 23154 11730
rect 23998 11678 24050 11730
rect 25342 11678 25394 11730
rect 27806 11678 27858 11730
rect 33406 11678 33458 11730
rect 34638 11678 34690 11730
rect 35870 11678 35922 11730
rect 44046 11678 44098 11730
rect 44494 11678 44546 11730
rect 46622 11678 46674 11730
rect 17502 11566 17554 11618
rect 23550 11566 23602 11618
rect 24222 11566 24274 11618
rect 30942 11566 30994 11618
rect 32286 11566 32338 11618
rect 33070 11566 33122 11618
rect 33742 11566 33794 11618
rect 34078 11566 34130 11618
rect 35198 11566 35250 11618
rect 48078 11566 48130 11618
rect 21086 11454 21138 11506
rect 21982 11454 22034 11506
rect 26350 11454 26402 11506
rect 27246 11454 27298 11506
rect 28254 11454 28306 11506
rect 28702 11454 28754 11506
rect 29150 11454 29202 11506
rect 30606 11454 30658 11506
rect 38782 11454 38834 11506
rect 39230 11454 39282 11506
rect 28142 11342 28194 11394
rect 28702 11230 28754 11282
rect 29262 11230 29314 11282
rect 4478 11062 4530 11114
rect 4582 11062 4634 11114
rect 4686 11062 4738 11114
rect 35198 11062 35250 11114
rect 35302 11062 35354 11114
rect 35406 11062 35458 11114
rect 27806 10894 27858 10946
rect 42590 10782 42642 10834
rect 20638 10670 20690 10722
rect 25902 10670 25954 10722
rect 28142 10670 28194 10722
rect 38782 10670 38834 10722
rect 16942 10558 16994 10610
rect 19070 10558 19122 10610
rect 21646 10558 21698 10610
rect 21982 10558 22034 10610
rect 22318 10558 22370 10610
rect 23438 10558 23490 10610
rect 25006 10558 25058 10610
rect 27134 10558 27186 10610
rect 30606 10558 30658 10610
rect 38334 10558 38386 10610
rect 39678 10558 39730 10610
rect 40126 10558 40178 10610
rect 16382 10446 16434 10498
rect 21310 10446 21362 10498
rect 22878 10446 22930 10498
rect 26910 10446 26962 10498
rect 27358 10446 27410 10498
rect 29374 10446 29426 10498
rect 29710 10446 29762 10498
rect 30046 10446 30098 10498
rect 33070 10446 33122 10498
rect 19742 10334 19794 10386
rect 24110 10334 24162 10386
rect 28590 10334 28642 10386
rect 34526 10334 34578 10386
rect 39230 10334 39282 10386
rect 42142 10334 42194 10386
rect 19838 10054 19890 10106
rect 19942 10054 19994 10106
rect 20046 10054 20098 10106
rect 50558 10054 50610 10106
rect 50662 10054 50714 10106
rect 50766 10054 50818 10106
rect 22430 9886 22482 9938
rect 23214 9886 23266 9938
rect 24670 9886 24722 9938
rect 23214 9774 23266 9826
rect 24222 9774 24274 9826
rect 24670 9774 24722 9826
rect 25342 9774 25394 9826
rect 26910 9774 26962 9826
rect 41918 9774 41970 9826
rect 20190 9662 20242 9714
rect 25902 9662 25954 9714
rect 26238 9662 26290 9714
rect 27470 9662 27522 9714
rect 28702 9662 28754 9714
rect 29598 9662 29650 9714
rect 42478 9662 42530 9714
rect 43038 9662 43090 9714
rect 43710 9662 43762 9714
rect 19630 9550 19682 9602
rect 19854 9550 19906 9602
rect 26574 9550 26626 9602
rect 28030 9550 28082 9602
rect 34750 9550 34802 9602
rect 36094 9550 36146 9602
rect 36542 9550 36594 9602
rect 38782 9550 38834 9602
rect 40238 9550 40290 9602
rect 40910 9550 40962 9602
rect 41246 9550 41298 9602
rect 41582 9550 41634 9602
rect 18510 9438 18562 9490
rect 18958 9438 19010 9490
rect 23662 9438 23714 9490
rect 32510 9438 32562 9490
rect 35198 9438 35250 9490
rect 35646 9438 35698 9490
rect 23662 9326 23714 9378
rect 24222 9326 24274 9378
rect 4478 9046 4530 9098
rect 4582 9046 4634 9098
rect 4686 9046 4738 9098
rect 35198 9046 35250 9098
rect 35302 9046 35354 9098
rect 35406 9046 35458 9098
rect 21310 8878 21362 8930
rect 35534 8878 35586 8930
rect 44046 8878 44098 8930
rect 28254 8766 28306 8818
rect 41134 8766 41186 8818
rect 19854 8654 19906 8706
rect 20302 8654 20354 8706
rect 22766 8654 22818 8706
rect 23326 8654 23378 8706
rect 30270 8654 30322 8706
rect 30718 8654 30770 8706
rect 36206 8654 36258 8706
rect 42030 8654 42082 8706
rect 19406 8542 19458 8594
rect 23662 8542 23714 8594
rect 23886 8542 23938 8594
rect 25006 8542 25058 8594
rect 29262 8542 29314 8594
rect 29822 8542 29874 8594
rect 31390 8542 31442 8594
rect 31614 8542 31666 8594
rect 32062 8542 32114 8594
rect 32734 8542 32786 8594
rect 37326 8542 37378 8594
rect 37662 8542 37714 8594
rect 40350 8542 40402 8594
rect 41806 8542 41858 8594
rect 43262 8542 43314 8594
rect 18958 8430 19010 8482
rect 20750 8430 20802 8482
rect 22206 8430 22258 8482
rect 24222 8430 24274 8482
rect 27246 8430 27298 8482
rect 31166 8430 31218 8482
rect 35086 8430 35138 8482
rect 40014 8430 40066 8482
rect 42254 8430 42306 8482
rect 19838 8038 19890 8090
rect 19942 8038 19994 8090
rect 20046 8038 20098 8090
rect 50558 8038 50610 8090
rect 50662 8038 50714 8090
rect 50766 8038 50818 8090
rect 30270 7870 30322 7922
rect 31278 7870 31330 7922
rect 37102 7870 37154 7922
rect 37662 7870 37714 7922
rect 24670 7758 24722 7810
rect 30270 7758 30322 7810
rect 30718 7758 30770 7810
rect 31166 7758 31218 7810
rect 34078 7758 34130 7810
rect 36654 7758 36706 7810
rect 37102 7758 37154 7810
rect 37550 7758 37602 7810
rect 40350 7758 40402 7810
rect 41022 7758 41074 7810
rect 41470 7758 41522 7810
rect 41918 7758 41970 7810
rect 25230 7646 25282 7698
rect 29262 7646 29314 7698
rect 33406 7646 33458 7698
rect 34526 7646 34578 7698
rect 35870 7646 35922 7698
rect 19406 7534 19458 7586
rect 19518 7534 19570 7586
rect 19966 7534 20018 7586
rect 20638 7534 20690 7586
rect 22990 7534 23042 7586
rect 25118 7534 25170 7586
rect 25902 7534 25954 7586
rect 26126 7534 26178 7586
rect 33070 7534 33122 7586
rect 33742 7534 33794 7586
rect 35198 7534 35250 7586
rect 31950 7422 32002 7474
rect 32398 7422 32450 7474
rect 23998 7310 24050 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 35758 6862 35810 6914
rect 32846 6750 32898 6802
rect 25678 6638 25730 6690
rect 21198 6526 21250 6578
rect 21534 6526 21586 6578
rect 21982 6526 22034 6578
rect 22654 6526 22706 6578
rect 29262 6526 29314 6578
rect 31838 6526 31890 6578
rect 33630 6526 33682 6578
rect 33854 6526 33906 6578
rect 28478 6414 28530 6466
rect 29934 6414 29986 6466
rect 34974 6414 35026 6466
rect 4174 6302 4226 6354
rect 4622 6302 4674 6354
rect 18174 6302 18226 6354
rect 20526 6302 20578 6354
rect 25342 6302 25394 6354
rect 33630 6302 33682 6354
rect 19838 6022 19890 6074
rect 19942 6022 19994 6074
rect 20046 6022 20098 6074
rect 50558 6022 50610 6074
rect 50662 6022 50714 6074
rect 50766 6022 50818 6074
rect 27022 5854 27074 5906
rect 27918 5854 27970 5906
rect 20078 5742 20130 5794
rect 20526 5742 20578 5794
rect 20974 5742 21026 5794
rect 22542 5742 22594 5794
rect 24334 5742 24386 5794
rect 25342 5742 25394 5794
rect 27022 5742 27074 5794
rect 27470 5742 27522 5794
rect 27918 5742 27970 5794
rect 28366 5742 28418 5794
rect 32398 5742 32450 5794
rect 21534 5630 21586 5682
rect 21870 5630 21922 5682
rect 22206 5630 22258 5682
rect 22990 5630 23042 5682
rect 23662 5630 23714 5682
rect 28814 5518 28866 5570
rect 29262 5518 29314 5570
rect 31838 5518 31890 5570
rect 33070 5518 33122 5570
rect 33630 5518 33682 5570
rect 25902 5406 25954 5458
rect 26350 5406 26402 5458
rect 31502 5406 31554 5458
rect 36094 5406 36146 5458
rect 25454 5294 25506 5346
rect 26126 5294 26178 5346
rect 26350 5294 26402 5346
rect 4478 5014 4530 5066
rect 4582 5014 4634 5066
rect 4686 5014 4738 5066
rect 35198 5014 35250 5066
rect 35302 5014 35354 5066
rect 35406 5014 35458 5066
rect 32398 4846 32450 4898
rect 32846 4846 32898 4898
rect 33518 4846 33570 4898
rect 23998 4622 24050 4674
rect 24670 4622 24722 4674
rect 25454 4622 25506 4674
rect 27694 4622 27746 4674
rect 28478 4622 28530 4674
rect 28926 4622 28978 4674
rect 32398 4622 32450 4674
rect 32846 4622 32898 4674
rect 33294 4622 33346 4674
rect 33742 4622 33794 4674
rect 19838 4006 19890 4058
rect 19942 4006 19994 4058
rect 20046 4006 20098 4058
rect 50558 4006 50610 4058
rect 50662 4006 50714 4058
rect 50766 4006 50818 4058
<< metal2 >>
rect 27552 59200 27664 60000
rect 27916 59276 28308 59332
rect 27580 59108 27636 59200
rect 27916 59108 27972 59276
rect 27580 59052 27972 59108
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 4476 55468 4740 55478
rect 4532 55412 4580 55468
rect 4636 55412 4684 55468
rect 4476 55402 4740 55412
rect 19836 54460 20100 54470
rect 19892 54404 19940 54460
rect 19996 54404 20044 54460
rect 19836 54394 20100 54404
rect 4476 53452 4740 53462
rect 4532 53396 4580 53452
rect 4636 53396 4684 53452
rect 4476 53386 4740 53396
rect 19836 52444 20100 52454
rect 19892 52388 19940 52444
rect 19996 52388 20044 52444
rect 19836 52378 20100 52388
rect 5852 52164 5908 52174
rect 5852 52070 5908 52108
rect 4476 51436 4740 51446
rect 4532 51380 4580 51436
rect 4636 51380 4684 51436
rect 4476 51370 4740 51380
rect 19836 50428 20100 50438
rect 19892 50372 19940 50428
rect 19996 50372 20044 50428
rect 19836 50362 20100 50372
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 19836 48412 20100 48422
rect 19892 48356 19940 48412
rect 19996 48356 20044 48412
rect 19836 48346 20100 48356
rect 6188 48130 6244 48142
rect 6188 48078 6190 48130
rect 6242 48078 6244 48130
rect 3388 47906 3444 47918
rect 3388 47854 3390 47906
rect 3442 47854 3444 47906
rect 3052 47794 3108 47806
rect 3052 47742 3054 47794
rect 3106 47742 3108 47794
rect 1820 45780 1876 45790
rect 1708 45778 1876 45780
rect 1708 45726 1822 45778
rect 1874 45726 1876 45778
rect 1708 45724 1876 45726
rect 1708 45332 1764 45724
rect 1820 45714 1876 45724
rect 1708 44436 1764 45276
rect 3052 45332 3108 47742
rect 3052 45266 3108 45276
rect 1820 44884 1876 44894
rect 1820 44882 1988 44884
rect 1820 44830 1822 44882
rect 1874 44830 1988 44882
rect 1820 44828 1988 44830
rect 1820 44818 1876 44828
rect 1820 44436 1876 44446
rect 1708 44380 1820 44436
rect 1820 44098 1876 44380
rect 1820 44046 1822 44098
rect 1874 44046 1876 44098
rect 1820 44034 1876 44046
rect 1932 43204 1988 44828
rect 2380 44882 2436 44894
rect 2380 44830 2382 44882
rect 2434 44830 2436 44882
rect 2380 44660 2436 44830
rect 2380 44594 2436 44604
rect 3388 44660 3444 47854
rect 3948 47906 4004 47918
rect 3948 47854 3950 47906
rect 4002 47854 4004 47906
rect 3948 47012 4004 47854
rect 4476 47404 4740 47414
rect 4532 47348 4580 47404
rect 4636 47348 4684 47404
rect 4476 47338 4740 47348
rect 3948 46946 4004 46956
rect 4508 47012 4564 47022
rect 4508 45890 4564 46956
rect 5628 47012 5684 47022
rect 5628 46918 5684 46956
rect 5740 47010 5796 47022
rect 5740 46958 5742 47010
rect 5794 46958 5796 47010
rect 5740 46898 5796 46958
rect 5740 46846 5742 46898
rect 5794 46846 5796 46898
rect 5740 46834 5796 46846
rect 6188 46674 6244 48078
rect 26012 47906 26068 47918
rect 26012 47854 26014 47906
rect 26066 47854 26068 47906
rect 24668 47796 24724 47806
rect 24668 47702 24724 47740
rect 25564 47796 25620 47806
rect 26012 47796 26068 47854
rect 25564 47794 26068 47796
rect 25564 47742 25566 47794
rect 25618 47742 26068 47794
rect 25564 47740 26068 47742
rect 25564 47730 25620 47740
rect 6524 47684 6580 47694
rect 6300 47682 6580 47684
rect 6300 47630 6526 47682
rect 6578 47630 6580 47682
rect 6300 47628 6580 47630
rect 6300 47122 6356 47628
rect 6524 47618 6580 47628
rect 6300 47070 6302 47122
rect 6354 47070 6356 47122
rect 6300 47058 6356 47070
rect 22540 46900 22596 46910
rect 22540 46898 22820 46900
rect 22540 46846 22542 46898
rect 22594 46846 22820 46898
rect 22540 46844 22820 46846
rect 22540 46834 22596 46844
rect 6188 46622 6190 46674
rect 6242 46622 6244 46674
rect 4508 45838 4510 45890
rect 4562 45838 4564 45890
rect 4508 45826 4564 45838
rect 5068 45892 5124 45902
rect 5068 45890 5684 45892
rect 5068 45838 5070 45890
rect 5122 45838 5684 45890
rect 5068 45836 5684 45838
rect 5068 45826 5124 45836
rect 4172 45780 4228 45790
rect 4172 45332 4228 45724
rect 4476 45388 4740 45398
rect 4532 45332 4580 45388
rect 4636 45332 4684 45388
rect 4228 45276 4340 45332
rect 4476 45322 4740 45332
rect 4172 45266 4228 45276
rect 4284 45108 4340 45276
rect 5628 45218 5684 45836
rect 6188 45780 6244 46622
rect 21644 46674 21700 46686
rect 21644 46622 21646 46674
rect 21698 46622 21700 46674
rect 19836 46396 20100 46406
rect 19892 46340 19940 46396
rect 19996 46340 20044 46396
rect 19836 46330 20100 46340
rect 6188 45714 6244 45724
rect 7196 46114 7252 46126
rect 7196 46062 7198 46114
rect 7250 46062 7252 46114
rect 7196 45780 7252 46062
rect 8428 45892 8484 45902
rect 8428 45890 8932 45892
rect 8428 45838 8430 45890
rect 8482 45838 8932 45890
rect 8428 45836 8932 45838
rect 8428 45826 8484 45836
rect 7196 45714 7252 45724
rect 5628 45166 5630 45218
rect 5682 45166 5684 45218
rect 4284 45052 4564 45108
rect 3388 44594 3444 44604
rect 4508 44660 4564 45052
rect 4508 44658 4900 44660
rect 4508 44606 4510 44658
rect 4562 44606 4900 44658
rect 4508 44604 4900 44606
rect 4508 44594 4564 44604
rect 4844 44098 4900 44604
rect 4844 44046 4846 44098
rect 4898 44046 4900 44098
rect 2156 43874 2212 43886
rect 2156 43822 2158 43874
rect 2210 43822 2212 43874
rect 2156 43708 2212 43822
rect 2716 43874 2772 43886
rect 2716 43822 2718 43874
rect 2770 43822 2772 43874
rect 2156 43652 2436 43708
rect 1932 43138 1988 43148
rect 1820 42868 1876 42878
rect 1708 42866 1876 42868
rect 1708 42814 1822 42866
rect 1874 42814 1876 42866
rect 1708 42812 1876 42814
rect 1708 40964 1764 42812
rect 1820 42802 1876 42812
rect 2380 42866 2436 43652
rect 2716 43204 2772 43822
rect 4476 43372 4740 43382
rect 4532 43316 4580 43372
rect 4636 43316 4684 43372
rect 4476 43306 4740 43316
rect 2716 43138 2772 43148
rect 2380 42814 2382 42866
rect 2434 42814 2436 42866
rect 2380 41972 2436 42814
rect 4620 42644 4676 42654
rect 4844 42644 4900 44046
rect 4956 44658 5012 44670
rect 4956 44606 4958 44658
rect 5010 44606 5012 44658
rect 4956 42868 5012 44606
rect 5628 43876 5684 45166
rect 5740 45668 5796 45678
rect 5740 44882 5796 45612
rect 7644 45668 7700 45678
rect 7644 45574 7700 45612
rect 8764 45668 8820 45678
rect 5740 44830 5742 44882
rect 5794 44830 5796 44882
rect 5740 44818 5796 44830
rect 6076 45556 6132 45566
rect 6076 44884 6132 45500
rect 8316 45556 8372 45566
rect 8316 45462 8372 45500
rect 6636 44884 6692 44894
rect 6076 44882 6356 44884
rect 6076 44830 6078 44882
rect 6130 44830 6356 44882
rect 6076 44828 6356 44830
rect 6076 44818 6132 44828
rect 6076 44660 6132 44670
rect 5740 43876 5796 43886
rect 5628 43874 5796 43876
rect 5628 43822 5742 43874
rect 5794 43822 5796 43874
rect 5628 43820 5796 43822
rect 5740 43810 5796 43820
rect 5292 43650 5348 43662
rect 5292 43598 5294 43650
rect 5346 43598 5348 43650
rect 5292 42868 5348 43598
rect 5628 43204 5684 43214
rect 5628 43110 5684 43148
rect 6076 43202 6132 44604
rect 6300 43874 6356 44828
rect 6636 44790 6692 44828
rect 8764 44660 8820 45612
rect 8540 44658 8820 44660
rect 8540 44606 8766 44658
rect 8818 44606 8820 44658
rect 8540 44604 8820 44606
rect 8540 44100 8596 44604
rect 8764 44594 8820 44604
rect 8540 44006 8596 44044
rect 8876 44098 8932 45836
rect 11676 45890 11732 45902
rect 11676 45838 11678 45890
rect 11730 45838 11732 45890
rect 9660 45780 9716 45790
rect 9660 45686 9716 45724
rect 11564 45554 11620 45566
rect 11564 45502 11566 45554
rect 11618 45502 11620 45554
rect 9548 44996 9604 45006
rect 9212 44660 9268 44670
rect 9212 44566 9268 44604
rect 8876 44046 8878 44098
rect 8930 44046 8932 44098
rect 8876 44034 8932 44046
rect 6300 43822 6302 43874
rect 6354 43822 6356 43874
rect 6300 43810 6356 43822
rect 9548 43708 9604 44940
rect 10220 44996 10276 45006
rect 9660 44884 9716 44894
rect 9716 44828 10164 44884
rect 9660 44790 9716 44828
rect 10108 44212 10164 44828
rect 10220 44882 10276 44940
rect 11564 44996 11620 45502
rect 11676 45108 11732 45838
rect 11676 45042 11732 45052
rect 12796 45108 12852 45118
rect 12796 45014 12852 45052
rect 11564 44930 11620 44940
rect 10220 44830 10222 44882
rect 10274 44830 10276 44882
rect 10220 44818 10276 44830
rect 10332 44660 10388 44670
rect 10220 44212 10276 44222
rect 10108 44210 10276 44212
rect 10108 44158 10222 44210
rect 10274 44158 10276 44210
rect 10108 44156 10276 44158
rect 10220 44146 10276 44156
rect 9884 44100 9940 44110
rect 9548 43652 9716 43708
rect 6076 43150 6078 43202
rect 6130 43150 6132 43202
rect 6076 43138 6132 43150
rect 5740 42868 5796 42878
rect 5292 42866 5796 42868
rect 5292 42814 5742 42866
rect 5794 42814 5796 42866
rect 5292 42812 5796 42814
rect 4956 42802 5012 42812
rect 5740 42802 5796 42812
rect 6188 42868 6244 42878
rect 6188 42774 6244 42812
rect 9660 42866 9716 43652
rect 9660 42814 9662 42866
rect 9714 42814 9716 42866
rect 9660 42802 9716 42814
rect 4620 42642 4900 42644
rect 4620 42590 4622 42642
rect 4674 42590 4900 42642
rect 4620 42588 4900 42590
rect 4956 42642 5012 42654
rect 4956 42590 4958 42642
rect 5010 42590 5012 42642
rect 4620 42578 4676 42588
rect 4956 42308 5012 42590
rect 3500 42252 5012 42308
rect 6636 42642 6692 42654
rect 6636 42590 6638 42642
rect 6690 42590 6692 42642
rect 3500 42082 3556 42252
rect 3500 42030 3502 42082
rect 3554 42030 3556 42082
rect 3500 42018 3556 42030
rect 6636 42082 6692 42590
rect 6636 42030 6638 42082
rect 6690 42030 6692 42082
rect 2380 41906 2436 41916
rect 3388 41972 3444 41982
rect 3388 41878 3444 41916
rect 3836 41858 3892 41870
rect 3836 41806 3838 41858
rect 3890 41806 3892 41858
rect 1820 41748 1876 41758
rect 1820 41746 1988 41748
rect 1820 41694 1822 41746
rect 1874 41694 1988 41746
rect 1820 41692 1988 41694
rect 1820 41682 1876 41692
rect 1708 40898 1764 40908
rect 1820 41524 1876 41534
rect 1820 40850 1876 41468
rect 1820 40798 1822 40850
rect 1874 40798 1876 40850
rect 1820 40786 1876 40798
rect 1820 40404 1876 40414
rect 1932 40404 1988 41692
rect 3052 41746 3108 41758
rect 3052 41694 3054 41746
rect 3106 41694 3108 41746
rect 2380 40964 2436 40974
rect 2380 40850 2436 40908
rect 2380 40798 2382 40850
rect 2434 40798 2436 40850
rect 2380 40786 2436 40798
rect 1876 40348 1988 40404
rect 3052 40404 3108 41694
rect 1820 40066 1876 40348
rect 3052 40338 3108 40348
rect 1820 40014 1822 40066
rect 1874 40014 1876 40066
rect 1820 40002 1876 40014
rect 3836 39956 3892 41806
rect 4396 41858 4452 41870
rect 4396 41806 4398 41858
rect 4450 41806 4452 41858
rect 4396 41524 4452 41806
rect 5740 41636 5796 41646
rect 4396 41458 4452 41468
rect 5628 41524 5684 41534
rect 4476 41356 4740 41366
rect 4532 41300 4580 41356
rect 4636 41300 4684 41356
rect 4476 41290 4740 41300
rect 5628 41186 5684 41468
rect 5628 41134 5630 41186
rect 5682 41134 5684 41186
rect 5628 41122 5684 41134
rect 5740 40850 5796 41580
rect 6076 40964 6132 40974
rect 6076 40870 6132 40908
rect 5740 40798 5742 40850
rect 5794 40798 5796 40850
rect 5740 40786 5796 40798
rect 4508 40626 4564 40638
rect 4508 40574 4510 40626
rect 4562 40574 4564 40626
rect 3836 39890 3892 39900
rect 4060 40404 4116 40414
rect 4060 40068 4116 40348
rect 4508 40068 4564 40574
rect 4956 40628 5012 40638
rect 4956 40534 5012 40572
rect 6188 40628 6244 40638
rect 6188 40534 6244 40572
rect 6636 40292 6692 42030
rect 9324 42644 9380 42654
rect 9884 42644 9940 44044
rect 10332 44098 10388 44604
rect 10332 44046 10334 44098
rect 10386 44046 10388 44098
rect 10332 44034 10388 44046
rect 12348 44658 12404 44670
rect 12348 44606 12350 44658
rect 12402 44606 12404 44658
rect 12348 44100 12404 44606
rect 19836 44380 20100 44390
rect 19892 44324 19940 44380
rect 19996 44324 20044 44380
rect 19836 44314 20100 44324
rect 13580 44100 13636 44110
rect 10892 43988 10948 43998
rect 10892 43874 10948 43932
rect 10892 43822 10894 43874
rect 10946 43822 10948 43874
rect 10892 43708 10948 43822
rect 10220 43652 10948 43708
rect 11452 43874 11508 43886
rect 11452 43822 11454 43874
rect 11506 43822 11508 43874
rect 10220 42866 10276 43652
rect 10220 42814 10222 42866
rect 10274 42814 10276 42866
rect 10220 42802 10276 42814
rect 10780 43204 10836 43214
rect 9324 42642 9940 42644
rect 9324 42590 9326 42642
rect 9378 42590 9940 42642
rect 9324 42588 9940 42590
rect 6972 41636 7028 41646
rect 6972 41542 7028 41580
rect 9324 40628 9380 42588
rect 10780 41858 10836 43148
rect 11452 43204 11508 43822
rect 11452 43138 11508 43148
rect 12348 43652 12404 44044
rect 13468 44098 13636 44100
rect 13468 44046 13582 44098
rect 13634 44046 13636 44098
rect 13468 44044 13636 44046
rect 12348 42642 12404 43596
rect 12796 43876 12852 43886
rect 12796 43090 12852 43820
rect 13468 43652 13524 44044
rect 13580 44034 13636 44044
rect 14476 43988 14532 43998
rect 14476 43894 14532 43932
rect 18172 43986 18228 43998
rect 18172 43934 18174 43986
rect 18226 43934 18228 43986
rect 14588 43876 14644 43886
rect 14588 43782 14644 43820
rect 17388 43874 17444 43886
rect 17388 43822 17390 43874
rect 17442 43822 17444 43874
rect 16828 43762 16884 43774
rect 16828 43710 16830 43762
rect 16882 43710 16884 43762
rect 16828 43708 16884 43710
rect 17388 43708 17444 43822
rect 18172 43708 18228 43934
rect 12796 43038 12798 43090
rect 12850 43038 12852 43090
rect 12796 43026 12852 43038
rect 13356 43596 13468 43652
rect 12348 42590 12350 42642
rect 12402 42590 12404 42642
rect 10780 41806 10782 41858
rect 10834 41806 10836 41858
rect 10780 41794 10836 41806
rect 11340 41858 11396 41870
rect 11340 41806 11342 41858
rect 11394 41806 11396 41858
rect 10444 41746 10500 41758
rect 10444 41694 10446 41746
rect 10498 41694 10500 41746
rect 9660 41636 9716 41646
rect 9660 40850 9716 41580
rect 9660 40798 9662 40850
rect 9714 40798 9716 40850
rect 9660 40786 9716 40798
rect 10220 40850 10276 40862
rect 10220 40798 10222 40850
rect 10274 40798 10276 40850
rect 10220 40740 10276 40798
rect 10220 40674 10276 40684
rect 9324 40534 9380 40572
rect 10444 40628 10500 41694
rect 11340 41636 11396 41806
rect 11340 41570 11396 41580
rect 6860 40292 6916 40302
rect 6636 40236 6860 40292
rect 4060 40012 4564 40068
rect 6860 40066 6916 40236
rect 6860 40014 6862 40066
rect 6914 40014 6916 40066
rect 3836 39732 3892 39742
rect 4060 39732 4116 40012
rect 4956 39956 5012 39966
rect 3836 39730 4116 39732
rect 3836 39678 3838 39730
rect 3890 39678 4116 39730
rect 3836 39676 4116 39678
rect 4172 39842 4228 39854
rect 4172 39790 4174 39842
rect 4226 39790 4228 39842
rect 3836 38724 3892 39676
rect 3836 38658 3892 38668
rect 3500 37826 3556 37838
rect 3500 37774 3502 37826
rect 3554 37774 3556 37826
rect 3164 37714 3220 37726
rect 3164 37662 3166 37714
rect 3218 37662 3220 37714
rect 2716 36036 2772 36046
rect 2716 35942 2772 35980
rect 3164 36036 3220 37662
rect 3164 35970 3220 35980
rect 3500 36148 3556 37774
rect 4060 37828 4116 37838
rect 4172 37828 4228 39790
rect 4732 39844 4788 39854
rect 4732 39842 4900 39844
rect 4732 39790 4734 39842
rect 4786 39790 4900 39842
rect 4732 39788 4900 39790
rect 4732 39778 4788 39788
rect 4060 37826 4228 37828
rect 4060 37774 4062 37826
rect 4114 37774 4228 37826
rect 4060 37772 4228 37774
rect 4060 37762 4116 37772
rect 4172 37156 4228 37772
rect 4284 39732 4340 39742
rect 4284 37828 4340 39676
rect 4476 39340 4740 39350
rect 4532 39284 4580 39340
rect 4636 39284 4684 39340
rect 4476 39274 4740 39284
rect 4620 38724 4676 38734
rect 4620 38630 4676 38668
rect 4844 38276 4900 39788
rect 4956 39172 5012 39900
rect 4956 39078 5012 39116
rect 5068 38724 5124 38734
rect 5740 38724 5796 38734
rect 5068 38722 5796 38724
rect 5068 38670 5070 38722
rect 5122 38670 5742 38722
rect 5794 38670 5796 38722
rect 5068 38668 5796 38670
rect 5068 38658 5124 38668
rect 5740 38658 5796 38668
rect 6076 38724 6132 38734
rect 6076 38610 6132 38668
rect 6860 38724 6916 40014
rect 10444 39730 10500 40572
rect 10780 40740 10836 40750
rect 10780 39842 10836 40684
rect 12348 40626 12404 42590
rect 13356 42644 13412 43596
rect 13468 43586 13524 43596
rect 14028 43650 14084 43662
rect 14028 43598 14030 43650
rect 14082 43598 14084 43650
rect 13468 43204 13524 43214
rect 13468 43110 13524 43148
rect 13580 42868 13636 42878
rect 14028 42868 14084 43598
rect 13580 42866 14084 42868
rect 13580 42814 13582 42866
rect 13634 42814 14084 42866
rect 13580 42812 14084 42814
rect 16716 43652 17444 43708
rect 18060 43652 18228 43708
rect 20188 43764 20244 43802
rect 20188 43698 20244 43708
rect 21644 43764 21700 46622
rect 22092 46674 22148 46686
rect 22092 46622 22094 46674
rect 22146 46622 22148 46674
rect 22092 45218 22148 46622
rect 22092 45166 22094 45218
rect 22146 45166 22148 45218
rect 22092 45154 22148 45166
rect 21644 43698 21700 43708
rect 22204 44996 22260 45006
rect 22204 43876 22260 44940
rect 22764 44884 22820 46844
rect 22764 44818 22820 44828
rect 22988 46898 23044 46910
rect 22988 46846 22990 46898
rect 23042 46846 23044 46898
rect 22988 45218 23044 46846
rect 25004 46898 25060 46910
rect 25004 46846 25006 46898
rect 25058 46846 25060 46898
rect 25004 45780 25060 46846
rect 25004 45714 25060 45724
rect 25788 46674 25844 46686
rect 25788 46622 25790 46674
rect 25842 46622 25844 46674
rect 22988 45166 22990 45218
rect 23042 45166 23044 45218
rect 16716 42868 16772 43652
rect 17052 42868 17108 42878
rect 16716 42866 17108 42868
rect 16716 42814 17054 42866
rect 17106 42814 17108 42866
rect 16716 42812 17108 42814
rect 13580 42802 13636 42812
rect 13356 42084 13412 42588
rect 16716 42644 16772 42812
rect 16716 42550 16772 42588
rect 13468 42084 13524 42094
rect 13356 42082 13524 42084
rect 13356 42030 13470 42082
rect 13522 42030 13524 42082
rect 13356 42028 13524 42030
rect 12348 40574 12350 40626
rect 12402 40574 12404 40626
rect 12348 40562 12404 40574
rect 12796 40628 12852 40638
rect 12796 40534 12852 40572
rect 13356 40516 13412 42028
rect 13468 42018 13524 42028
rect 13916 41860 13972 41870
rect 14476 41860 14532 41870
rect 13916 41858 14532 41860
rect 13916 41806 13918 41858
rect 13970 41806 14478 41858
rect 14530 41806 14532 41858
rect 13916 41804 14532 41806
rect 13916 41794 13972 41804
rect 14476 41794 14532 41804
rect 14364 41636 14420 41646
rect 14364 41542 14420 41580
rect 17052 41186 17108 42812
rect 17836 42644 17892 42654
rect 17052 41134 17054 41186
rect 17106 41134 17108 41186
rect 17052 40964 17108 41134
rect 17388 42642 17892 42644
rect 17388 42590 17838 42642
rect 17890 42590 17892 42642
rect 17388 42588 17892 42590
rect 17164 40964 17220 40974
rect 17052 40962 17220 40964
rect 17052 40910 17166 40962
rect 17218 40910 17220 40962
rect 17052 40908 17220 40910
rect 17164 40898 17220 40908
rect 13468 40740 13524 40750
rect 13468 40646 13524 40684
rect 13580 40628 13636 40638
rect 13580 40534 13636 40572
rect 13356 40460 13524 40516
rect 13468 40068 13524 40460
rect 17388 40178 17444 42588
rect 17836 42578 17892 42588
rect 17836 42420 17892 42430
rect 17612 41186 17668 41198
rect 17612 41134 17614 41186
rect 17666 41134 17668 41186
rect 17612 40962 17668 41134
rect 17612 40910 17614 40962
rect 17666 40910 17668 40962
rect 17612 40852 17668 40910
rect 17612 40786 17668 40796
rect 17388 40126 17390 40178
rect 17442 40126 17444 40178
rect 17388 40114 17444 40126
rect 13468 40066 14420 40068
rect 13468 40014 13470 40066
rect 13522 40014 14420 40066
rect 13468 40012 14420 40014
rect 13468 40002 13524 40012
rect 10780 39790 10782 39842
rect 10834 39790 10836 39842
rect 10780 39778 10836 39790
rect 11340 39844 11396 39854
rect 11340 39750 11396 39788
rect 11676 39844 11732 39854
rect 10444 39678 10446 39730
rect 10498 39678 10500 39730
rect 6860 38658 6916 38668
rect 7308 39618 7364 39630
rect 7308 39566 7310 39618
rect 7362 39566 7364 39618
rect 6076 38558 6078 38610
rect 6130 38558 6132 38610
rect 4844 38210 4900 38220
rect 5516 38276 5572 38286
rect 5572 38220 5684 38276
rect 5516 38210 5572 38220
rect 4284 37762 4340 37772
rect 4476 37324 4740 37334
rect 4532 37268 4580 37324
rect 4636 37268 4684 37324
rect 4476 37258 4740 37268
rect 4396 37156 4452 37166
rect 4172 37154 4452 37156
rect 4172 37102 4398 37154
rect 4450 37102 4452 37154
rect 4172 37100 4452 37102
rect 4396 37090 4452 37100
rect 4508 37156 4564 37166
rect 4508 36818 4564 37100
rect 4508 36766 4510 36818
rect 4562 36766 4564 36818
rect 4508 36754 4564 36766
rect 5628 36818 5684 38220
rect 5628 36766 5630 36818
rect 5682 36766 5684 36818
rect 5628 36754 5684 36766
rect 6076 38052 6132 38558
rect 7084 38276 7140 38286
rect 6300 38164 6356 38174
rect 6188 38052 6244 38062
rect 6076 38050 6244 38052
rect 6076 37998 6190 38050
rect 6242 37998 6244 38050
rect 6076 37996 6244 37998
rect 4060 36594 4116 36606
rect 4060 36542 4062 36594
rect 4114 36542 4116 36594
rect 3724 36148 3780 36158
rect 3500 36146 3780 36148
rect 3500 36094 3726 36146
rect 3778 36094 3780 36146
rect 3500 36092 3780 36094
rect 3052 35810 3108 35822
rect 3052 35758 3054 35810
rect 3106 35758 3108 35810
rect 2380 34916 2436 34926
rect 1820 34802 1876 34814
rect 1820 34750 1822 34802
rect 1874 34750 1876 34802
rect 1820 34130 1876 34750
rect 2380 34802 2436 34860
rect 3052 34916 3108 35758
rect 3500 35812 3556 36092
rect 3724 36082 3780 36092
rect 4060 36036 4116 36542
rect 4956 36596 5012 36606
rect 4956 36502 5012 36540
rect 4844 36482 4900 36494
rect 4844 36430 4846 36482
rect 4898 36430 4900 36482
rect 3612 35812 3668 35822
rect 3500 35810 3668 35812
rect 3500 35758 3614 35810
rect 3666 35758 3668 35810
rect 3500 35756 3668 35758
rect 3612 35746 3668 35756
rect 3052 34850 3108 34860
rect 2380 34750 2382 34802
rect 2434 34750 2436 34802
rect 2380 34738 2436 34750
rect 4060 34692 4116 35980
rect 4172 36372 4228 36382
rect 4172 35028 4228 36316
rect 4508 36148 4564 36158
rect 4844 36148 4900 36430
rect 4508 36146 4900 36148
rect 4508 36094 4510 36146
rect 4562 36094 4900 36146
rect 4508 36092 4900 36094
rect 4508 36082 4564 36092
rect 5852 36036 5908 36046
rect 6076 36036 6132 37996
rect 6188 37986 6244 37996
rect 6188 36820 6244 36830
rect 6300 36820 6356 38108
rect 7084 38162 7140 38220
rect 7084 38110 7086 38162
rect 7138 38110 7140 38162
rect 7084 38098 7140 38110
rect 7196 38052 7252 38062
rect 7308 38052 7364 39566
rect 8316 39172 8372 39182
rect 8316 38834 8372 39116
rect 8316 38782 8318 38834
rect 8370 38782 8372 38834
rect 8316 38770 8372 38782
rect 8876 38834 8932 38846
rect 8876 38782 8878 38834
rect 8930 38782 8932 38834
rect 7532 38164 7588 38174
rect 7532 38070 7588 38108
rect 8876 38164 8932 38782
rect 8876 38098 8932 38108
rect 7196 38050 7364 38052
rect 7196 37998 7198 38050
rect 7250 37998 7364 38050
rect 7196 37996 7364 37998
rect 7196 37986 7252 37996
rect 7644 37826 7700 37838
rect 7644 37774 7646 37826
rect 7698 37774 7700 37826
rect 6636 37602 6692 37614
rect 6636 37550 6638 37602
rect 6690 37550 6692 37602
rect 6636 37156 6692 37550
rect 6636 37090 6692 37100
rect 7644 36932 7700 37774
rect 10444 37716 10500 39678
rect 11676 37826 11732 39788
rect 12684 39844 12740 39854
rect 12684 39170 12740 39788
rect 12684 39118 12686 39170
rect 12738 39118 12740 39170
rect 12684 39106 12740 39118
rect 12796 39620 12852 39630
rect 12796 38834 12852 39564
rect 13916 39620 13972 39630
rect 13916 39526 13972 39564
rect 12796 38782 12798 38834
rect 12850 38782 12852 38834
rect 12796 38770 12852 38782
rect 11676 37774 11678 37826
rect 11730 37774 11732 37826
rect 11676 37762 11732 37774
rect 12236 38724 12292 38734
rect 12236 37826 12292 38668
rect 13468 38724 13524 38734
rect 13468 38630 13524 38668
rect 12236 37774 12238 37826
rect 12290 37774 12292 37826
rect 12236 37762 12292 37774
rect 13580 38610 13636 38622
rect 13580 38558 13582 38610
rect 13634 38558 13636 38610
rect 11340 37716 11396 37726
rect 10444 37714 11396 37716
rect 10444 37662 11342 37714
rect 11394 37662 11396 37714
rect 10444 37660 11396 37662
rect 7644 36866 7700 36876
rect 8764 36932 8820 36942
rect 8764 36838 8820 36876
rect 6188 36818 6356 36820
rect 6188 36766 6190 36818
rect 6242 36766 6356 36818
rect 6188 36764 6356 36766
rect 6188 36754 6244 36764
rect 5852 36034 6132 36036
rect 5852 35982 5854 36034
rect 5906 35982 6132 36034
rect 5852 35980 6132 35982
rect 6188 36596 6244 36606
rect 6188 36034 6244 36540
rect 8316 36596 8372 36606
rect 8316 36502 8372 36540
rect 11004 36596 11060 36606
rect 6188 35982 6190 36034
rect 6242 35982 6244 36034
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4172 34962 4228 34972
rect 5628 34916 5684 34926
rect 5628 34822 5684 34860
rect 4060 34626 4116 34636
rect 4620 34692 4676 34702
rect 4620 34578 4676 34636
rect 5516 34692 5572 34702
rect 4620 34526 4622 34578
rect 4674 34526 4676 34578
rect 4620 34514 4676 34526
rect 4956 34580 5012 34590
rect 4956 34486 5012 34524
rect 1820 34078 1822 34130
rect 1874 34078 1876 34130
rect 1820 34066 1876 34078
rect 2716 34132 2772 34142
rect 2716 34130 3332 34132
rect 2716 34078 2718 34130
rect 2770 34078 3332 34130
rect 2716 34076 3332 34078
rect 2716 34066 2772 34076
rect 2716 33794 2772 33806
rect 2716 33742 2718 33794
rect 2770 33742 2772 33794
rect 1820 33684 1876 33694
rect 2380 33684 2436 33694
rect 1820 33682 2436 33684
rect 1820 33630 1822 33682
rect 1874 33630 2382 33682
rect 2434 33630 2436 33682
rect 1820 33628 2436 33630
rect 1820 33618 1876 33628
rect 2268 31948 2324 33628
rect 2380 33618 2436 33628
rect 2716 33124 2772 33742
rect 3276 33794 3332 34076
rect 3276 33742 3278 33794
rect 3330 33742 3332 33794
rect 3276 33348 3332 33742
rect 5516 34018 5572 34636
rect 5852 34692 5908 35980
rect 6188 35970 6244 35982
rect 9772 36484 9828 36494
rect 9772 34802 9828 36428
rect 10780 35810 10836 35822
rect 10780 35758 10782 35810
rect 10834 35758 10836 35810
rect 10108 35586 10164 35598
rect 10108 35534 10110 35586
rect 10162 35534 10164 35586
rect 10108 35140 10164 35534
rect 10108 35084 10500 35140
rect 9772 34750 9774 34802
rect 9826 34750 9828 34802
rect 9772 34738 9828 34750
rect 10444 34802 10500 35084
rect 10444 34750 10446 34802
rect 10498 34750 10500 34802
rect 10444 34738 10500 34750
rect 5852 34626 5908 34636
rect 8540 34692 8596 34702
rect 8540 34598 8596 34636
rect 9324 34692 9380 34702
rect 5740 34580 5796 34590
rect 5740 34486 5796 34524
rect 8988 34580 9044 34590
rect 8988 34486 9044 34524
rect 9324 34578 9380 34636
rect 9884 34692 9940 34702
rect 9884 34598 9940 34636
rect 9324 34526 9326 34578
rect 9378 34526 9380 34578
rect 5516 33966 5518 34018
rect 5570 33966 5572 34018
rect 4284 33684 4340 33694
rect 3276 33292 3444 33348
rect 2716 33058 2772 33068
rect 3276 33124 3332 33134
rect 2268 31892 2996 31948
rect 2380 31890 2436 31892
rect 2380 31838 2382 31890
rect 2434 31838 2436 31890
rect 2380 31826 2436 31838
rect 2716 31778 2772 31790
rect 2716 31726 2718 31778
rect 2770 31726 2772 31778
rect 2380 30884 2436 30894
rect 1820 30770 1876 30782
rect 1820 30718 1822 30770
rect 1874 30718 1876 30770
rect 1820 30100 1876 30718
rect 2380 30770 2436 30828
rect 2716 30884 2772 31726
rect 2716 30818 2772 30828
rect 2380 30718 2382 30770
rect 2434 30718 2436 30770
rect 2380 30706 2436 30718
rect 1820 30034 1876 30044
rect 1932 29764 1988 29774
rect 1820 29650 1876 29662
rect 1820 29598 1822 29650
rect 1874 29598 1876 29650
rect 1820 27860 1876 29598
rect 1932 28978 1988 29708
rect 1932 28926 1934 28978
rect 1986 28926 1988 28978
rect 1932 28914 1988 28926
rect 2940 29650 2996 31892
rect 3276 31778 3332 33068
rect 3388 32788 3444 33292
rect 4284 33012 4340 33628
rect 4476 33292 4740 33302
rect 4532 33236 4580 33292
rect 4636 33236 4684 33292
rect 4476 33226 4740 33236
rect 4844 33124 4900 33134
rect 4844 33030 4900 33068
rect 4284 32956 4564 33012
rect 3388 32722 3444 32732
rect 4396 32788 4452 32798
rect 4396 32674 4452 32732
rect 4508 32786 4564 32956
rect 4508 32734 4510 32786
rect 4562 32734 4564 32786
rect 4508 32722 4564 32734
rect 4396 32622 4398 32674
rect 4450 32622 4452 32674
rect 4396 32610 4452 32622
rect 4956 32562 5012 32574
rect 4956 32510 4958 32562
rect 5010 32510 5012 32562
rect 4956 31892 5012 32510
rect 5516 32002 5572 33966
rect 5852 33684 5908 33694
rect 5852 33590 5908 33628
rect 5516 31950 5518 32002
rect 5570 31950 5572 32002
rect 5516 31948 5572 31950
rect 4956 31826 5012 31836
rect 5180 31892 5572 31948
rect 5852 31892 5908 31902
rect 3276 31726 3278 31778
rect 3330 31726 3332 31778
rect 3276 31714 3332 31726
rect 4476 31276 4740 31286
rect 4532 31220 4580 31276
rect 4636 31220 4684 31276
rect 4476 31210 4740 31220
rect 4620 30548 4676 30558
rect 4956 30548 5012 30558
rect 4620 30546 4900 30548
rect 4620 30494 4622 30546
rect 4674 30494 4900 30546
rect 4620 30492 4900 30494
rect 4620 30482 4676 30492
rect 4732 30324 4788 30334
rect 4844 30324 4900 30492
rect 4956 30454 5012 30492
rect 4844 30268 5124 30324
rect 3836 30100 3892 30110
rect 2940 29598 2942 29650
rect 2994 29598 2996 29650
rect 1820 27766 1876 27804
rect 2380 28530 2436 28542
rect 2380 28478 2382 28530
rect 2434 28478 2436 28530
rect 2380 27860 2436 28478
rect 2380 27794 2436 27804
rect 2940 27860 2996 29598
rect 3388 29762 3444 29774
rect 3388 29710 3390 29762
rect 3442 29710 3444 29762
rect 3388 29540 3444 29710
rect 3724 29764 3780 29774
rect 3724 29670 3780 29708
rect 3388 29474 3444 29484
rect 3276 29428 3332 29438
rect 3276 29334 3332 29372
rect 3836 28980 3892 30044
rect 4732 29986 4788 30268
rect 4732 29934 4734 29986
rect 4786 29934 4788 29986
rect 4732 29922 4788 29934
rect 5068 29988 5124 30268
rect 5180 29988 5236 31892
rect 5852 31798 5908 31836
rect 5628 30884 5684 30894
rect 5628 30790 5684 30828
rect 5740 30548 5796 30558
rect 5740 30454 5796 30492
rect 6076 30546 6132 30558
rect 6076 30494 6078 30546
rect 6130 30494 6132 30546
rect 6076 30324 6132 30494
rect 9324 30548 9380 34526
rect 10108 34580 10164 34590
rect 10108 34486 10164 34524
rect 9436 34468 9492 34478
rect 9436 34374 9492 34412
rect 10332 34468 10388 34478
rect 10332 33906 10388 34412
rect 10332 33854 10334 33906
rect 10386 33854 10388 33906
rect 10332 33842 10388 33854
rect 10780 33908 10836 35758
rect 11004 35812 11060 36540
rect 11340 35812 11396 37660
rect 13580 36932 13636 38558
rect 14364 38052 14420 40012
rect 16828 39956 16884 39966
rect 17836 39956 17892 42364
rect 17948 40852 18004 40862
rect 17948 40758 18004 40796
rect 16828 39954 17892 39956
rect 16828 39902 16830 39954
rect 16882 39902 17838 39954
rect 17890 39902 17892 39954
rect 16828 39900 17892 39902
rect 16828 39890 16884 39900
rect 17836 39890 17892 39900
rect 16492 39732 16548 39742
rect 16492 39638 16548 39676
rect 18060 39170 18116 43652
rect 19852 42866 19908 42878
rect 19852 42814 19854 42866
rect 19906 42814 19908 42866
rect 19852 42532 19908 42814
rect 19852 42466 19908 42476
rect 21420 42644 21476 42654
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 21420 42084 21476 42588
rect 21868 42642 21924 42654
rect 21868 42590 21870 42642
rect 21922 42590 21924 42642
rect 21868 42530 21924 42590
rect 22204 42644 22260 43820
rect 22652 44658 22708 44670
rect 22652 44606 22654 44658
rect 22706 44606 22708 44658
rect 22540 43764 22596 43774
rect 22652 43764 22708 44606
rect 22988 44660 23044 45166
rect 23436 44884 23492 44894
rect 23100 44660 23156 44670
rect 22988 44658 23156 44660
rect 22988 44606 23102 44658
rect 23154 44606 23156 44658
rect 22988 44604 23156 44606
rect 22596 43708 22708 43764
rect 22540 43540 22596 43708
rect 22316 42756 22372 42766
rect 22316 42662 22372 42700
rect 22540 42754 22596 43484
rect 23100 43652 23156 44604
rect 23436 43708 23492 44828
rect 23996 44882 24052 44894
rect 23996 44830 23998 44882
rect 24050 44830 24052 44882
rect 23996 44100 24052 44830
rect 23996 44034 24052 44044
rect 24668 44100 24724 44110
rect 23884 43764 23940 43774
rect 23436 43652 23828 43708
rect 22540 42702 22542 42754
rect 22594 42702 22596 42754
rect 22204 42578 22260 42588
rect 21868 42478 21870 42530
rect 21922 42478 21924 42530
rect 21868 42466 21924 42478
rect 22428 42532 22484 42542
rect 22540 42532 22596 42702
rect 22764 42754 22820 42766
rect 22764 42702 22766 42754
rect 22818 42702 22820 42754
rect 22764 42644 22820 42702
rect 23100 42756 23156 43596
rect 23772 42866 23828 43652
rect 23884 43540 23940 43708
rect 24668 43652 24724 44044
rect 25788 43708 25844 46622
rect 26012 46676 26068 47740
rect 26572 47906 26628 47918
rect 26572 47854 26574 47906
rect 26626 47854 26628 47906
rect 26572 47796 26628 47854
rect 26572 47124 26628 47740
rect 26572 47058 26628 47068
rect 27580 47012 27636 47022
rect 26348 46676 26404 46686
rect 26012 46674 26404 46676
rect 26012 46622 26350 46674
rect 26402 46622 26404 46674
rect 26012 46620 26404 46622
rect 26348 46004 26404 46620
rect 27580 46674 27636 46956
rect 27580 46622 27582 46674
rect 27634 46622 27636 46674
rect 27580 46004 27636 46622
rect 26348 45948 26628 46004
rect 26460 45780 26516 45790
rect 26348 44884 26404 44894
rect 26460 44884 26516 45724
rect 26572 45666 26628 45948
rect 27580 45938 27636 45948
rect 27804 46676 27860 46686
rect 27804 46114 27860 46620
rect 27804 46062 27806 46114
rect 27858 46062 27860 46114
rect 26572 45614 26574 45666
rect 26626 45614 26628 45666
rect 26572 45602 26628 45614
rect 26908 45778 26964 45790
rect 26908 45726 26910 45778
rect 26962 45726 26964 45778
rect 26908 45666 26964 45726
rect 26908 45614 26910 45666
rect 26962 45614 26964 45666
rect 26908 45602 26964 45614
rect 27356 45778 27412 45790
rect 27356 45726 27358 45778
rect 27410 45726 27412 45778
rect 27356 45666 27412 45726
rect 27356 45614 27358 45666
rect 27410 45614 27412 45666
rect 27356 45602 27412 45614
rect 26684 44884 26740 44894
rect 26460 44882 26740 44884
rect 26460 44830 26686 44882
rect 26738 44830 26740 44882
rect 26460 44828 26740 44830
rect 26348 44790 26404 44828
rect 26684 43764 26740 44828
rect 27804 44884 27860 46062
rect 27804 44818 27860 44828
rect 28140 45890 28196 45902
rect 28140 45838 28142 45890
rect 28194 45838 28196 45890
rect 28140 45666 28196 45838
rect 28140 45614 28142 45666
rect 28194 45614 28196 45666
rect 28140 44884 28196 45614
rect 27804 44546 27860 44558
rect 27804 44494 27806 44546
rect 27858 44494 27860 44546
rect 27244 44100 27300 44110
rect 27244 44006 27300 44044
rect 27692 43988 27748 43998
rect 27692 43708 27748 43932
rect 25788 43652 26516 43708
rect 26684 43698 26740 43708
rect 24668 43586 24724 43596
rect 23884 43474 23940 43484
rect 23772 42814 23774 42866
rect 23826 42814 23828 42866
rect 23100 42690 23156 42700
rect 23436 42756 23492 42766
rect 23492 42700 23604 42756
rect 23436 42662 23492 42700
rect 22764 42578 22820 42588
rect 22428 42530 22596 42532
rect 22428 42478 22430 42530
rect 22482 42478 22596 42530
rect 22428 42476 22596 42478
rect 22428 42466 22484 42476
rect 21868 42140 22148 42196
rect 21476 42028 21812 42084
rect 21420 41990 21476 42028
rect 18508 41972 18564 41982
rect 18508 41858 18564 41916
rect 20524 41972 20580 41982
rect 20524 41878 20580 41916
rect 18508 41806 18510 41858
rect 18562 41806 18564 41858
rect 18508 41794 18564 41806
rect 21308 41858 21364 41870
rect 21308 41806 21310 41858
rect 21362 41806 21364 41858
rect 18172 41746 18228 41758
rect 18172 41694 18174 41746
rect 18226 41694 18228 41746
rect 18172 40852 18228 41694
rect 21308 41076 21364 41806
rect 21756 41524 21812 42028
rect 21868 41970 21924 42140
rect 21868 41918 21870 41970
rect 21922 41918 21924 41970
rect 21868 41906 21924 41918
rect 21980 41972 22036 41982
rect 21756 41468 21924 41524
rect 21308 40982 21364 41020
rect 18172 40786 18228 40796
rect 18956 40852 19012 40862
rect 18732 40628 18788 40638
rect 18732 40626 18900 40628
rect 18732 40574 18734 40626
rect 18786 40574 18900 40626
rect 18732 40572 18900 40574
rect 18732 40562 18788 40572
rect 18060 39118 18062 39170
rect 18114 39118 18116 39170
rect 18060 39106 18116 39118
rect 18396 39954 18452 39966
rect 18396 39902 18398 39954
rect 18450 39902 18452 39954
rect 18396 39732 18452 39902
rect 17388 39060 17444 39070
rect 17388 38948 17444 39004
rect 18396 38948 18452 39676
rect 18508 39732 18564 39742
rect 18508 39730 18788 39732
rect 18508 39678 18510 39730
rect 18562 39678 18788 39730
rect 18508 39676 18788 39678
rect 18508 39666 18564 39676
rect 18732 39060 18788 39676
rect 17388 38946 17556 38948
rect 17388 38894 17390 38946
rect 17442 38894 17556 38946
rect 17388 38892 17556 38894
rect 18396 38892 18676 38948
rect 17388 38882 17444 38892
rect 16604 38722 16660 38734
rect 16604 38670 16606 38722
rect 16658 38670 16660 38722
rect 16604 38668 16660 38670
rect 16604 38612 16884 38668
rect 14364 38050 14756 38052
rect 14364 37998 14366 38050
rect 14418 37998 14756 38050
rect 14364 37996 14756 37998
rect 14364 37986 14420 37996
rect 13580 36866 13636 36876
rect 14700 36930 14756 37996
rect 16828 37716 16884 38556
rect 17052 38610 17108 38622
rect 17052 38558 17054 38610
rect 17106 38558 17108 38610
rect 17052 38052 17108 38558
rect 17052 37986 17108 37996
rect 17500 38050 17556 38892
rect 17836 38724 17892 38734
rect 17836 38630 17892 38668
rect 18508 38724 18564 38734
rect 18508 38630 18564 38668
rect 17500 37998 17502 38050
rect 17554 37998 17556 38050
rect 17500 37940 17556 37998
rect 17948 38052 18004 38062
rect 17948 37958 18004 37996
rect 17500 37874 17556 37884
rect 18396 37828 18452 37838
rect 18396 37734 18452 37772
rect 16828 37622 16884 37660
rect 14700 36878 14702 36930
rect 14754 36878 14756 36930
rect 14700 36820 14756 36878
rect 14700 36754 14756 36764
rect 14812 37602 14868 37614
rect 14812 37550 14814 37602
rect 14866 37550 14868 37602
rect 14812 36932 14868 37550
rect 13580 36594 13636 36606
rect 13580 36542 13582 36594
rect 13634 36542 13636 36594
rect 13468 36484 13524 36494
rect 13468 36390 13524 36428
rect 12124 35924 12180 35934
rect 12124 35830 12180 35868
rect 11004 35810 11396 35812
rect 11004 35758 11342 35810
rect 11394 35758 11396 35810
rect 11004 35756 11396 35758
rect 11340 35746 11396 35756
rect 10892 35698 10948 35710
rect 10892 35646 10894 35698
rect 10946 35646 10948 35698
rect 10892 34132 10948 35646
rect 13580 35026 13636 36542
rect 14812 36260 14868 36876
rect 15036 36820 15092 36830
rect 15036 36726 15092 36764
rect 15484 36820 15540 36830
rect 14812 36204 15204 36260
rect 14476 35924 14532 35934
rect 14476 35830 14532 35868
rect 14588 35812 14644 35822
rect 14588 35718 14644 35756
rect 14140 35588 14196 35598
rect 13580 34974 13582 35026
rect 13634 34974 13636 35026
rect 13580 34962 13636 34974
rect 13692 35586 14196 35588
rect 13692 35534 14142 35586
rect 14194 35534 14196 35586
rect 13692 35532 14196 35534
rect 13468 34802 13524 34814
rect 13468 34750 13470 34802
rect 13522 34750 13524 34802
rect 12124 34692 12180 34702
rect 12124 34598 12180 34636
rect 13468 34692 13524 34750
rect 13468 34626 13524 34636
rect 13692 34802 13748 35532
rect 14140 35522 14196 35532
rect 13692 34750 13694 34802
rect 13746 34750 13748 34802
rect 10892 34066 10948 34076
rect 11900 34468 11956 34478
rect 11004 33908 11060 33918
rect 10780 33906 11060 33908
rect 10780 33854 11006 33906
rect 11058 33854 11060 33906
rect 10780 33852 11060 33854
rect 11004 33572 11060 33852
rect 11004 33506 11060 33516
rect 11900 32786 11956 34412
rect 12908 34468 12964 34478
rect 12572 34356 12628 34366
rect 12124 34132 12180 34142
rect 12124 34038 12180 34076
rect 12572 34130 12628 34300
rect 12572 34078 12574 34130
rect 12626 34078 12628 34130
rect 12572 34066 12628 34078
rect 12908 33684 12964 34412
rect 13020 34132 13076 34142
rect 13020 33906 13076 34076
rect 13020 33854 13022 33906
rect 13074 33854 13076 33906
rect 13020 33842 13076 33854
rect 13580 33908 13636 33918
rect 13580 33814 13636 33852
rect 13692 33908 13748 34750
rect 15036 34020 15092 34030
rect 14364 33964 14756 34020
rect 14140 33908 14196 33918
rect 14364 33908 14420 33964
rect 13692 33906 14420 33908
rect 13692 33854 13694 33906
rect 13746 33854 14142 33906
rect 14194 33854 14420 33906
rect 13692 33852 14420 33854
rect 14700 33906 14756 33964
rect 15036 33926 15092 33964
rect 14700 33854 14702 33906
rect 14754 33854 14756 33906
rect 13692 33842 13748 33852
rect 12908 33618 12964 33628
rect 12460 33572 12516 33582
rect 12460 33010 12516 33516
rect 12460 32958 12462 33010
rect 12514 32958 12516 33010
rect 12460 32946 12516 32958
rect 11900 32734 11902 32786
rect 11954 32734 11956 32786
rect 11900 32722 11956 32734
rect 12796 32674 12852 32686
rect 12796 32622 12798 32674
rect 12850 32622 12852 32674
rect 12796 32564 12852 32622
rect 14140 32674 14196 33852
rect 14700 33842 14756 33854
rect 14476 33796 14532 33806
rect 14476 33702 14532 33740
rect 14364 33684 14420 33694
rect 14364 33590 14420 33628
rect 14700 33012 14756 33022
rect 14700 32918 14756 32956
rect 14588 32788 14644 32798
rect 14140 32622 14142 32674
rect 14194 32622 14196 32674
rect 14140 32610 14196 32622
rect 14476 32732 14588 32788
rect 12796 32498 12852 32508
rect 14476 32562 14532 32732
rect 14476 32510 14478 32562
rect 14530 32510 14532 32562
rect 14476 32498 14532 32510
rect 10780 32452 10836 32462
rect 10780 31778 10836 32396
rect 11788 32452 11844 32462
rect 11788 32358 11844 32396
rect 13468 32002 13524 32014
rect 13468 31950 13470 32002
rect 13522 31950 13524 32002
rect 11340 31892 11396 31902
rect 11340 31780 11396 31836
rect 10780 31726 10782 31778
rect 10834 31726 10836 31778
rect 10780 31714 10836 31726
rect 10892 31778 11396 31780
rect 10892 31726 11342 31778
rect 11394 31726 11396 31778
rect 10892 31724 11396 31726
rect 10444 31666 10500 31678
rect 10444 31614 10446 31666
rect 10498 31614 10500 31666
rect 6076 30258 6132 30268
rect 6188 30434 6244 30446
rect 6188 30382 6190 30434
rect 6242 30382 6244 30434
rect 5068 29986 5236 29988
rect 5068 29934 5182 29986
rect 5234 29934 5236 29986
rect 5068 29932 5236 29934
rect 4172 29764 4228 29774
rect 3836 28914 3892 28924
rect 3948 29762 4228 29764
rect 3948 29710 4174 29762
rect 4226 29710 4228 29762
rect 3948 29708 4228 29710
rect 3836 27972 3892 27982
rect 3948 27972 4004 29708
rect 4172 29698 4228 29708
rect 4284 29426 4340 29438
rect 4284 29374 4286 29426
rect 4338 29374 4340 29426
rect 4284 29092 4340 29374
rect 5068 29428 5124 29438
rect 4476 29260 4740 29270
rect 4532 29204 4580 29260
rect 4636 29204 4684 29260
rect 4476 29194 4740 29204
rect 4284 29026 4340 29036
rect 4508 28980 4564 28990
rect 4508 28754 4564 28924
rect 4508 28702 4510 28754
rect 4562 28702 4564 28754
rect 4508 28690 4564 28702
rect 5068 28756 5124 29372
rect 5068 28662 5124 28700
rect 3836 27970 4004 27972
rect 3836 27918 3838 27970
rect 3890 27918 4004 27970
rect 3836 27916 4004 27918
rect 4284 27970 4340 27982
rect 4284 27918 4286 27970
rect 4338 27918 4340 27970
rect 3836 27906 3892 27916
rect 2940 27794 2996 27804
rect 3388 27860 3444 27870
rect 3388 27766 3444 27804
rect 4284 27860 4340 27918
rect 4284 27794 4340 27804
rect 5068 27860 5124 27870
rect 5180 27860 5236 29932
rect 6188 29876 6244 30382
rect 6188 29810 6244 29820
rect 6748 30436 6804 30446
rect 5516 29092 5572 29102
rect 5572 29036 5684 29092
rect 5516 29026 5572 29036
rect 5628 28754 5684 29036
rect 6748 28980 6804 30380
rect 8540 29988 8596 29998
rect 8540 29894 8596 29932
rect 9324 29988 9380 30492
rect 9660 30770 9716 30782
rect 10220 30772 10276 30782
rect 9660 30718 9662 30770
rect 9714 30718 9716 30770
rect 9660 30100 9716 30718
rect 9660 30034 9716 30044
rect 9884 30770 10276 30772
rect 9884 30718 10222 30770
rect 10274 30718 10276 30770
rect 9884 30716 10276 30718
rect 6748 28914 6804 28924
rect 6972 29876 7028 29886
rect 5628 28702 5630 28754
rect 5682 28702 5684 28754
rect 5628 28082 5684 28702
rect 6188 28756 6244 28766
rect 6188 28662 6244 28700
rect 5628 28030 5630 28082
rect 5682 28030 5684 28082
rect 5628 28018 5684 28030
rect 6300 28084 6356 28094
rect 6300 28082 6468 28084
rect 6300 28030 6302 28082
rect 6354 28030 6468 28082
rect 6300 28028 6468 28030
rect 6300 28018 6356 28028
rect 5124 27804 5236 27860
rect 5740 27860 5796 27870
rect 5068 27794 5124 27804
rect 4476 27244 4740 27254
rect 4532 27188 4580 27244
rect 4636 27188 4684 27244
rect 4476 27178 4740 27188
rect 5740 26850 5796 27804
rect 6412 27746 6468 28028
rect 6412 27694 6414 27746
rect 6466 27694 6468 27746
rect 6412 27682 6468 27694
rect 6972 27746 7028 29820
rect 7308 29876 7364 29886
rect 7308 29762 7364 29820
rect 7308 29710 7310 29762
rect 7362 29710 7364 29762
rect 7308 29698 7364 29710
rect 7868 29762 7924 29774
rect 7868 29710 7870 29762
rect 7922 29710 7924 29762
rect 7868 29428 7924 29710
rect 8988 29762 9044 29774
rect 8988 29710 8990 29762
rect 9042 29710 9044 29762
rect 7868 29362 7924 29372
rect 8764 29540 8820 29550
rect 8764 28978 8820 29484
rect 8876 29428 8932 29438
rect 8876 29334 8932 29372
rect 8764 28926 8766 28978
rect 8818 28926 8820 28978
rect 8764 28914 8820 28926
rect 8988 28644 9044 29710
rect 9324 28868 9380 29932
rect 9884 29426 9940 30716
rect 10220 30706 10276 30716
rect 10444 30548 10500 31614
rect 10444 30482 10500 30492
rect 10332 30100 10388 30110
rect 10220 30044 10332 30100
rect 9996 29764 10052 29774
rect 9996 29670 10052 29708
rect 9884 29374 9886 29426
rect 9938 29374 9940 29426
rect 8988 28578 9044 28588
rect 9100 28866 9380 28868
rect 9100 28814 9326 28866
rect 9378 28814 9380 28866
rect 9100 28812 9380 28814
rect 8428 28532 8484 28542
rect 8428 28438 8484 28476
rect 9100 28532 9156 28812
rect 9324 28802 9380 28812
rect 9660 29092 9716 29102
rect 9660 28754 9716 29036
rect 9660 28702 9662 28754
rect 9714 28702 9716 28754
rect 9660 28690 9716 28702
rect 8988 27972 9044 27982
rect 9100 27972 9156 28476
rect 8988 27970 9156 27972
rect 8988 27918 8990 27970
rect 9042 27918 9156 27970
rect 8988 27916 9156 27918
rect 8988 27906 9044 27916
rect 6972 27694 6974 27746
rect 7026 27694 7028 27746
rect 6972 27682 7028 27694
rect 9660 27748 9716 27758
rect 9884 27748 9940 29374
rect 9660 27746 9940 27748
rect 9660 27694 9662 27746
rect 9714 27694 9940 27746
rect 9660 27692 9940 27694
rect 10108 29428 10164 29438
rect 10108 27748 10164 29372
rect 10220 28754 10276 30044
rect 10332 30006 10388 30044
rect 10444 29762 10500 29774
rect 10444 29710 10446 29762
rect 10498 29710 10500 29762
rect 10444 28980 10500 29710
rect 10780 29764 10836 29774
rect 10892 29764 10948 31724
rect 11340 31714 11396 31724
rect 13468 31332 13524 31950
rect 14364 31892 14420 31902
rect 14364 31798 14420 31836
rect 13916 31780 13972 31790
rect 13916 31686 13972 31724
rect 14476 31780 14532 31790
rect 14476 31686 14532 31724
rect 12460 30548 12516 30558
rect 10780 29762 10948 29764
rect 10780 29710 10782 29762
rect 10834 29710 10948 29762
rect 10780 29708 10948 29710
rect 11340 29762 11396 29774
rect 11340 29710 11342 29762
rect 11394 29710 11396 29762
rect 10780 29698 10836 29708
rect 11340 29092 11396 29710
rect 11340 29026 11396 29036
rect 10444 28914 10500 28924
rect 10220 28702 10222 28754
rect 10274 28702 10276 28754
rect 10220 28690 10276 28702
rect 12460 28530 12516 30492
rect 12796 30548 12852 30558
rect 13468 30548 13524 31276
rect 14588 30772 14644 32732
rect 15148 32786 15204 36204
rect 15484 34916 15540 36764
rect 17836 36818 17892 36830
rect 17836 36766 17838 36818
rect 17890 36766 17892 36818
rect 17836 36708 17892 36766
rect 15820 36596 15876 36606
rect 15820 36502 15876 36540
rect 16604 35476 16660 35486
rect 16156 34916 16212 34926
rect 15484 34914 15876 34916
rect 15484 34862 15486 34914
rect 15538 34862 15876 34914
rect 15484 34860 15876 34862
rect 15484 34850 15540 34860
rect 15820 34802 15876 34860
rect 15820 34750 15822 34802
rect 15874 34750 15876 34802
rect 15820 34738 15876 34750
rect 16156 34020 16212 34860
rect 16604 34690 16660 35420
rect 17836 35364 17892 36652
rect 18508 36708 18564 36718
rect 18508 36614 18564 36652
rect 18060 36596 18116 36606
rect 18060 36502 18116 36540
rect 18620 35924 18676 38892
rect 18732 38834 18788 39004
rect 18732 38782 18734 38834
rect 18786 38782 18788 38834
rect 18732 38770 18788 38782
rect 18844 38162 18900 40572
rect 18956 39842 19012 40796
rect 20188 40852 20244 40862
rect 19836 40348 20100 40358
rect 19892 40292 19940 40348
rect 19996 40292 20044 40348
rect 19836 40282 20100 40292
rect 19740 39956 19796 39966
rect 18956 39790 18958 39842
rect 19010 39790 19012 39842
rect 18956 39778 19012 39790
rect 19516 39954 19796 39956
rect 19516 39902 19742 39954
rect 19794 39902 19796 39954
rect 19516 39900 19796 39902
rect 19516 39170 19572 39900
rect 19740 39890 19796 39900
rect 19516 39118 19518 39170
rect 19570 39118 19572 39170
rect 19516 39106 19572 39118
rect 19964 38836 20020 38846
rect 19964 38742 20020 38780
rect 18956 38722 19012 38734
rect 18956 38670 18958 38722
rect 19010 38670 19012 38722
rect 18956 38668 19012 38670
rect 18956 38612 19124 38668
rect 18844 38110 18846 38162
rect 18898 38110 18900 38162
rect 18844 38098 18900 38110
rect 19068 38052 19124 38612
rect 19836 38332 20100 38342
rect 19892 38276 19940 38332
rect 19996 38276 20044 38332
rect 19836 38266 20100 38276
rect 19404 38162 19460 38174
rect 19404 38110 19406 38162
rect 19458 38110 19460 38162
rect 19404 38052 19460 38110
rect 19516 38052 19572 38062
rect 19404 38050 19572 38052
rect 19404 37998 19518 38050
rect 19570 37998 19572 38050
rect 19404 37996 19572 37998
rect 18844 37714 18900 37726
rect 18844 37662 18846 37714
rect 18898 37662 18900 37714
rect 18844 37044 18900 37662
rect 18844 36978 18900 36988
rect 19068 36820 19124 37996
rect 19516 37986 19572 37996
rect 19404 37828 19460 37838
rect 19404 37734 19460 37772
rect 19964 37828 20020 37838
rect 20188 37828 20244 40796
rect 20748 40852 20804 40862
rect 20748 40758 20804 40796
rect 21420 40626 21476 40638
rect 21420 40574 21422 40626
rect 21474 40574 21476 40626
rect 21420 40516 21476 40574
rect 21420 40068 21476 40460
rect 21868 40626 21924 41468
rect 21868 40574 21870 40626
rect 21922 40574 21924 40626
rect 21868 40514 21924 40574
rect 21868 40462 21870 40514
rect 21922 40462 21924 40514
rect 21868 40450 21924 40462
rect 21980 40178 22036 41916
rect 21980 40126 21982 40178
rect 22034 40126 22036 40178
rect 21980 40114 22036 40126
rect 21420 40012 21812 40068
rect 21644 39844 21700 39854
rect 20412 39060 20468 39070
rect 20020 37772 20244 37828
rect 20300 39004 20412 39060
rect 20300 37826 20356 39004
rect 20412 38994 20468 39004
rect 21644 39060 21700 39788
rect 21756 39620 21812 40012
rect 21756 39618 21924 39620
rect 21756 39566 21758 39618
rect 21810 39566 21924 39618
rect 21756 39564 21924 39566
rect 21756 39554 21812 39564
rect 21644 38966 21700 39004
rect 21868 38836 21924 39564
rect 20412 38722 20468 38734
rect 20412 38670 20414 38722
rect 20466 38670 20468 38722
rect 20412 38612 20468 38670
rect 20636 38724 20692 38734
rect 21308 38724 21364 38734
rect 20636 38722 21364 38724
rect 20636 38670 20638 38722
rect 20690 38670 21310 38722
rect 21362 38670 21364 38722
rect 20636 38668 21364 38670
rect 20636 38658 20692 38668
rect 20412 38546 20468 38556
rect 20412 37940 20468 37950
rect 20412 37846 20468 37884
rect 20300 37774 20302 37826
rect 20354 37774 20356 37826
rect 19964 37734 20020 37772
rect 20300 37762 20356 37774
rect 20636 37828 20692 37838
rect 19964 37044 20020 37054
rect 19068 36706 19124 36764
rect 19068 36654 19070 36706
rect 19122 36654 19124 36706
rect 19068 36642 19124 36654
rect 19180 36932 19236 36942
rect 18956 35924 19012 35934
rect 18620 35922 19012 35924
rect 18620 35870 18958 35922
rect 19010 35870 19012 35922
rect 18620 35868 19012 35870
rect 18396 35810 18452 35822
rect 18396 35758 18398 35810
rect 18450 35758 18452 35810
rect 17948 35476 18004 35486
rect 17948 35382 18004 35420
rect 16604 34638 16606 34690
rect 16658 34638 16660 34690
rect 16604 34626 16660 34638
rect 17500 35308 17892 35364
rect 16156 33906 16212 33964
rect 16156 33854 16158 33906
rect 16210 33854 16212 33906
rect 15932 33796 15988 33806
rect 15932 33702 15988 33740
rect 16044 33458 16100 33470
rect 16044 33406 16046 33458
rect 16098 33406 16100 33458
rect 15708 32900 15764 32910
rect 15148 32734 15150 32786
rect 15202 32734 15204 32786
rect 15148 32722 15204 32734
rect 15372 32788 15428 32798
rect 15372 32694 15428 32732
rect 15708 32674 15764 32844
rect 15708 32622 15710 32674
rect 15762 32622 15764 32674
rect 15708 32610 15764 32622
rect 16044 32340 16100 33406
rect 16044 32274 16100 32284
rect 15932 31890 15988 31902
rect 15932 31838 15934 31890
rect 15986 31838 15988 31890
rect 15372 31780 15428 31790
rect 15372 31686 15428 31724
rect 14924 31668 14980 31678
rect 14924 31574 14980 31612
rect 15932 31108 15988 31838
rect 16044 31892 16100 31902
rect 16156 31892 16212 33854
rect 16044 31890 16212 31892
rect 16044 31838 16046 31890
rect 16098 31838 16212 31890
rect 16044 31836 16212 31838
rect 16044 31826 16100 31836
rect 15932 31042 15988 31052
rect 15036 30996 15092 31006
rect 15036 30902 15092 30940
rect 16156 30882 16212 31836
rect 16380 33794 16436 33806
rect 16380 33742 16382 33794
rect 16434 33742 16436 33794
rect 16380 31780 16436 33742
rect 17276 32788 17332 32798
rect 17500 32788 17556 35308
rect 18396 34804 18452 35758
rect 18956 35364 19012 35868
rect 19068 35924 19124 35934
rect 19180 35924 19236 36876
rect 19964 36708 20020 36988
rect 20412 37044 20468 37054
rect 20076 36932 20132 36942
rect 20132 36876 20244 36932
rect 20076 36866 20132 36876
rect 20076 36708 20132 36718
rect 19964 36706 20132 36708
rect 19964 36654 20078 36706
rect 20130 36654 20132 36706
rect 19964 36652 20132 36654
rect 20076 36642 20132 36652
rect 19836 36316 20100 36326
rect 19892 36260 19940 36316
rect 19996 36260 20044 36316
rect 19836 36250 20100 36260
rect 20076 36148 20132 36158
rect 19964 36092 20076 36148
rect 19068 35922 19236 35924
rect 19068 35870 19070 35922
rect 19122 35870 19236 35922
rect 19068 35868 19236 35870
rect 19740 35924 19796 35934
rect 19068 35858 19124 35868
rect 19740 35830 19796 35868
rect 18956 35298 19012 35308
rect 19516 35810 19572 35822
rect 19516 35758 19518 35810
rect 19570 35758 19572 35810
rect 19180 35028 19236 35038
rect 19180 34914 19236 34972
rect 19180 34862 19182 34914
rect 19234 34862 19236 34914
rect 19180 34850 19236 34862
rect 19516 34916 19572 35758
rect 19628 35812 19684 35822
rect 19628 35718 19684 35756
rect 19964 35810 20020 36092
rect 20076 36082 20132 36092
rect 19964 35758 19966 35810
rect 20018 35758 20020 35810
rect 19964 35746 20020 35758
rect 19516 34850 19572 34860
rect 18620 34804 18676 34814
rect 18396 34802 18676 34804
rect 18396 34750 18622 34802
rect 18674 34750 18676 34802
rect 18396 34748 18676 34750
rect 18396 33796 18452 33806
rect 17948 33460 18004 33470
rect 17276 32786 17556 32788
rect 17276 32734 17278 32786
rect 17330 32734 17556 32786
rect 17276 32732 17556 32734
rect 17612 33458 18004 33460
rect 17612 33406 17950 33458
rect 18002 33406 18004 33458
rect 17612 33404 18004 33406
rect 17612 32786 17668 33404
rect 17948 33394 18004 33404
rect 17612 32734 17614 32786
rect 17666 32734 17668 32786
rect 17276 32722 17332 32732
rect 17612 32722 17668 32734
rect 18396 32788 18452 33740
rect 18396 32722 18452 32732
rect 18508 32786 18564 34748
rect 18620 34738 18676 34748
rect 20188 34802 20244 36876
rect 20412 36818 20468 36988
rect 20412 36766 20414 36818
rect 20466 36766 20468 36818
rect 20412 36754 20468 36766
rect 20524 35698 20580 35710
rect 20524 35646 20526 35698
rect 20578 35646 20580 35698
rect 20524 35364 20580 35646
rect 20524 35298 20580 35308
rect 20188 34750 20190 34802
rect 20242 34750 20244 34802
rect 20188 34738 20244 34750
rect 20300 35028 20356 35038
rect 19852 34692 19908 34702
rect 19292 34690 19908 34692
rect 19292 34638 19854 34690
rect 19906 34638 19908 34690
rect 19292 34636 19908 34638
rect 18956 33906 19012 33918
rect 18956 33854 18958 33906
rect 19010 33854 19012 33906
rect 18956 32900 19012 33854
rect 19068 33908 19124 33918
rect 19292 33908 19348 34636
rect 19852 34626 19908 34636
rect 20300 34690 20356 34972
rect 20300 34638 20302 34690
rect 20354 34638 20356 34690
rect 20300 34626 20356 34638
rect 19404 34468 19460 34478
rect 19404 34466 19684 34468
rect 19404 34414 19406 34466
rect 19458 34414 19684 34466
rect 19404 34412 19684 34414
rect 19404 34402 19460 34412
rect 19068 33906 19348 33908
rect 19068 33854 19070 33906
rect 19122 33854 19348 33906
rect 19068 33852 19348 33854
rect 19068 33842 19124 33852
rect 18956 32834 19012 32844
rect 19292 33012 19348 33852
rect 18508 32734 18510 32786
rect 18562 32734 18564 32786
rect 18508 32722 18564 32734
rect 16940 32676 16996 32686
rect 19068 32676 19124 32686
rect 16940 32674 17220 32676
rect 16940 32622 16942 32674
rect 16994 32622 17220 32674
rect 16940 32620 17220 32622
rect 16940 32610 16996 32620
rect 16380 31714 16436 31724
rect 16828 31666 16884 31678
rect 16828 31614 16830 31666
rect 16882 31614 16884 31666
rect 16828 31332 16884 31614
rect 16828 31266 16884 31276
rect 17164 31108 17220 32620
rect 18732 32674 19124 32676
rect 18732 32622 19070 32674
rect 19122 32622 19124 32674
rect 18732 32620 19124 32622
rect 17948 32564 18004 32574
rect 17948 32470 18004 32508
rect 17724 31556 17780 31566
rect 17836 31556 17892 31566
rect 17724 31554 17836 31556
rect 17724 31502 17726 31554
rect 17778 31502 17836 31554
rect 17724 31500 17836 31502
rect 17724 31490 17780 31500
rect 17276 31108 17332 31118
rect 17164 31106 17332 31108
rect 17164 31054 17278 31106
rect 17330 31054 17332 31106
rect 17164 31052 17332 31054
rect 17276 31042 17332 31052
rect 16156 30830 16158 30882
rect 16210 30830 16212 30882
rect 16156 30818 16212 30830
rect 17836 30772 17892 31500
rect 18732 31106 18788 32620
rect 19068 32610 19124 32620
rect 18732 31054 18734 31106
rect 18786 31054 18788 31106
rect 18732 31042 18788 31054
rect 19180 30884 19236 30894
rect 17948 30772 18004 30782
rect 14588 30770 14980 30772
rect 14588 30718 14590 30770
rect 14642 30718 14980 30770
rect 14588 30716 14980 30718
rect 17836 30770 18004 30772
rect 17836 30718 17950 30770
rect 18002 30718 18004 30770
rect 17836 30716 18004 30718
rect 14588 30706 14644 30716
rect 12796 30546 12964 30548
rect 12796 30494 12798 30546
rect 12850 30494 12964 30546
rect 12796 30492 12964 30494
rect 12796 30482 12852 30492
rect 12908 29764 12964 30492
rect 13468 29986 13524 30492
rect 13916 30660 13972 30670
rect 13580 30436 13636 30446
rect 13580 30342 13636 30380
rect 13916 29988 13972 30604
rect 13468 29934 13470 29986
rect 13522 29934 13524 29986
rect 13468 29922 13524 29934
rect 13580 29986 13972 29988
rect 13580 29934 13918 29986
rect 13970 29934 13972 29986
rect 13580 29932 13972 29934
rect 12796 28980 12852 28990
rect 12796 28886 12852 28924
rect 12908 28756 12964 29708
rect 13468 29092 13524 29102
rect 13468 28998 13524 29036
rect 12908 28690 12964 28700
rect 13580 28754 13636 29932
rect 13916 29922 13972 29932
rect 14028 30658 14084 30670
rect 14028 30606 14030 30658
rect 14082 30606 14084 30658
rect 13580 28702 13582 28754
rect 13634 28702 13636 28754
rect 13580 28690 13636 28702
rect 13916 29652 13972 29662
rect 13916 28756 13972 29596
rect 14028 28980 14084 30606
rect 14476 30658 14532 30670
rect 14476 30606 14478 30658
rect 14530 30606 14532 30658
rect 14476 30548 14532 30606
rect 14588 30548 14644 30558
rect 14476 30492 14588 30548
rect 14588 30482 14644 30492
rect 14252 30212 14308 30222
rect 14252 30098 14308 30156
rect 14252 30046 14254 30098
rect 14306 30046 14308 30098
rect 14252 30034 14308 30046
rect 14028 28914 14084 28924
rect 14700 29762 14756 29774
rect 14700 29710 14702 29762
rect 14754 29710 14756 29762
rect 14028 28756 14084 28766
rect 13916 28754 14084 28756
rect 13916 28702 14030 28754
rect 14082 28702 14084 28754
rect 13916 28700 14084 28702
rect 14028 28690 14084 28700
rect 14476 28756 14532 28766
rect 14476 28662 14532 28700
rect 12460 28478 12462 28530
rect 12514 28478 12516 28530
rect 12460 27970 12516 28478
rect 12460 27918 12462 27970
rect 12514 27918 12516 27970
rect 12460 27906 12516 27918
rect 12796 28644 12852 28654
rect 12796 27970 12852 28588
rect 14700 28644 14756 29710
rect 14924 29764 14980 30716
rect 17948 30706 18004 30716
rect 19180 30770 19236 30828
rect 19180 30718 19182 30770
rect 19234 30718 19236 30770
rect 15484 30660 15540 30670
rect 15484 30566 15540 30604
rect 16044 30658 16100 30670
rect 16044 30606 16046 30658
rect 16098 30606 16100 30658
rect 16044 30436 16100 30606
rect 16044 30370 16100 30380
rect 17724 30658 17780 30670
rect 17724 30606 17726 30658
rect 17778 30606 17780 30658
rect 17724 30548 17780 30606
rect 17724 30100 17780 30492
rect 18284 30658 18340 30670
rect 18284 30606 18286 30658
rect 18338 30606 18340 30658
rect 18284 30436 18340 30606
rect 18284 30370 18340 30380
rect 17724 30034 17780 30044
rect 15260 29876 15316 29886
rect 15260 29782 15316 29820
rect 19180 29876 19236 30718
rect 19292 30772 19348 32956
rect 19628 32004 19684 34412
rect 19836 34300 20100 34310
rect 19892 34244 19940 34300
rect 19996 34244 20044 34300
rect 19836 34234 20100 34244
rect 20524 33684 20580 33694
rect 20412 33012 20468 33022
rect 20412 32918 20468 32956
rect 19740 32562 19796 32574
rect 19740 32510 19742 32562
rect 19794 32510 19796 32562
rect 19740 32452 19796 32510
rect 19740 32396 20244 32452
rect 19836 32284 20100 32294
rect 19892 32228 19940 32284
rect 19996 32228 20044 32284
rect 19836 32218 20100 32228
rect 19740 32004 19796 32014
rect 19628 32002 19796 32004
rect 19628 31950 19742 32002
rect 19794 31950 19796 32002
rect 19628 31948 19796 31950
rect 19740 31938 19796 31948
rect 20188 31892 20244 32396
rect 20188 31826 20244 31836
rect 20412 31780 20468 31790
rect 20524 31780 20580 33628
rect 20412 31778 20580 31780
rect 20412 31726 20414 31778
rect 20466 31726 20580 31778
rect 20412 31724 20580 31726
rect 20188 31332 20244 31342
rect 20412 31332 20468 31724
rect 20244 31276 20468 31332
rect 20188 31266 20244 31276
rect 19404 30772 19460 30782
rect 19292 30770 19460 30772
rect 19292 30718 19406 30770
rect 19458 30718 19460 30770
rect 19292 30716 19460 30718
rect 19404 30706 19460 30716
rect 19180 29810 19236 29820
rect 19628 30658 19684 30670
rect 19628 30606 19630 30658
rect 19682 30606 19684 30658
rect 19628 29876 19684 30606
rect 19836 30268 20100 30278
rect 19892 30212 19940 30268
rect 19996 30212 20044 30268
rect 19836 30202 20100 30212
rect 14924 29762 15092 29764
rect 14924 29710 14926 29762
rect 14978 29710 15092 29762
rect 14924 29708 15092 29710
rect 14924 29698 14980 29708
rect 15036 28868 15092 29708
rect 15148 28868 15204 28878
rect 15036 28866 15204 28868
rect 15036 28814 15150 28866
rect 15202 28814 15204 28866
rect 15036 28812 15204 28814
rect 15148 28802 15204 28812
rect 19628 28868 19684 29820
rect 19628 28802 19684 28812
rect 19516 28756 19572 28766
rect 14700 28578 14756 28588
rect 15036 28644 15092 28654
rect 15036 28550 15092 28588
rect 17836 28644 17892 28654
rect 12796 27918 12798 27970
rect 12850 27918 12852 27970
rect 12796 27906 12852 27918
rect 10220 27748 10276 27758
rect 10108 27746 10276 27748
rect 10108 27694 10222 27746
rect 10274 27694 10276 27746
rect 10108 27692 10276 27694
rect 9660 27682 9716 27692
rect 10220 27682 10276 27692
rect 17388 27746 17444 27758
rect 17388 27694 17390 27746
rect 17442 27694 17444 27746
rect 5740 26798 5742 26850
rect 5794 26798 5796 26850
rect 5740 26786 5796 26798
rect 15932 26740 15988 26750
rect 15932 26646 15988 26684
rect 16380 26626 16436 26638
rect 16380 26574 16382 26626
rect 16434 26574 16436 26626
rect 14588 25844 14644 25854
rect 13468 25730 13524 25742
rect 13468 25678 13470 25730
rect 13522 25678 13524 25730
rect 4476 25228 4740 25238
rect 4532 25172 4580 25228
rect 4636 25172 4684 25228
rect 4476 25162 4740 25172
rect 13468 24722 13524 25678
rect 13468 24670 13470 24722
rect 13522 24670 13524 24722
rect 11676 23716 11732 23726
rect 11676 23622 11732 23660
rect 13468 23716 13524 24670
rect 14588 23826 14644 25788
rect 14588 23774 14590 23826
rect 14642 23774 14644 23826
rect 14588 23762 14644 23774
rect 13468 23650 13524 23660
rect 15148 23716 15204 23726
rect 4476 23212 4740 23222
rect 4532 23156 4580 23212
rect 4636 23156 4684 23212
rect 4476 23146 4740 23156
rect 15148 22706 15204 23660
rect 16380 23044 16436 26574
rect 16940 26626 16996 26638
rect 16940 26574 16942 26626
rect 16994 26574 16996 26626
rect 16716 25956 16772 25966
rect 16716 25862 16772 25900
rect 16940 24834 16996 26574
rect 17052 26628 17108 26638
rect 17388 26628 17444 27694
rect 17724 27636 17780 27646
rect 17836 27636 17892 28588
rect 17724 27634 17892 27636
rect 17724 27582 17726 27634
rect 17778 27582 17892 27634
rect 17724 27580 17892 27582
rect 17724 27570 17780 27580
rect 17724 26628 17780 26638
rect 17388 26626 17780 26628
rect 17388 26574 17726 26626
rect 17778 26574 17780 26626
rect 17388 26572 17780 26574
rect 17052 26534 17108 26572
rect 17724 26068 17780 26572
rect 17836 26626 17892 27580
rect 19516 27746 19572 28700
rect 20300 28756 20356 28766
rect 20300 28662 20356 28700
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19516 27694 19518 27746
rect 19570 27694 19572 27746
rect 17836 26574 17838 26626
rect 17890 26574 17892 26626
rect 17836 26562 17892 26574
rect 17948 26628 18004 26638
rect 19516 26628 19572 27694
rect 19852 26628 19908 26638
rect 19516 26626 19908 26628
rect 19516 26574 19854 26626
rect 19906 26574 19908 26626
rect 19516 26572 19908 26574
rect 17724 26002 17780 26012
rect 17612 25844 17668 25854
rect 17612 25750 17668 25788
rect 17948 25730 18004 26572
rect 18956 26404 19012 26414
rect 18172 25956 18228 25966
rect 18172 25842 18228 25900
rect 18172 25790 18174 25842
rect 18226 25790 18228 25842
rect 18172 25778 18228 25790
rect 17948 25678 17950 25730
rect 18002 25678 18004 25730
rect 17948 25666 18004 25678
rect 18956 25618 19012 26348
rect 19852 26404 19908 26572
rect 19852 26338 19908 26348
rect 19836 26236 20100 26246
rect 19892 26180 19940 26236
rect 19996 26180 20044 26236
rect 19836 26170 20100 26180
rect 20524 25956 20580 25966
rect 20636 25956 20692 37772
rect 20748 36932 20804 38668
rect 21308 38658 21364 38668
rect 21532 38612 21588 38622
rect 21308 37940 21364 37950
rect 21084 37826 21140 37838
rect 21084 37774 21086 37826
rect 21138 37774 21140 37826
rect 21084 37716 21140 37774
rect 21308 37826 21364 37884
rect 21308 37774 21310 37826
rect 21362 37774 21364 37826
rect 21308 37762 21364 37774
rect 21532 37938 21588 38556
rect 21532 37886 21534 37938
rect 21586 37886 21588 37938
rect 21084 37650 21140 37660
rect 21196 37492 21252 37502
rect 21196 37490 21476 37492
rect 21196 37438 21198 37490
rect 21250 37438 21476 37490
rect 21196 37436 21476 37438
rect 21196 37426 21252 37436
rect 21420 36932 21476 37436
rect 21532 37156 21588 37886
rect 21756 37938 21812 37950
rect 21756 37886 21758 37938
rect 21810 37886 21812 37938
rect 21532 37100 21700 37156
rect 20748 36930 21364 36932
rect 20748 36878 20750 36930
rect 20802 36878 21364 36930
rect 20748 36876 21364 36878
rect 20748 35924 20804 36876
rect 21308 36818 21364 36876
rect 21420 36866 21476 36876
rect 21308 36766 21310 36818
rect 21362 36766 21364 36818
rect 21308 36754 21364 36766
rect 21644 36820 21700 37100
rect 21756 37044 21812 37886
rect 21756 36978 21812 36988
rect 21644 36764 21812 36820
rect 21420 36708 21476 36718
rect 21308 36036 21364 36046
rect 21420 36036 21476 36652
rect 21644 36596 21700 36606
rect 21644 36502 21700 36540
rect 21308 36034 21476 36036
rect 21308 35982 21310 36034
rect 21362 35982 21476 36034
rect 21308 35980 21476 35982
rect 21756 36036 21812 36764
rect 21308 35970 21364 35980
rect 21756 35942 21812 35980
rect 20748 35858 20804 35868
rect 21868 34020 21924 38780
rect 22092 38668 22148 42140
rect 22316 41074 22372 41086
rect 22316 41022 22318 41074
rect 22370 41022 22372 41074
rect 22316 40626 22372 41022
rect 22540 40740 22596 42476
rect 23548 40964 23604 42700
rect 23772 41972 23828 42814
rect 26348 42642 26404 42654
rect 26348 42590 26350 42642
rect 26402 42590 26404 42642
rect 26124 41972 26180 41982
rect 23772 41906 23828 41916
rect 26012 41916 26124 41972
rect 26012 41636 26068 41916
rect 26124 41878 26180 41916
rect 26348 41972 26404 42590
rect 26348 41906 26404 41916
rect 26460 41970 26516 43652
rect 27356 43652 27748 43708
rect 27356 42644 27412 43652
rect 27804 42868 27860 44494
rect 28140 43988 28196 44828
rect 28140 43874 28196 43932
rect 28140 43822 28142 43874
rect 28194 43822 28196 43874
rect 28140 43810 28196 43822
rect 28252 43708 28308 59276
rect 29568 59200 29680 60000
rect 28700 47794 28756 47806
rect 28700 47742 28702 47794
rect 28754 47742 28756 47794
rect 28588 46004 28644 46014
rect 28588 44994 28644 45948
rect 28588 44942 28590 44994
rect 28642 44942 28644 44994
rect 28588 43988 28644 44942
rect 28588 43922 28644 43932
rect 27804 42802 27860 42812
rect 28140 43652 28308 43708
rect 28700 43708 28756 47742
rect 29260 46674 29316 46686
rect 29260 46622 29262 46674
rect 29314 46622 29316 46674
rect 29260 46562 29316 46622
rect 29260 46510 29262 46562
rect 29314 46510 29316 46562
rect 29260 45780 29316 46510
rect 29260 45714 29316 45724
rect 29484 44884 29540 44894
rect 29484 44790 29540 44828
rect 28812 43988 28868 43998
rect 28812 43894 28868 43932
rect 28700 43652 29316 43708
rect 27804 42644 27860 42654
rect 27356 42642 27860 42644
rect 27356 42590 27358 42642
rect 27410 42590 27806 42642
rect 27858 42590 27860 42642
rect 27356 42588 27860 42590
rect 26460 41918 26462 41970
rect 26514 41918 26516 41970
rect 26460 41906 26516 41918
rect 26908 42084 26964 42094
rect 26796 41858 26852 41870
rect 26796 41806 26798 41858
rect 26850 41806 26852 41858
rect 26796 41748 26852 41806
rect 26796 41682 26852 41692
rect 23548 40962 24276 40964
rect 23548 40910 23550 40962
rect 23602 40910 24276 40962
rect 23548 40908 24276 40910
rect 23548 40898 23604 40908
rect 24220 40852 24276 40908
rect 26012 40852 26068 41580
rect 24220 40850 24724 40852
rect 24220 40798 24222 40850
rect 24274 40798 24724 40850
rect 24220 40796 24724 40798
rect 24220 40786 24276 40796
rect 22540 40674 22596 40684
rect 23100 40740 23156 40750
rect 22316 40574 22318 40626
rect 22370 40574 22372 40626
rect 22316 38836 22372 40574
rect 23100 40626 23156 40684
rect 23884 40740 23940 40750
rect 23940 40684 24164 40740
rect 23884 40646 23940 40684
rect 23100 40574 23102 40626
rect 23154 40574 23156 40626
rect 22428 40514 22484 40526
rect 22428 40462 22430 40514
rect 22482 40462 22484 40514
rect 22428 39954 22484 40462
rect 22428 39902 22430 39954
rect 22482 39902 22484 39954
rect 22428 39890 22484 39902
rect 22876 39954 22932 39966
rect 22876 39902 22878 39954
rect 22930 39902 22932 39954
rect 22652 39844 22708 39854
rect 22652 39750 22708 39788
rect 22652 38836 22708 38846
rect 22316 38834 22708 38836
rect 22316 38782 22654 38834
rect 22706 38782 22708 38834
rect 22316 38780 22708 38782
rect 22652 38770 22708 38780
rect 22876 38668 22932 39902
rect 22092 38612 22260 38668
rect 22204 38610 22260 38612
rect 22204 38558 22206 38610
rect 22258 38558 22260 38610
rect 22092 37940 22148 37950
rect 22092 37846 22148 37884
rect 22204 37716 22260 38558
rect 22204 37650 22260 37660
rect 22652 38612 22932 38668
rect 22988 38724 23044 38734
rect 23100 38724 23156 40574
rect 24108 40068 24164 40684
rect 24220 40068 24276 40078
rect 24108 40066 24276 40068
rect 24108 40014 24222 40066
rect 24274 40014 24276 40066
rect 24108 40012 24276 40014
rect 24220 39956 24276 40012
rect 24668 40068 24724 40796
rect 25564 40850 26068 40852
rect 25564 40798 26014 40850
rect 26066 40798 26068 40850
rect 25564 40796 26068 40798
rect 24668 39974 24724 40012
rect 25116 40628 25172 40638
rect 24220 39890 24276 39900
rect 25116 39956 25172 40572
rect 25116 39862 25172 39900
rect 25452 40068 25508 40078
rect 25452 39954 25508 40012
rect 25452 39902 25454 39954
rect 25506 39902 25508 39954
rect 25452 39890 25508 39902
rect 25452 39060 25508 39070
rect 25564 39060 25620 40796
rect 26012 40786 26068 40796
rect 26572 40404 26628 40414
rect 23044 38668 23156 38724
rect 24780 39058 25620 39060
rect 24780 39006 25454 39058
rect 25506 39006 25620 39058
rect 24780 39004 25620 39006
rect 26460 39844 26516 39854
rect 22988 38658 23044 38668
rect 23436 38612 23492 38622
rect 22652 37826 22708 38612
rect 22652 37774 22654 37826
rect 22706 37774 22708 37826
rect 22652 37716 22708 37774
rect 22652 37650 22708 37660
rect 23100 38610 23492 38612
rect 23100 38558 23438 38610
rect 23490 38558 23492 38610
rect 23100 38556 23492 38558
rect 22204 37492 22260 37502
rect 22204 37490 22372 37492
rect 22204 37438 22206 37490
rect 22258 37438 22372 37490
rect 22204 37436 22372 37438
rect 22204 37426 22260 37436
rect 21980 36932 22036 36942
rect 21980 36708 22036 36876
rect 21980 36614 22036 36652
rect 22204 36708 22260 36718
rect 22316 36708 22372 37436
rect 22540 37490 22596 37502
rect 22540 37438 22542 37490
rect 22594 37438 22596 37490
rect 22428 36708 22484 36718
rect 22316 36706 22484 36708
rect 22316 36654 22430 36706
rect 22482 36654 22484 36706
rect 22316 36652 22484 36654
rect 22204 36614 22260 36652
rect 21980 36036 22036 36046
rect 21980 35942 22036 35980
rect 22092 35476 22148 35486
rect 22316 35476 22372 35486
rect 22092 35474 22372 35476
rect 22092 35422 22094 35474
rect 22146 35422 22318 35474
rect 22370 35422 22372 35474
rect 22092 35420 22372 35422
rect 22092 35410 22148 35420
rect 22316 35410 22372 35420
rect 22428 34692 22484 36652
rect 22540 36708 22596 37438
rect 23100 37154 23156 38556
rect 23436 38546 23492 38556
rect 23548 37940 23604 37950
rect 23548 37846 23604 37884
rect 23100 37102 23102 37154
rect 23154 37102 23156 37154
rect 23100 37090 23156 37102
rect 23212 37714 23268 37726
rect 23212 37662 23214 37714
rect 23266 37662 23268 37714
rect 22540 36642 22596 36652
rect 22652 36706 22708 36718
rect 22652 36654 22654 36706
rect 22706 36654 22708 36706
rect 22540 35700 22596 35710
rect 22540 35028 22596 35644
rect 22652 35474 22708 36654
rect 22764 36484 22820 36494
rect 22764 36482 22932 36484
rect 22764 36430 22766 36482
rect 22818 36430 22932 36482
rect 22764 36428 22932 36430
rect 22764 36418 22820 36428
rect 22876 36148 22932 36428
rect 22876 35922 22932 36092
rect 23212 36036 23268 37662
rect 24780 36932 24836 39004
rect 25452 38994 25508 39004
rect 25116 38836 25172 38846
rect 25116 37828 25172 38780
rect 26124 38500 26180 38510
rect 25452 38498 26180 38500
rect 25452 38446 26126 38498
rect 26178 38446 26180 38498
rect 25452 38444 26180 38446
rect 25452 38050 25508 38444
rect 26124 38434 26180 38444
rect 25452 37998 25454 38050
rect 25506 37998 25508 38050
rect 25452 37986 25508 37998
rect 26012 38276 26068 38286
rect 25004 37826 25172 37828
rect 25004 37774 25118 37826
rect 25170 37774 25172 37826
rect 25004 37772 25172 37774
rect 23548 36930 24836 36932
rect 23548 36878 24782 36930
rect 24834 36878 24836 36930
rect 23548 36876 24836 36878
rect 23548 36818 23604 36876
rect 24780 36866 24836 36876
rect 24892 37716 24948 37726
rect 23548 36766 23550 36818
rect 23602 36766 23604 36818
rect 23548 36754 23604 36766
rect 23996 36706 24052 36718
rect 23996 36654 23998 36706
rect 24050 36654 24052 36706
rect 22876 35870 22878 35922
rect 22930 35870 22932 35922
rect 22876 35858 22932 35870
rect 23100 35980 23268 36036
rect 23548 36596 23604 36606
rect 23100 35700 23156 35980
rect 23100 35634 23156 35644
rect 23212 35812 23268 35822
rect 23212 35700 23268 35756
rect 23212 35698 23380 35700
rect 23212 35646 23214 35698
rect 23266 35646 23380 35698
rect 23212 35644 23380 35646
rect 23212 35634 23268 35644
rect 22652 35422 22654 35474
rect 22706 35422 22708 35474
rect 22652 35410 22708 35422
rect 22876 35474 22932 35486
rect 22876 35422 22878 35474
rect 22930 35422 22932 35474
rect 22876 35364 22932 35422
rect 22876 35308 23044 35364
rect 22540 34962 22596 34972
rect 22876 34916 22932 34926
rect 22652 34914 22932 34916
rect 22652 34862 22878 34914
rect 22930 34862 22932 34914
rect 22652 34860 22932 34862
rect 22540 34804 22596 34814
rect 22540 34710 22596 34748
rect 22428 34626 22484 34636
rect 21868 33964 22148 34020
rect 21980 33794 22036 33806
rect 21980 33742 21982 33794
rect 22034 33742 22036 33794
rect 21532 33684 21588 33694
rect 21532 33590 21588 33628
rect 21980 33684 22036 33742
rect 21980 33618 22036 33628
rect 21084 33012 21140 33022
rect 20748 32674 20804 32686
rect 20748 32622 20750 32674
rect 20802 32622 20804 32674
rect 20748 31556 20804 32622
rect 20972 31892 21028 31902
rect 20972 31798 21028 31836
rect 21084 31890 21140 32956
rect 21084 31838 21086 31890
rect 21138 31838 21140 31890
rect 21084 31826 21140 31838
rect 21868 31892 21924 31902
rect 21868 31798 21924 31836
rect 20748 31490 20804 31500
rect 20860 31780 20916 31790
rect 20860 31444 20916 31724
rect 21308 31784 21364 31796
rect 21308 31732 21310 31784
rect 21362 31780 21364 31784
rect 21420 31780 21476 31790
rect 21362 31732 21420 31780
rect 21308 31724 21420 31732
rect 21308 31720 21364 31724
rect 21420 31714 21476 31724
rect 21756 31778 21812 31790
rect 21756 31726 21758 31778
rect 21810 31726 21812 31778
rect 21756 31556 21812 31726
rect 21756 31490 21812 31500
rect 20860 31378 20916 31388
rect 21308 28756 21364 28766
rect 21308 28662 21364 28700
rect 20748 28644 20804 28654
rect 20748 28550 20804 28588
rect 21756 28644 21812 28654
rect 21812 28588 21924 28644
rect 21756 28578 21812 28588
rect 21644 28530 21700 28542
rect 21644 28478 21646 28530
rect 21698 28478 21700 28530
rect 21644 27858 21700 28478
rect 21644 27806 21646 27858
rect 21698 27806 21700 27858
rect 21644 27794 21700 27806
rect 20860 27748 20916 27758
rect 20860 27654 20916 27692
rect 21756 27746 21812 27758
rect 21756 27694 21758 27746
rect 21810 27694 21812 27746
rect 21644 27412 21700 27422
rect 21644 26626 21700 27356
rect 21756 26740 21812 27694
rect 21868 26908 21924 28588
rect 21868 26852 22036 26908
rect 21868 26740 21924 26750
rect 21756 26738 21924 26740
rect 21756 26686 21870 26738
rect 21922 26686 21924 26738
rect 21756 26684 21924 26686
rect 21644 26574 21646 26626
rect 21698 26574 21700 26626
rect 21644 26562 21700 26574
rect 21868 26628 21924 26684
rect 20748 26516 20804 26526
rect 20748 26422 20804 26460
rect 18956 25566 18958 25618
rect 19010 25566 19012 25618
rect 18620 25396 18676 25406
rect 18620 25302 18676 25340
rect 16940 24782 16942 24834
rect 16994 24782 16996 24834
rect 16940 24770 16996 24782
rect 18956 24836 19012 25566
rect 20300 25954 20692 25956
rect 20300 25902 20526 25954
rect 20578 25902 20692 25954
rect 20300 25900 20692 25902
rect 20972 26404 21028 26414
rect 19180 24836 19236 24846
rect 18956 24834 19236 24836
rect 18956 24782 19182 24834
rect 19234 24782 19236 24834
rect 18956 24780 19236 24782
rect 17500 23716 17556 23726
rect 16604 23044 16660 23054
rect 16380 23042 16660 23044
rect 16380 22990 16606 23042
rect 16658 22990 16660 23042
rect 16380 22988 16660 22990
rect 16604 22978 16660 22988
rect 17500 22820 17556 23660
rect 18844 23716 18900 23726
rect 18956 23716 19012 24780
rect 19180 24770 19236 24780
rect 19404 24836 19460 24846
rect 19180 23828 19236 23838
rect 19236 23772 19348 23828
rect 19180 23734 19236 23772
rect 18900 23660 19012 23716
rect 18844 23622 18900 23660
rect 17612 22820 17668 22830
rect 17500 22818 17668 22820
rect 17500 22766 17614 22818
rect 17666 22766 17668 22818
rect 17500 22764 17668 22766
rect 19292 22820 19348 23772
rect 19404 23826 19460 24780
rect 20300 24834 20356 25900
rect 20524 25890 20580 25900
rect 20300 24782 20302 24834
rect 20354 24782 20356 24834
rect 20188 24612 20244 24622
rect 19852 24498 19908 24510
rect 19852 24446 19854 24498
rect 19906 24446 19908 24498
rect 19852 24386 19908 24446
rect 19852 24334 19854 24386
rect 19906 24334 19908 24386
rect 19852 24322 19908 24334
rect 19836 24220 20100 24230
rect 19892 24164 19940 24220
rect 19996 24164 20044 24220
rect 19836 24154 20100 24164
rect 19404 23774 19406 23826
rect 19458 23774 19460 23826
rect 19404 23762 19460 23774
rect 19404 22820 19460 22830
rect 19852 22820 19908 22830
rect 19292 22818 19908 22820
rect 19292 22766 19406 22818
rect 19458 22766 19854 22818
rect 19906 22766 19908 22818
rect 19292 22764 19908 22766
rect 20188 22820 20244 24556
rect 20300 24388 20356 24782
rect 20972 25618 21028 26348
rect 20972 25566 20974 25618
rect 21026 25566 21028 25618
rect 20972 24724 21028 25566
rect 21420 26068 21476 26078
rect 21420 25732 21476 26012
rect 21868 26068 21924 26572
rect 21868 26002 21924 26012
rect 21420 25618 21476 25676
rect 21420 25566 21422 25618
rect 21474 25566 21476 25618
rect 21420 25554 21476 25566
rect 21868 25844 21924 25854
rect 21980 25844 22036 26852
rect 22092 26852 22148 33964
rect 22652 34018 22708 34860
rect 22876 34850 22932 34860
rect 22876 34692 22932 34702
rect 22988 34692 23044 35308
rect 23324 34802 23380 35644
rect 23324 34750 23326 34802
rect 23378 34750 23380 34802
rect 23324 34738 23380 34750
rect 23548 34804 23604 36540
rect 23772 35924 23828 35934
rect 23996 35924 24052 36654
rect 24220 36706 24276 36718
rect 24220 36654 24222 36706
rect 24274 36654 24276 36706
rect 24220 36596 24276 36654
rect 24220 36530 24276 36540
rect 24892 36484 24948 37660
rect 23772 35922 24052 35924
rect 23772 35870 23774 35922
rect 23826 35870 24052 35922
rect 23772 35868 24052 35870
rect 24332 36428 24948 36484
rect 23772 35700 23828 35868
rect 24108 35812 24164 35822
rect 24108 35718 24164 35756
rect 24332 35810 24388 36428
rect 24780 36036 24836 36046
rect 24780 35942 24836 35980
rect 24332 35758 24334 35810
rect 24386 35758 24388 35810
rect 23772 35634 23828 35644
rect 23548 34710 23604 34748
rect 22876 34690 23044 34692
rect 22876 34638 22878 34690
rect 22930 34638 23044 34690
rect 22876 34636 23044 34638
rect 23772 34692 23828 34702
rect 22876 34626 22932 34636
rect 23772 34598 23828 34636
rect 22652 33966 22654 34018
rect 22706 33966 22708 34018
rect 22652 33954 22708 33966
rect 23100 34578 23156 34590
rect 23100 34526 23102 34578
rect 23154 34526 23156 34578
rect 22428 33684 22484 33694
rect 22428 32898 22484 33628
rect 22428 32846 22430 32898
rect 22482 32846 22484 32898
rect 22428 32834 22484 32846
rect 22764 33684 22820 33694
rect 22764 32562 22820 33628
rect 22764 32510 22766 32562
rect 22818 32510 22820 32562
rect 22540 31892 22596 31902
rect 22764 31892 22820 32510
rect 22876 32564 22932 32574
rect 23100 32564 23156 34526
rect 23212 34580 23268 34590
rect 23212 33796 23268 34524
rect 23212 32786 23268 33740
rect 23212 32734 23214 32786
rect 23266 32734 23268 32786
rect 23212 32722 23268 32734
rect 23996 34578 24052 34590
rect 23996 34526 23998 34578
rect 24050 34526 24052 34578
rect 23996 32674 24052 34526
rect 23996 32622 23998 32674
rect 24050 32622 24052 32674
rect 23996 32610 24052 32622
rect 24220 34578 24276 34590
rect 24220 34526 24222 34578
rect 24274 34526 24276 34578
rect 22876 32562 23156 32564
rect 22876 32510 22878 32562
rect 22930 32510 23156 32562
rect 22876 32508 23156 32510
rect 22876 32498 22932 32508
rect 22540 31890 22820 31892
rect 22540 31838 22542 31890
rect 22594 31838 22820 31890
rect 22540 31836 22820 31838
rect 22876 32002 22932 32014
rect 22876 31950 22878 32002
rect 22930 31950 22932 32002
rect 22540 31826 22596 31836
rect 22764 31668 22820 31678
rect 22764 30658 22820 31612
rect 22876 31556 22932 31950
rect 22876 31490 22932 31500
rect 22988 30772 23044 32508
rect 23884 32340 23940 32350
rect 23660 32002 23716 32014
rect 23660 31950 23662 32002
rect 23714 31950 23716 32002
rect 23212 31780 23268 31790
rect 23212 31686 23268 31724
rect 23660 31666 23716 31950
rect 23884 31890 23940 32284
rect 24220 32004 24276 34526
rect 24332 33460 24388 35758
rect 24444 35812 24500 35822
rect 24444 34802 24500 35756
rect 24444 34750 24446 34802
rect 24498 34750 24500 34802
rect 24444 34738 24500 34750
rect 24668 33684 24724 33694
rect 24668 33590 24724 33628
rect 24332 33404 24724 33460
rect 24220 31938 24276 31948
rect 23884 31838 23886 31890
rect 23938 31838 23940 31890
rect 23884 31826 23940 31838
rect 24108 31892 24164 31902
rect 24108 31798 24164 31836
rect 23660 31614 23662 31666
rect 23714 31614 23716 31666
rect 23660 31602 23716 31614
rect 24332 31778 24388 31790
rect 24332 31726 24334 31778
rect 24386 31726 24388 31778
rect 24108 31556 24164 31566
rect 23772 31444 23828 31454
rect 24108 31444 24164 31500
rect 24332 31444 24388 31726
rect 23828 31388 23940 31444
rect 23772 31378 23828 31388
rect 23884 31106 23940 31388
rect 23884 31054 23886 31106
rect 23938 31054 23940 31106
rect 23884 31042 23940 31054
rect 24108 31388 24388 31444
rect 24556 31666 24612 31678
rect 24556 31614 24558 31666
rect 24610 31614 24612 31666
rect 23548 30772 23604 30782
rect 22988 30770 23604 30772
rect 22988 30718 23550 30770
rect 23602 30718 23604 30770
rect 22988 30716 23604 30718
rect 23548 30706 23604 30716
rect 23772 30770 23828 30782
rect 23772 30718 23774 30770
rect 23826 30718 23828 30770
rect 22764 30606 22766 30658
rect 22818 30606 22820 30658
rect 22764 30594 22820 30606
rect 22652 30548 22708 30558
rect 22316 28756 22372 28766
rect 22316 28662 22372 28700
rect 22652 28082 22708 30492
rect 23100 30546 23156 30558
rect 23100 30494 23102 30546
rect 23154 30494 23156 30546
rect 23100 29988 23156 30494
rect 23100 29922 23156 29932
rect 22988 28756 23044 28766
rect 22652 28030 22654 28082
rect 22706 28030 22708 28082
rect 22652 28018 22708 28030
rect 22764 28530 22820 28542
rect 22764 28478 22766 28530
rect 22818 28478 22820 28530
rect 22204 27748 22260 27758
rect 22204 27654 22260 27692
rect 22540 26852 22596 26862
rect 22092 26796 22260 26852
rect 22092 26626 22148 26638
rect 22092 26574 22094 26626
rect 22146 26574 22148 26626
rect 22092 26516 22148 26574
rect 22092 26450 22148 26460
rect 21868 25842 22036 25844
rect 21868 25790 21870 25842
rect 21922 25790 22036 25842
rect 21868 25788 22036 25790
rect 21868 24948 21924 25788
rect 21644 24892 21924 24948
rect 21644 24836 21700 24892
rect 21644 24742 21700 24780
rect 22092 24836 22148 24846
rect 22092 24742 22148 24780
rect 21084 24724 21140 24734
rect 20972 24668 21084 24724
rect 20300 24322 20356 24332
rect 20748 24498 20804 24510
rect 20748 24446 20750 24498
rect 20802 24446 20804 24498
rect 20748 24386 20804 24446
rect 20748 24334 20750 24386
rect 20802 24334 20804 24386
rect 20748 23940 20804 24334
rect 20748 23874 20804 23884
rect 21084 23938 21140 24668
rect 22204 24724 22260 26796
rect 22540 26758 22596 26796
rect 22764 26516 22820 28478
rect 22988 27972 23044 28700
rect 23436 27972 23492 27982
rect 22988 27970 23492 27972
rect 22988 27918 22990 27970
rect 23042 27918 23438 27970
rect 23490 27918 23492 27970
rect 22988 27916 23492 27918
rect 22988 27906 23044 27916
rect 23436 27906 23492 27916
rect 23660 27748 23716 27758
rect 23548 27692 23660 27748
rect 22876 27412 22932 27422
rect 22876 27318 22932 27356
rect 23548 26852 23604 27692
rect 23660 27682 23716 27692
rect 23772 27524 23828 30718
rect 23996 30772 24052 30782
rect 23996 30678 24052 30716
rect 24108 30548 24164 31388
rect 23884 30492 24164 30548
rect 24220 30770 24276 30782
rect 24220 30718 24222 30770
rect 24274 30718 24276 30770
rect 23884 29874 23940 30492
rect 24220 30324 24276 30718
rect 23884 29822 23886 29874
rect 23938 29822 23940 29874
rect 23884 29540 23940 29822
rect 23996 30268 24276 30324
rect 24556 30770 24612 31614
rect 24556 30718 24558 30770
rect 24610 30718 24612 30770
rect 23996 29652 24052 30268
rect 24444 30098 24500 30110
rect 24444 30046 24446 30098
rect 24498 30046 24500 30098
rect 24332 29988 24388 29998
rect 24220 29874 24276 29886
rect 24220 29822 24222 29874
rect 24274 29822 24276 29874
rect 23996 29596 24164 29652
rect 23884 29474 23940 29484
rect 23996 27746 24052 27758
rect 23996 27694 23998 27746
rect 24050 27694 24052 27746
rect 23884 27524 23940 27534
rect 23772 27522 23940 27524
rect 23772 27470 23886 27522
rect 23938 27470 23940 27522
rect 23772 27468 23940 27470
rect 23884 27458 23940 27468
rect 23884 26964 23940 26974
rect 23996 26964 24052 27694
rect 23884 26962 24052 26964
rect 23884 26910 23886 26962
rect 23938 26910 24052 26962
rect 23884 26908 24052 26910
rect 23884 26898 23940 26908
rect 24108 26852 24164 29596
rect 24220 29204 24276 29822
rect 24332 29764 24388 29932
rect 24444 29876 24500 30046
rect 24556 29988 24612 30718
rect 24556 29922 24612 29932
rect 24668 29876 24724 33404
rect 24780 32340 24836 32350
rect 24780 30770 24836 32284
rect 25004 31556 25060 37772
rect 25116 37762 25172 37772
rect 25788 37940 25844 37950
rect 25564 37716 25620 37726
rect 25452 37714 25620 37716
rect 25452 37662 25566 37714
rect 25618 37662 25620 37714
rect 25452 37660 25620 37662
rect 25340 36708 25396 36718
rect 25116 36596 25172 36606
rect 25116 35810 25172 36540
rect 25340 36034 25396 36652
rect 25340 35982 25342 36034
rect 25394 35982 25396 36034
rect 25340 35970 25396 35982
rect 25116 35758 25118 35810
rect 25170 35758 25172 35810
rect 25116 35746 25172 35758
rect 25228 33906 25284 33918
rect 25228 33854 25230 33906
rect 25282 33854 25284 33906
rect 25228 33684 25284 33854
rect 25228 33618 25284 33628
rect 25340 32004 25396 32014
rect 25340 31890 25396 31948
rect 25340 31838 25342 31890
rect 25394 31838 25396 31890
rect 25228 31778 25284 31790
rect 25228 31726 25230 31778
rect 25282 31726 25284 31778
rect 25228 31668 25284 31726
rect 25228 31602 25284 31612
rect 24780 30718 24782 30770
rect 24834 30718 24836 30770
rect 24780 30706 24836 30718
rect 24892 31500 25004 31556
rect 24444 29810 24500 29820
rect 24663 29820 24724 29876
rect 24780 29874 24836 29886
rect 24780 29822 24782 29874
rect 24834 29822 24836 29874
rect 24663 29764 24719 29820
rect 24332 29698 24388 29708
rect 24556 29708 24719 29764
rect 24220 29138 24276 29148
rect 24220 28980 24276 28990
rect 24556 28980 24612 29708
rect 24220 27746 24276 28924
rect 24220 27694 24222 27746
rect 24274 27694 24276 27746
rect 24220 27682 24276 27694
rect 24332 28924 24612 28980
rect 24332 26908 24388 28924
rect 24780 28866 24836 29822
rect 24780 28814 24782 28866
rect 24834 28814 24836 28866
rect 24780 28802 24836 28814
rect 24444 28756 24500 28766
rect 24444 28754 24724 28756
rect 24444 28702 24446 28754
rect 24498 28702 24724 28754
rect 24444 28700 24724 28702
rect 24444 28690 24500 28700
rect 24668 28644 24724 28700
rect 24892 28644 24948 31500
rect 25004 31490 25060 31500
rect 25116 31108 25172 31118
rect 25116 31014 25172 31052
rect 25004 30660 25060 30670
rect 25004 30566 25060 30604
rect 25228 29874 25284 29886
rect 25228 29822 25230 29874
rect 25282 29822 25284 29874
rect 25004 29764 25060 29774
rect 25004 28980 25060 29708
rect 25228 29540 25284 29822
rect 25228 29474 25284 29484
rect 25004 28914 25060 28924
rect 25228 28866 25284 28878
rect 25228 28814 25230 28866
rect 25282 28814 25284 28866
rect 25116 28756 25172 28766
rect 25116 28662 25172 28700
rect 24668 28588 24948 28644
rect 24556 28530 24612 28542
rect 24556 28478 24558 28530
rect 24610 28478 24612 28530
rect 24444 27748 24500 27758
rect 24444 27654 24500 27692
rect 24332 26852 24500 26908
rect 22428 26460 22820 26516
rect 22876 26796 23604 26852
rect 23996 26796 24164 26852
rect 22428 25732 22484 26460
rect 21756 24500 21812 24510
rect 21084 23886 21086 23938
rect 21138 23886 21140 23938
rect 21084 23874 21140 23886
rect 21532 23940 21588 23950
rect 20300 22820 20356 22830
rect 20748 22820 20804 22830
rect 20188 22818 20804 22820
rect 20188 22766 20302 22818
rect 20354 22766 20750 22818
rect 20802 22766 20804 22818
rect 20188 22764 20804 22766
rect 17612 22754 17668 22764
rect 19404 22754 19460 22764
rect 15148 22654 15150 22706
rect 15202 22654 15204 22706
rect 15148 22642 15204 22654
rect 19852 22372 19908 22764
rect 19852 22316 20244 22372
rect 19836 22204 20100 22214
rect 19892 22148 19940 22204
rect 19996 22148 20044 22204
rect 19836 22138 20100 22148
rect 19852 21700 19908 21710
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 18508 20692 18564 20702
rect 17724 19682 17780 19694
rect 17724 19630 17726 19682
rect 17778 19630 17780 19682
rect 4476 19180 4740 19190
rect 4532 19124 4580 19180
rect 4636 19124 4684 19180
rect 4476 19114 4740 19124
rect 17500 18676 17556 18686
rect 17500 18582 17556 18620
rect 16604 18564 16660 18574
rect 16604 18470 16660 18508
rect 17724 18564 17780 19630
rect 18396 19124 18452 19134
rect 18284 19068 18396 19124
rect 18284 18676 18340 19068
rect 18396 19058 18452 19068
rect 18284 18582 18340 18620
rect 17052 18450 17108 18462
rect 17052 18398 17054 18450
rect 17106 18398 17108 18450
rect 16828 17556 16884 17566
rect 17052 17556 17108 18398
rect 16884 17500 17108 17556
rect 17612 17668 17668 17678
rect 17724 17668 17780 18508
rect 18060 18562 18116 18574
rect 18060 18510 18062 18562
rect 18114 18510 18116 18562
rect 18060 18452 18116 18510
rect 18508 18564 18564 20636
rect 19292 20580 19348 20590
rect 19292 19458 19348 20524
rect 19740 20468 19796 20478
rect 19740 20374 19796 20412
rect 19852 20356 19908 21644
rect 19852 20290 19908 20300
rect 20188 21698 20244 22316
rect 20300 21924 20356 22764
rect 20748 22754 20804 22764
rect 20300 21858 20356 21868
rect 21532 21812 21588 23884
rect 21756 23938 21812 24444
rect 21756 23886 21758 23938
rect 21810 23886 21812 23938
rect 21756 23874 21812 23886
rect 21868 23828 21924 23838
rect 21868 23268 21924 23772
rect 21644 23212 21924 23268
rect 21644 22818 21700 23212
rect 21644 22766 21646 22818
rect 21698 22766 21700 22818
rect 21644 22754 21700 22766
rect 22092 22820 22148 22830
rect 22204 22820 22260 24668
rect 22316 25676 22428 25732
rect 22316 24612 22372 25676
rect 22428 25638 22484 25676
rect 22540 26292 22596 26302
rect 22428 24724 22484 24734
rect 22540 24724 22596 26236
rect 22764 26068 22820 26078
rect 22764 25974 22820 26012
rect 22876 24834 22932 26796
rect 23772 26738 23828 26750
rect 23772 26686 23774 26738
rect 23826 26686 23828 26738
rect 23548 26628 23604 26638
rect 23548 26534 23604 26572
rect 23324 26516 23380 26526
rect 23772 26516 23828 26686
rect 23324 26422 23380 26460
rect 23660 26460 23772 26516
rect 23212 26404 23268 26414
rect 22876 24782 22878 24834
rect 22930 24782 22932 24834
rect 22876 24770 22932 24782
rect 23100 25730 23156 25742
rect 23100 25678 23102 25730
rect 23154 25678 23156 25730
rect 22428 24722 22596 24724
rect 22428 24670 22430 24722
rect 22482 24670 22596 24722
rect 22428 24668 22596 24670
rect 22428 24658 22484 24668
rect 22316 23828 22372 24556
rect 22540 24500 22596 24510
rect 22316 23762 22372 23772
rect 22428 24498 22596 24500
rect 22428 24446 22542 24498
rect 22594 24446 22596 24498
rect 22428 24444 22596 24446
rect 22092 22818 22260 22820
rect 22092 22766 22094 22818
rect 22146 22766 22260 22818
rect 22092 22764 22260 22766
rect 22092 22754 22148 22764
rect 21532 21810 21700 21812
rect 21532 21758 21534 21810
rect 21586 21758 21700 21810
rect 21532 21756 21700 21758
rect 21532 21746 21588 21756
rect 20188 21646 20190 21698
rect 20242 21646 20244 21698
rect 19836 20188 20100 20198
rect 19892 20132 19940 20188
rect 19996 20132 20044 20188
rect 19836 20122 20100 20132
rect 19292 19406 19294 19458
rect 19346 19406 19348 19458
rect 19292 19394 19348 19406
rect 20188 19796 20244 21646
rect 20300 20692 20356 20702
rect 20300 20468 20356 20636
rect 21420 20578 21476 20590
rect 21420 20526 21422 20578
rect 21474 20526 21476 20578
rect 20748 20468 20804 20478
rect 20300 20466 20804 20468
rect 20300 20414 20302 20466
rect 20354 20414 20750 20466
rect 20802 20414 20804 20466
rect 20300 20412 20804 20414
rect 20300 20402 20356 20412
rect 20748 20244 20804 20412
rect 20748 20178 20804 20188
rect 20636 20132 20692 20142
rect 20636 19908 20692 20076
rect 20636 19906 21028 19908
rect 20636 19854 20638 19906
rect 20690 19854 21028 19906
rect 20636 19852 21028 19854
rect 20636 19842 20692 19852
rect 20188 19236 20244 19740
rect 20972 19682 21028 19852
rect 21084 19796 21140 19806
rect 21084 19702 21140 19740
rect 20972 19630 20974 19682
rect 21026 19630 21028 19682
rect 20972 19618 21028 19630
rect 20188 19180 20468 19236
rect 19516 19124 19572 19134
rect 18508 18498 18564 18508
rect 18956 18674 19012 18686
rect 18956 18622 18958 18674
rect 19010 18622 19012 18674
rect 18956 18564 19012 18622
rect 18956 18498 19012 18508
rect 18284 18452 18340 18462
rect 18060 18396 18284 18452
rect 17612 17666 17780 17668
rect 17612 17614 17614 17666
rect 17666 17614 17780 17666
rect 17612 17612 17780 17614
rect 18284 17666 18340 18396
rect 19180 18452 19236 18462
rect 19180 18358 19236 18396
rect 19516 18450 19572 19068
rect 20188 19124 20244 19180
rect 20188 19058 20244 19068
rect 20300 19012 20356 19022
rect 19740 18676 19796 18686
rect 19740 18582 19796 18620
rect 19516 18398 19518 18450
rect 19570 18398 19572 18450
rect 19516 18386 19572 18398
rect 20076 18450 20132 18462
rect 20076 18398 20078 18450
rect 20130 18398 20132 18450
rect 18732 18340 18788 18350
rect 20076 18340 20132 18398
rect 18732 18338 19124 18340
rect 18732 18286 18734 18338
rect 18786 18286 19124 18338
rect 18732 18284 19124 18286
rect 20076 18284 20244 18340
rect 18732 18274 18788 18284
rect 19068 18004 19124 18284
rect 19836 18172 20100 18182
rect 19892 18116 19940 18172
rect 19996 18116 20044 18172
rect 19836 18106 20100 18116
rect 20188 18004 20244 18284
rect 19068 17948 19796 18004
rect 19740 17778 19796 17948
rect 19740 17726 19742 17778
rect 19794 17726 19796 17778
rect 19740 17714 19796 17726
rect 19852 17948 20244 18004
rect 18284 17614 18286 17666
rect 18338 17614 18340 17666
rect 16828 17462 16884 17500
rect 4476 17164 4740 17174
rect 4532 17108 4580 17164
rect 4636 17108 4684 17164
rect 4476 17098 4740 17108
rect 15036 16660 15092 16670
rect 15036 16566 15092 16604
rect 17612 16660 17668 17612
rect 17612 16594 17668 16604
rect 18284 17556 18340 17614
rect 18172 15538 18228 15550
rect 18172 15486 18174 15538
rect 18226 15486 18228 15538
rect 18172 15426 18228 15486
rect 18172 15374 18174 15426
rect 18226 15374 18228 15426
rect 18172 15362 18228 15374
rect 4476 15148 4740 15158
rect 4532 15092 4580 15148
rect 4636 15092 4684 15148
rect 4476 15082 4740 15092
rect 17612 13524 17668 13534
rect 4476 13132 4740 13142
rect 4532 13076 4580 13132
rect 4636 13076 4684 13132
rect 4476 13066 4740 13076
rect 17612 12628 17668 13468
rect 17500 12626 17668 12628
rect 17500 12574 17614 12626
rect 17666 12574 17668 12626
rect 17500 12572 17668 12574
rect 17500 11618 17556 12572
rect 17612 12562 17668 12572
rect 18284 12514 18340 17500
rect 18732 17556 18788 17566
rect 18732 17462 18788 17500
rect 19852 16884 19908 17948
rect 20300 17892 20356 18956
rect 20412 18786 20468 19180
rect 21420 19012 21476 20526
rect 21532 20580 21588 20590
rect 21532 20486 21588 20524
rect 21420 18946 21476 18956
rect 20412 18734 20414 18786
rect 20466 18734 20468 18786
rect 20412 18722 20468 18734
rect 21420 18788 21476 18798
rect 21644 18788 21700 21756
rect 22092 20580 22148 20590
rect 22092 20486 22148 20524
rect 22204 19908 22260 22764
rect 22428 21028 22484 24444
rect 22540 24434 22596 24444
rect 22876 24500 22932 24510
rect 22876 24406 22932 24444
rect 22652 24388 22708 24398
rect 22540 23940 22596 23950
rect 22540 22818 22596 23884
rect 22652 23714 22708 24332
rect 23100 24052 23156 25678
rect 23212 24722 23268 26348
rect 23436 25844 23492 25854
rect 23436 25750 23492 25788
rect 23212 24670 23214 24722
rect 23266 24670 23268 24722
rect 23212 24658 23268 24670
rect 23324 24724 23380 24734
rect 23324 24630 23380 24668
rect 23548 24498 23604 24510
rect 23548 24446 23550 24498
rect 23602 24446 23604 24498
rect 23548 24388 23604 24446
rect 23548 24322 23604 24332
rect 23100 23996 23268 24052
rect 22652 23662 22654 23714
rect 22706 23662 22708 23714
rect 22652 23650 22708 23662
rect 23100 23828 23156 23838
rect 22540 22766 22542 22818
rect 22594 22766 22596 22818
rect 22540 22754 22596 22766
rect 22988 22482 23044 22494
rect 22988 22430 22990 22482
rect 23042 22430 23044 22482
rect 22652 21698 22708 21710
rect 22652 21646 22654 21698
rect 22706 21646 22708 21698
rect 22540 21028 22596 21038
rect 22428 21026 22596 21028
rect 22428 20974 22542 21026
rect 22594 20974 22596 21026
rect 22428 20972 22596 20974
rect 22652 21028 22708 21646
rect 22764 21028 22820 21038
rect 22652 21026 22820 21028
rect 22652 20974 22766 21026
rect 22818 20974 22820 21026
rect 22652 20972 22820 20974
rect 22540 20962 22596 20972
rect 22764 20962 22820 20972
rect 22876 20804 22932 20814
rect 22988 20804 23044 22430
rect 23100 21476 23156 23772
rect 23212 23604 23268 23996
rect 23548 23940 23604 23950
rect 23548 23714 23604 23884
rect 23548 23662 23550 23714
rect 23602 23662 23604 23714
rect 23548 23650 23604 23662
rect 23660 23716 23716 26460
rect 23772 26450 23828 26460
rect 23884 25732 23940 25742
rect 23660 23650 23716 23660
rect 23772 25730 23940 25732
rect 23772 25678 23886 25730
rect 23938 25678 23940 25730
rect 23772 25676 23940 25678
rect 23212 23538 23268 23548
rect 23772 21922 23828 25676
rect 23884 25666 23940 25676
rect 23884 24612 23940 24622
rect 23884 24518 23940 24556
rect 23996 24388 24052 26796
rect 24444 26738 24500 26852
rect 24556 26852 24612 28478
rect 24892 27972 24948 28588
rect 25004 28532 25060 28542
rect 25004 28438 25060 28476
rect 25228 28196 25284 28814
rect 25340 28644 25396 31838
rect 25452 31892 25508 37660
rect 25564 37650 25620 37660
rect 25564 35924 25620 35934
rect 25564 35830 25620 35868
rect 25788 35922 25844 37884
rect 26012 37826 26068 38220
rect 26460 37938 26516 39788
rect 26572 38834 26628 40348
rect 26572 38782 26574 38834
rect 26626 38782 26628 38834
rect 26572 38770 26628 38782
rect 26460 37886 26462 37938
rect 26514 37886 26516 37938
rect 26460 37874 26516 37886
rect 26012 37774 26014 37826
rect 26066 37774 26068 37826
rect 26012 37762 26068 37774
rect 26348 37716 26404 37726
rect 26348 37622 26404 37660
rect 25788 35870 25790 35922
rect 25842 35870 25844 35922
rect 25564 34020 25620 34030
rect 25564 34018 25732 34020
rect 25564 33966 25566 34018
rect 25618 33966 25732 34018
rect 25564 33964 25732 33966
rect 25564 33954 25620 33964
rect 25676 33124 25732 33964
rect 25788 33348 25844 35870
rect 25900 35812 25956 35822
rect 25900 35718 25956 35756
rect 26236 35810 26292 35822
rect 26236 35758 26238 35810
rect 26290 35758 26292 35810
rect 25900 34580 25956 34590
rect 26236 34580 26292 35758
rect 25956 34524 26292 34580
rect 25900 34486 25956 34524
rect 26796 34020 26852 34030
rect 26572 33964 26796 34020
rect 25788 33282 25844 33292
rect 26460 33908 26516 33918
rect 26460 33682 26516 33852
rect 26460 33630 26462 33682
rect 26514 33630 26516 33682
rect 25676 33068 26404 33124
rect 25564 31892 25620 31902
rect 25452 31890 25620 31892
rect 25452 31838 25566 31890
rect 25618 31838 25620 31890
rect 25452 31836 25620 31838
rect 25564 31826 25620 31836
rect 25676 31668 25732 33068
rect 26124 32900 26180 32910
rect 26012 32786 26068 32798
rect 26012 32734 26014 32786
rect 26066 32734 26068 32786
rect 25564 31612 25732 31668
rect 25900 31890 25956 31902
rect 25900 31838 25902 31890
rect 25954 31838 25956 31890
rect 25564 30660 25620 31612
rect 25788 31554 25844 31566
rect 25788 31502 25790 31554
rect 25842 31502 25844 31554
rect 25788 30884 25844 31502
rect 25788 30818 25844 30828
rect 25900 30772 25956 31838
rect 26012 31780 26068 32734
rect 26012 31714 26068 31724
rect 26124 30994 26180 32844
rect 26348 32674 26404 33068
rect 26348 32622 26350 32674
rect 26402 32622 26404 32674
rect 26124 30942 26126 30994
rect 26178 30942 26180 30994
rect 26124 30930 26180 30942
rect 26236 31890 26292 31902
rect 26236 31838 26238 31890
rect 26290 31838 26292 31890
rect 26236 30884 26292 31838
rect 26348 31890 26404 32622
rect 26348 31838 26350 31890
rect 26402 31838 26404 31890
rect 26348 31826 26404 31838
rect 26460 31892 26516 33630
rect 26460 31826 26516 31836
rect 26348 31556 26404 31566
rect 26404 31500 26516 31556
rect 26348 31490 26404 31500
rect 26236 30818 26292 30828
rect 25564 30566 25620 30604
rect 25676 30658 25732 30670
rect 25676 30606 25678 30658
rect 25730 30606 25732 30658
rect 25676 30212 25732 30606
rect 25900 30548 25956 30716
rect 26460 30770 26516 31500
rect 26460 30718 26462 30770
rect 26514 30718 26516 30770
rect 26460 30706 26516 30718
rect 26348 30660 26404 30670
rect 26348 30566 26404 30604
rect 26012 30548 26068 30558
rect 25900 30546 26068 30548
rect 25900 30494 26014 30546
rect 26066 30494 26068 30546
rect 25900 30492 26068 30494
rect 26012 30324 26068 30492
rect 26012 30258 26068 30268
rect 26460 30436 26516 30446
rect 25788 30212 25844 30222
rect 25676 30156 25788 30212
rect 25788 30146 25844 30156
rect 25564 30100 25620 30110
rect 25564 30006 25620 30044
rect 26460 30098 26516 30380
rect 26572 30324 26628 33964
rect 26796 33926 26852 33964
rect 26908 33908 26964 42028
rect 27132 41972 27188 41982
rect 27132 41878 27188 41916
rect 27020 41636 27076 41646
rect 27356 41636 27412 42588
rect 27804 42578 27860 42588
rect 28028 42644 28084 42654
rect 28028 42084 28084 42588
rect 28028 41970 28084 42028
rect 28028 41918 28030 41970
rect 28082 41918 28084 41970
rect 28028 41906 28084 41918
rect 27468 41860 27524 41870
rect 27468 41858 27748 41860
rect 27468 41806 27470 41858
rect 27522 41806 27748 41858
rect 27468 41804 27748 41806
rect 27468 41794 27524 41804
rect 27076 41580 27524 41636
rect 27020 41570 27076 41580
rect 27020 40514 27076 40526
rect 27020 40462 27022 40514
rect 27074 40462 27076 40514
rect 27020 40404 27076 40462
rect 27020 40338 27076 40348
rect 27132 40068 27188 41580
rect 27468 40850 27524 41580
rect 27468 40798 27470 40850
rect 27522 40798 27524 40850
rect 27468 40786 27524 40798
rect 27132 39954 27188 40012
rect 27132 39902 27134 39954
rect 27186 39902 27188 39954
rect 27132 39890 27188 39902
rect 27580 40626 27636 40638
rect 27580 40574 27582 40626
rect 27634 40574 27636 40626
rect 27580 39844 27636 40574
rect 27692 39956 27748 41804
rect 27692 39890 27748 39900
rect 27580 39778 27636 39788
rect 27916 39620 27972 39630
rect 27020 39618 27972 39620
rect 27020 39566 27918 39618
rect 27970 39566 27972 39618
rect 27020 39564 27972 39566
rect 27020 37938 27076 39564
rect 27916 39554 27972 39564
rect 27132 39284 27188 39294
rect 27132 38722 27188 39228
rect 28028 38948 28084 38958
rect 27916 38946 28084 38948
rect 27916 38894 28030 38946
rect 28082 38894 28084 38946
rect 27916 38892 28084 38894
rect 27580 38836 27636 38846
rect 27580 38742 27636 38780
rect 27132 38670 27134 38722
rect 27186 38670 27188 38722
rect 27132 38658 27188 38670
rect 27244 38722 27300 38734
rect 27244 38670 27246 38722
rect 27298 38670 27300 38722
rect 27020 37886 27022 37938
rect 27074 37886 27076 37938
rect 27020 37874 27076 37886
rect 27244 37716 27300 38670
rect 27804 38612 27860 38622
rect 27468 38610 27860 38612
rect 27468 38558 27806 38610
rect 27858 38558 27860 38610
rect 27468 38556 27860 38558
rect 27468 38162 27524 38556
rect 27804 38546 27860 38556
rect 27468 38110 27470 38162
rect 27522 38110 27524 38162
rect 27468 38098 27524 38110
rect 27244 37650 27300 37660
rect 27356 36708 27412 36718
rect 27356 36148 27412 36652
rect 27020 35924 27076 35934
rect 27020 35830 27076 35868
rect 27132 35364 27188 35374
rect 27132 34690 27188 35308
rect 27356 34802 27412 36092
rect 27356 34750 27358 34802
rect 27410 34750 27412 34802
rect 27356 34738 27412 34750
rect 27132 34638 27134 34690
rect 27186 34638 27188 34690
rect 27132 34626 27188 34638
rect 27580 34690 27636 34702
rect 27580 34638 27582 34690
rect 27634 34638 27636 34690
rect 27580 34020 27636 34638
rect 27580 33954 27636 33964
rect 27132 33908 27188 33918
rect 26908 33852 27132 33908
rect 27132 33814 27188 33852
rect 27692 33796 27748 33806
rect 27692 33702 27748 33740
rect 27916 33570 27972 38892
rect 28028 38882 28084 38892
rect 28140 38724 28196 43652
rect 28588 42868 28644 42878
rect 28588 41970 28644 42812
rect 29260 42082 29316 43652
rect 29260 42030 29262 42082
rect 29314 42030 29316 42082
rect 29260 42018 29316 42030
rect 29372 42642 29428 42654
rect 29372 42590 29374 42642
rect 29426 42590 29428 42642
rect 28588 41918 28590 41970
rect 28642 41918 28644 41970
rect 28588 41906 28644 41918
rect 29372 40852 29428 42590
rect 29260 40796 29428 40852
rect 29484 40852 29540 40862
rect 29260 40516 29316 40796
rect 29372 40628 29428 40638
rect 29372 40534 29428 40572
rect 29260 40450 29316 40460
rect 28476 40068 28532 40078
rect 28476 39842 28532 40012
rect 29260 39956 29316 39966
rect 29260 39862 29316 39900
rect 28476 39790 28478 39842
rect 28530 39790 28532 39842
rect 28364 39618 28420 39630
rect 28364 39566 28366 39618
rect 28418 39566 28420 39618
rect 28364 39284 28420 39566
rect 28364 39218 28420 39228
rect 28476 39060 28532 39790
rect 28812 39508 28868 39518
rect 28028 38668 28196 38724
rect 28364 39004 28532 39060
rect 28588 39506 28868 39508
rect 28588 39454 28814 39506
rect 28866 39454 28868 39506
rect 28588 39452 28868 39454
rect 28364 38948 28420 39004
rect 28028 35364 28084 38668
rect 28252 38610 28308 38622
rect 28252 38558 28254 38610
rect 28306 38558 28308 38610
rect 28252 38388 28308 38558
rect 28252 38322 28308 38332
rect 28364 38164 28420 38892
rect 28476 38836 28532 38846
rect 28588 38836 28644 39452
rect 28812 39442 28868 39452
rect 29372 38948 29428 38958
rect 29484 38948 29540 40796
rect 29372 38946 29540 38948
rect 29372 38894 29374 38946
rect 29426 38894 29540 38946
rect 29372 38892 29540 38894
rect 29372 38882 29428 38892
rect 28476 38834 28644 38836
rect 28476 38782 28478 38834
rect 28530 38782 28644 38834
rect 28476 38780 28644 38782
rect 28476 38770 28532 38780
rect 29596 38668 29652 59200
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 35196 55468 35460 55478
rect 35252 55412 35300 55468
rect 35356 55412 35404 55468
rect 35196 55402 35460 55412
rect 50556 54460 50820 54470
rect 50612 54404 50660 54460
rect 50716 54404 50764 54460
rect 50556 54394 50820 54404
rect 55244 54178 55300 54190
rect 55244 54126 55246 54178
rect 55298 54126 55300 54178
rect 55244 53844 55300 54126
rect 55244 53778 55300 53788
rect 35196 53452 35460 53462
rect 35252 53396 35300 53452
rect 35356 53396 35404 53452
rect 35196 53386 35460 53396
rect 50556 52444 50820 52454
rect 50612 52388 50660 52444
rect 50716 52388 50764 52444
rect 50556 52378 50820 52388
rect 35196 51436 35460 51446
rect 35252 51380 35300 51436
rect 35356 51380 35404 51436
rect 35196 51370 35460 51380
rect 50556 50428 50820 50438
rect 50612 50372 50660 50428
rect 50716 50372 50764 50428
rect 50556 50362 50820 50372
rect 36988 49810 37044 49822
rect 36988 49758 36990 49810
rect 37042 49758 37044 49810
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 36988 49028 37044 49758
rect 41356 49810 41412 49822
rect 41356 49758 41358 49810
rect 41410 49758 41412 49810
rect 36764 48972 36988 49028
rect 31276 48916 31332 48926
rect 30828 48804 30884 48814
rect 30828 48710 30884 48748
rect 30492 46786 30548 46798
rect 30492 46734 30494 46786
rect 30546 46734 30548 46786
rect 29708 46676 29764 46686
rect 29708 46582 29764 46620
rect 30156 46676 30212 46686
rect 30492 46676 30548 46734
rect 30156 46674 30996 46676
rect 30156 46622 30158 46674
rect 30210 46622 30996 46674
rect 30156 46620 30996 46622
rect 30156 46562 30212 46620
rect 30156 46510 30158 46562
rect 30210 46510 30212 46562
rect 30156 46498 30212 46510
rect 30940 46114 30996 46620
rect 30940 46062 30942 46114
rect 30994 46062 30996 46114
rect 30940 45444 30996 46062
rect 30940 45378 30996 45388
rect 30268 45332 30324 45342
rect 29932 44884 29988 44894
rect 29932 44790 29988 44828
rect 30268 44882 30324 45276
rect 30268 44830 30270 44882
rect 30322 44830 30324 44882
rect 29932 43988 29988 43998
rect 29932 43708 29988 43932
rect 30268 43708 30324 44830
rect 29932 43652 30324 43708
rect 31276 45332 31332 48860
rect 32732 48916 32788 48926
rect 32732 48822 32788 48860
rect 31948 48804 32004 48814
rect 31500 46786 31556 46798
rect 31500 46734 31502 46786
rect 31554 46734 31556 46786
rect 31500 46676 31556 46734
rect 31500 46610 31556 46620
rect 31948 45780 32004 48748
rect 34860 48690 34916 48702
rect 34860 48638 34862 48690
rect 34914 48638 34916 48690
rect 34860 47236 34916 48638
rect 36428 48690 36484 48702
rect 36428 48638 36430 48690
rect 36482 48638 36484 48690
rect 35420 47794 35476 47806
rect 35420 47742 35422 47794
rect 35474 47742 35476 47794
rect 35420 47570 35476 47742
rect 35868 47796 35924 47806
rect 36316 47796 36372 47806
rect 36428 47796 36484 48638
rect 36764 47908 36820 48972
rect 36988 48962 37044 48972
rect 37436 49028 37492 49038
rect 37436 48802 37492 48972
rect 37436 48750 37438 48802
rect 37490 48750 37492 48802
rect 37436 48738 37492 48750
rect 40348 49028 40404 49038
rect 38108 48690 38164 48702
rect 38108 48638 38110 48690
rect 38162 48638 38164 48690
rect 35868 47794 36036 47796
rect 35868 47742 35870 47794
rect 35922 47742 36036 47794
rect 35868 47740 36036 47742
rect 35868 47730 35924 47740
rect 35420 47518 35422 47570
rect 35474 47518 35476 47570
rect 35420 47506 35476 47518
rect 35868 47570 35924 47582
rect 35868 47518 35870 47570
rect 35922 47518 35924 47570
rect 35196 47404 35460 47414
rect 35252 47348 35300 47404
rect 35356 47348 35404 47404
rect 35196 47338 35460 47348
rect 34860 47234 35028 47236
rect 34860 47182 34862 47234
rect 34914 47182 35028 47234
rect 34860 47180 35028 47182
rect 34860 47170 34916 47180
rect 31276 43764 31332 45276
rect 31836 45666 31892 45678
rect 31836 45614 31838 45666
rect 31890 45614 31892 45666
rect 31836 44324 31892 45614
rect 31948 44884 32004 45724
rect 31948 44818 32004 44828
rect 32620 46676 32676 46686
rect 32620 44882 32676 46620
rect 33180 45780 33236 45790
rect 33292 45780 33348 45790
rect 33180 45778 33292 45780
rect 33180 45726 33182 45778
rect 33234 45726 33292 45778
rect 33180 45724 33292 45726
rect 33180 45714 33236 45724
rect 32620 44830 32622 44882
rect 32674 44830 32676 44882
rect 32620 44818 32676 44830
rect 33180 45332 33236 45342
rect 33180 44882 33236 45276
rect 33180 44830 33182 44882
rect 33234 44830 33236 44882
rect 31836 44268 32116 44324
rect 32060 43988 32116 44268
rect 33180 44100 33236 44830
rect 32060 43932 32452 43988
rect 31276 43698 31332 43708
rect 32284 43764 32340 43802
rect 32284 43698 32340 43708
rect 31388 43652 31444 43662
rect 29820 42644 29876 42654
rect 29820 42550 29876 42588
rect 29820 40740 29876 40750
rect 29932 40740 29988 43652
rect 31388 43650 31780 43652
rect 31388 43598 31390 43650
rect 31442 43598 31780 43650
rect 31388 43596 31780 43598
rect 31388 43586 31444 43596
rect 31724 42866 31780 43596
rect 31724 42814 31726 42866
rect 31778 42814 31780 42866
rect 31724 42802 31780 42814
rect 32396 42866 32452 43932
rect 33180 43764 33236 44044
rect 33292 44098 33348 45724
rect 34636 45780 34692 45790
rect 34636 45686 34692 45724
rect 34972 45220 35028 47180
rect 35084 45892 35140 45902
rect 35084 45798 35140 45836
rect 35868 45890 35924 47518
rect 35868 45838 35870 45890
rect 35922 45838 35924 45890
rect 35532 45778 35588 45790
rect 35532 45726 35534 45778
rect 35586 45726 35588 45778
rect 35196 45388 35460 45398
rect 35252 45332 35300 45388
rect 35356 45332 35404 45388
rect 35196 45322 35460 45332
rect 34972 45164 35252 45220
rect 33292 44046 33294 44098
rect 33346 44046 33348 44098
rect 33292 44034 33348 44046
rect 33628 44658 33684 44670
rect 33628 44606 33630 44658
rect 33682 44606 33684 44658
rect 33516 43876 33572 43886
rect 33516 43782 33572 43820
rect 33180 43698 33236 43708
rect 33628 43708 33684 44606
rect 34412 44100 34468 44110
rect 34300 43988 34356 43998
rect 34412 43988 34468 44044
rect 34300 43986 34468 43988
rect 34300 43934 34302 43986
rect 34354 43934 34468 43986
rect 34300 43932 34468 43934
rect 34300 43922 34356 43932
rect 33628 43652 33908 43708
rect 32396 42814 32398 42866
rect 32450 42814 32452 42866
rect 32396 42802 32452 42814
rect 33852 42866 33908 43652
rect 33852 42814 33854 42866
rect 33906 42814 33908 42866
rect 33852 42802 33908 42814
rect 32060 42754 32116 42766
rect 32060 42702 32062 42754
rect 32114 42702 32116 42754
rect 32060 41972 32116 42702
rect 33292 42756 33348 42766
rect 33292 42662 33348 42700
rect 32060 41906 32116 41916
rect 32732 42642 32788 42654
rect 32732 42590 32734 42642
rect 32786 42590 32788 42642
rect 30044 41860 30100 41870
rect 30100 41804 30436 41860
rect 30044 41766 30100 41804
rect 30380 40964 30436 41804
rect 30492 41748 30548 41758
rect 30548 41692 30660 41748
rect 30492 41654 30548 41692
rect 30380 40852 30436 40908
rect 30492 40852 30548 40862
rect 30380 40850 30548 40852
rect 30380 40798 30494 40850
rect 30546 40798 30548 40850
rect 30380 40796 30548 40798
rect 30492 40786 30548 40796
rect 29876 40684 29988 40740
rect 29820 40646 29876 40684
rect 30268 40626 30324 40638
rect 30268 40574 30270 40626
rect 30322 40574 30324 40626
rect 29820 40404 29876 40414
rect 29820 39954 29876 40348
rect 29820 39902 29822 39954
rect 29874 39902 29876 39954
rect 29820 39890 29876 39902
rect 30268 40292 30324 40574
rect 30268 39956 30324 40236
rect 30380 39956 30436 39966
rect 30268 39954 30436 39956
rect 30268 39902 30382 39954
rect 30434 39902 30436 39954
rect 30268 39900 30436 39902
rect 29932 39732 29988 39742
rect 29372 38612 29652 38668
rect 29820 39730 29988 39732
rect 29820 39678 29934 39730
rect 29986 39678 29988 39730
rect 29820 39676 29988 39678
rect 28252 38108 28644 38164
rect 28140 38052 28196 38062
rect 28252 38052 28308 38108
rect 28140 38050 28308 38052
rect 28140 37998 28142 38050
rect 28194 37998 28308 38050
rect 28140 37996 28308 37998
rect 28588 38050 28644 38108
rect 28588 37998 28590 38050
rect 28642 37998 28644 38050
rect 28140 37986 28196 37996
rect 28588 37986 28644 37998
rect 29372 36820 29428 38612
rect 29260 36708 29316 36718
rect 29260 36614 29316 36652
rect 29372 36706 29428 36764
rect 29372 36654 29374 36706
rect 29426 36654 29428 36706
rect 29372 36642 29428 36654
rect 28588 36594 28644 36606
rect 28588 36542 28590 36594
rect 28642 36542 28644 36594
rect 28084 35308 28196 35364
rect 28028 35298 28084 35308
rect 28028 34468 28084 34478
rect 28028 34374 28084 34412
rect 28140 34018 28196 35308
rect 28140 33966 28142 34018
rect 28194 33966 28196 34018
rect 28140 33954 28196 33966
rect 28588 34580 28644 36542
rect 29372 35812 29428 35822
rect 29260 35810 29428 35812
rect 29260 35758 29374 35810
rect 29426 35758 29428 35810
rect 29260 35756 29428 35758
rect 28588 33796 28644 34524
rect 29036 35586 29092 35598
rect 29036 35534 29038 35586
rect 29090 35534 29092 35586
rect 28700 33796 28756 33806
rect 28588 33740 28700 33796
rect 28700 33702 28756 33740
rect 29036 33684 29092 35534
rect 29260 34802 29316 35756
rect 29372 35746 29428 35756
rect 29260 34750 29262 34802
rect 29314 34750 29316 34802
rect 29260 34580 29316 34750
rect 29260 34514 29316 34524
rect 29484 34468 29540 34478
rect 29484 34018 29540 34412
rect 29484 33966 29486 34018
rect 29538 33966 29540 34018
rect 29484 33954 29540 33966
rect 29036 33618 29092 33628
rect 27916 33518 27918 33570
rect 27970 33518 27972 33570
rect 27916 33506 27972 33518
rect 27244 33458 27300 33470
rect 27244 33406 27246 33458
rect 27298 33406 27300 33458
rect 27020 32788 27076 32798
rect 27020 32694 27076 32732
rect 27244 32786 27300 33406
rect 27916 33124 27972 33134
rect 27244 32734 27246 32786
rect 27298 32734 27300 32786
rect 27244 32722 27300 32734
rect 27804 33068 27916 33124
rect 27804 32786 27860 33068
rect 27916 33058 27972 33068
rect 28364 33124 28420 33134
rect 28364 32898 28420 33068
rect 28364 32846 28366 32898
rect 28418 32846 28420 32898
rect 28364 32834 28420 32846
rect 28588 32788 28644 32798
rect 27804 32734 27806 32786
rect 27858 32734 27860 32786
rect 27804 32722 27860 32734
rect 28476 32732 28588 32788
rect 26684 32674 26740 32686
rect 26684 32622 26686 32674
rect 26738 32622 26740 32674
rect 26684 31108 26740 32622
rect 27580 32674 27636 32686
rect 27580 32622 27582 32674
rect 27634 32622 27636 32674
rect 26796 32564 26852 32574
rect 26796 32562 26964 32564
rect 26796 32510 26798 32562
rect 26850 32510 26964 32562
rect 26796 32508 26964 32510
rect 26796 32498 26852 32508
rect 26908 32004 26964 32508
rect 26684 31042 26740 31052
rect 26796 31948 26964 32004
rect 27020 32228 27076 32238
rect 26684 30548 26740 30558
rect 26684 30454 26740 30492
rect 26796 30324 26852 31948
rect 27020 31834 27076 32172
rect 27580 32228 27636 32622
rect 27692 32452 27748 32462
rect 27692 32358 27748 32396
rect 27636 32172 27972 32228
rect 27580 32134 27636 32172
rect 27020 31782 27022 31834
rect 27074 31782 27076 31834
rect 27356 32004 27412 32014
rect 27356 31792 27412 31948
rect 27916 32004 27972 32172
rect 28364 32004 28420 32014
rect 28476 32004 28532 32732
rect 28588 32722 28644 32732
rect 27916 32002 28084 32004
rect 27916 31950 27918 32002
rect 27970 31950 28084 32002
rect 27916 31948 28084 31950
rect 27916 31938 27972 31948
rect 27580 31892 27636 31902
rect 27020 31770 27076 31782
rect 27242 31778 27412 31792
rect 27242 31726 27246 31778
rect 27298 31736 27412 31778
rect 27468 31890 27636 31892
rect 27468 31838 27582 31890
rect 27634 31838 27636 31890
rect 27468 31836 27636 31838
rect 27468 31780 27524 31836
rect 27580 31826 27636 31836
rect 27298 31726 27300 31736
rect 27242 31724 27300 31726
rect 27244 31714 27300 31724
rect 27020 31668 27076 31678
rect 26908 31444 26964 31454
rect 26908 31350 26964 31388
rect 26908 30660 26964 30670
rect 26908 30566 26964 30604
rect 27020 30658 27076 31612
rect 27020 30606 27022 30658
rect 27074 30606 27076 30658
rect 26572 30268 26740 30324
rect 26460 30046 26462 30098
rect 26514 30046 26516 30098
rect 26460 30034 26516 30046
rect 25788 29988 25844 29998
rect 25564 29876 25620 29886
rect 25564 29782 25620 29820
rect 25676 29874 25732 29886
rect 25676 29822 25678 29874
rect 25730 29822 25732 29874
rect 25676 29764 25732 29822
rect 25676 29698 25732 29708
rect 25452 28644 25508 28654
rect 25676 28644 25732 28654
rect 25340 28642 25508 28644
rect 25340 28590 25454 28642
rect 25506 28590 25508 28642
rect 25340 28588 25508 28590
rect 25452 28578 25508 28588
rect 25564 28642 25732 28644
rect 25564 28590 25678 28642
rect 25730 28590 25732 28642
rect 25564 28588 25732 28590
rect 24892 27906 24948 27916
rect 25116 28140 25284 28196
rect 24668 27748 24724 27758
rect 24668 27654 24724 27692
rect 24556 26786 24612 26796
rect 25116 26850 25172 28140
rect 25564 28084 25620 28588
rect 25676 28578 25732 28588
rect 25788 28418 25844 29932
rect 26012 29932 26292 29988
rect 26012 28866 26068 29932
rect 26012 28814 26014 28866
rect 26066 28814 26068 28866
rect 26012 28802 26068 28814
rect 26124 29762 26180 29774
rect 26124 29710 26126 29762
rect 26178 29710 26180 29762
rect 26124 28644 26180 29710
rect 26236 29762 26292 29932
rect 26236 29710 26238 29762
rect 26290 29710 26292 29762
rect 26236 29698 26292 29710
rect 26572 29874 26628 29886
rect 26572 29822 26574 29874
rect 26626 29822 26628 29874
rect 26572 29764 26628 29822
rect 26572 29698 26628 29708
rect 26348 28868 26404 28878
rect 26348 28754 26404 28812
rect 26348 28702 26350 28754
rect 26402 28702 26404 28754
rect 26348 28690 26404 28702
rect 26124 28588 26292 28644
rect 25900 28532 25956 28542
rect 25900 28438 25956 28476
rect 25788 28366 25790 28418
rect 25842 28366 25844 28418
rect 25788 28354 25844 28366
rect 26124 28420 26180 28430
rect 25340 28028 25620 28084
rect 25228 27972 25284 27982
rect 25228 27878 25284 27916
rect 25116 26798 25118 26850
rect 25170 26798 25172 26850
rect 25116 26786 25172 26798
rect 25228 27076 25284 27086
rect 24444 26686 24446 26738
rect 24498 26686 24500 26738
rect 24220 26626 24276 26638
rect 24220 26574 24222 26626
rect 24274 26574 24276 26626
rect 24220 26292 24276 26574
rect 24332 26404 24388 26414
rect 24332 26310 24388 26348
rect 24220 26226 24276 26236
rect 24444 26068 24500 26686
rect 24668 26740 24724 26750
rect 24668 26646 24724 26684
rect 25004 26740 25060 26750
rect 24444 26002 24500 26012
rect 24556 26628 24612 26638
rect 24444 25842 24500 25854
rect 24444 25790 24446 25842
rect 24498 25790 24500 25842
rect 23772 21870 23774 21922
rect 23826 21870 23828 21922
rect 23772 21858 23828 21870
rect 23884 24332 24052 24388
rect 24108 24722 24164 24734
rect 24108 24670 24110 24722
rect 24162 24670 24164 24722
rect 23212 21810 23268 21822
rect 23212 21758 23214 21810
rect 23266 21758 23268 21810
rect 23212 21700 23268 21758
rect 23212 21634 23268 21644
rect 23100 21420 23380 21476
rect 22876 20802 23044 20804
rect 22876 20750 22878 20802
rect 22930 20750 23044 20802
rect 22876 20748 23044 20750
rect 23324 20804 23380 21420
rect 23772 20804 23828 20814
rect 23324 20802 23772 20804
rect 23324 20750 23326 20802
rect 23378 20750 23772 20802
rect 23324 20748 23772 20750
rect 22764 20244 22820 20254
rect 22204 19842 22260 19852
rect 22316 20132 22372 20142
rect 21756 19796 21812 19806
rect 21812 19740 21924 19796
rect 21756 19730 21812 19740
rect 21476 18732 21700 18788
rect 21868 18786 21924 19740
rect 22316 18788 22372 20076
rect 22764 19794 22820 20188
rect 22876 20132 22932 20748
rect 23324 20738 23380 20748
rect 23772 20710 23828 20748
rect 22876 20066 22932 20076
rect 22764 19742 22766 19794
rect 22818 19742 22820 19794
rect 22764 19730 22820 19742
rect 22764 19348 22820 19358
rect 21868 18734 21870 18786
rect 21922 18734 21924 18786
rect 20076 17836 20356 17892
rect 20748 18564 20804 18574
rect 20748 17890 20804 18508
rect 21420 18562 21476 18732
rect 21420 18510 21422 18562
rect 21474 18510 21476 18562
rect 21420 18004 21476 18510
rect 20748 17838 20750 17890
rect 20802 17838 20804 17890
rect 19516 16828 19908 16884
rect 19964 17668 20020 17678
rect 19292 16772 19348 16782
rect 18620 16660 18676 16670
rect 18620 15538 18676 16604
rect 19180 16324 19236 16334
rect 19180 16230 19236 16268
rect 19292 15762 19348 16716
rect 19292 15710 19294 15762
rect 19346 15710 19348 15762
rect 19292 15698 19348 15710
rect 18956 15652 19012 15662
rect 19516 15652 19572 16828
rect 19964 16772 20020 17612
rect 19628 16716 20020 16772
rect 20076 17666 20132 17836
rect 20748 17826 20804 17838
rect 21196 17948 21476 18004
rect 20076 17614 20078 17666
rect 20130 17614 20132 17666
rect 20076 16772 20132 17614
rect 20412 17668 20468 17678
rect 20412 17574 20468 17612
rect 19628 15876 19684 16716
rect 20076 16706 20132 16716
rect 20748 16770 20804 16782
rect 20748 16718 20750 16770
rect 20802 16718 20804 16770
rect 20524 16660 20580 16670
rect 20188 16436 20244 16446
rect 20188 16342 20244 16380
rect 19836 16156 20100 16166
rect 19892 16100 19940 16156
rect 19996 16100 20044 16156
rect 19836 16090 20100 16100
rect 19964 15876 20020 15886
rect 19628 15874 20020 15876
rect 19628 15822 19966 15874
rect 20018 15822 20020 15874
rect 19628 15820 20020 15822
rect 19964 15810 20020 15820
rect 20524 15762 20580 16604
rect 20748 15876 20804 16718
rect 20748 15810 20804 15820
rect 21084 16324 21140 16334
rect 20524 15710 20526 15762
rect 20578 15710 20580 15762
rect 20524 15698 20580 15710
rect 21084 15762 21140 16268
rect 21084 15710 21086 15762
rect 21138 15710 21140 15762
rect 21084 15698 21140 15710
rect 19628 15652 19684 15662
rect 18956 15650 19124 15652
rect 18956 15598 18958 15650
rect 19010 15598 19124 15650
rect 18956 15596 19124 15598
rect 19516 15650 19684 15652
rect 19516 15598 19630 15650
rect 19682 15598 19684 15650
rect 19516 15596 19684 15598
rect 18956 15586 19012 15596
rect 18620 15486 18622 15538
rect 18674 15486 18676 15538
rect 18620 15426 18676 15486
rect 18620 15374 18622 15426
rect 18674 15374 18676 15426
rect 18620 14642 18676 15374
rect 19068 14978 19124 15596
rect 19628 15586 19684 15596
rect 20860 15652 20916 15662
rect 21196 15652 21252 17948
rect 21868 17892 21924 18734
rect 21420 17836 21924 17892
rect 22204 18786 22372 18788
rect 22204 18734 22318 18786
rect 22370 18734 22372 18786
rect 22204 18732 22372 18734
rect 21308 17666 21364 17678
rect 21308 17614 21310 17666
rect 21362 17614 21364 17666
rect 21308 16660 21364 17614
rect 21308 16594 21364 16604
rect 21420 16658 21476 17836
rect 21868 17668 21924 17678
rect 21420 16606 21422 16658
rect 21474 16606 21476 16658
rect 21308 15652 21364 15662
rect 21196 15596 21308 15652
rect 19068 14926 19070 14978
rect 19122 14926 19124 14978
rect 19068 14914 19124 14926
rect 20300 14756 20356 14766
rect 20300 14662 20356 14700
rect 18620 14590 18622 14642
rect 18674 14590 18676 14642
rect 18620 13524 18676 14590
rect 19852 14420 19908 14430
rect 19852 14326 19908 14364
rect 20748 14420 20804 14430
rect 20860 14420 20916 15596
rect 21308 15586 21364 15596
rect 20748 14418 20916 14420
rect 20748 14366 20750 14418
rect 20802 14366 20916 14418
rect 20748 14364 20916 14366
rect 20748 14354 20804 14364
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 18620 13458 18676 13468
rect 19404 13524 19460 13534
rect 19404 13430 19460 13468
rect 20524 13522 20580 13534
rect 20524 13470 20526 13522
rect 20578 13470 20580 13522
rect 18284 12462 18286 12514
rect 18338 12462 18340 12514
rect 18284 12292 18340 12462
rect 17948 11732 18004 11742
rect 18284 11732 18340 12236
rect 19836 12124 20100 12134
rect 19892 12068 19940 12124
rect 19996 12068 20044 12124
rect 19836 12058 20100 12068
rect 17948 11730 18340 11732
rect 17948 11678 17950 11730
rect 18002 11678 18340 11730
rect 17948 11676 18340 11678
rect 17948 11666 18004 11676
rect 17500 11566 17502 11618
rect 17554 11566 17556 11618
rect 4476 11116 4740 11126
rect 4532 11060 4580 11116
rect 4636 11060 4684 11116
rect 4476 11050 4740 11060
rect 16940 10610 16996 10622
rect 16940 10558 16942 10610
rect 16994 10558 16996 10610
rect 16380 10498 16436 10510
rect 16380 10446 16382 10498
rect 16434 10446 16436 10498
rect 16380 10164 16436 10446
rect 16380 10098 16436 10108
rect 16940 10052 16996 10558
rect 17500 10164 17556 11566
rect 17500 10098 17556 10108
rect 16940 9986 16996 9996
rect 18284 10052 18340 11676
rect 19852 11730 19908 11742
rect 19852 11678 19854 11730
rect 19906 11678 19908 11730
rect 19068 10612 19124 10622
rect 19068 10518 19124 10556
rect 19852 10612 19908 11678
rect 19852 10546 19908 10556
rect 19740 10388 19796 10398
rect 19740 10294 19796 10332
rect 18396 10164 18452 10174
rect 18452 10108 18564 10164
rect 18396 10098 18452 10108
rect 18284 9492 18340 9996
rect 18284 9426 18340 9436
rect 18508 9490 18564 10108
rect 19836 10108 20100 10118
rect 19892 10052 19940 10108
rect 19996 10052 20044 10108
rect 19836 10042 20100 10052
rect 20188 9714 20244 9726
rect 20188 9662 20190 9714
rect 20242 9662 20244 9714
rect 19628 9604 19684 9614
rect 19852 9604 19908 9614
rect 19292 9548 19628 9604
rect 18508 9438 18510 9490
rect 18562 9438 18564 9490
rect 4476 9100 4740 9110
rect 4532 9044 4580 9100
rect 4636 9044 4684 9100
rect 4476 9034 4740 9044
rect 18508 8484 18564 9438
rect 18956 9492 19012 9502
rect 18956 9398 19012 9436
rect 18956 8484 19012 8522
rect 18508 8428 18956 8484
rect 18956 8418 19012 8428
rect 19292 8428 19348 9548
rect 19628 9510 19684 9548
rect 19740 9602 19908 9604
rect 19740 9550 19854 9602
rect 19906 9550 19908 9602
rect 19740 9548 19908 9550
rect 19516 8820 19572 8830
rect 19404 8596 19460 8606
rect 19516 8596 19572 8764
rect 19404 8594 19572 8596
rect 19404 8542 19406 8594
rect 19458 8542 19572 8594
rect 19404 8540 19572 8542
rect 19404 8530 19460 8540
rect 19292 8372 19460 8428
rect 19404 7586 19460 8372
rect 19404 7534 19406 7586
rect 19458 7534 19460 7586
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4620 6804 4676 6814
rect 4172 6356 4228 6366
rect 4172 6262 4228 6300
rect 4620 6354 4676 6748
rect 19404 6580 19460 7534
rect 19516 7586 19572 8540
rect 19740 8484 19796 9548
rect 19852 9538 19908 9548
rect 20188 9492 20244 9662
rect 19852 8708 19908 8718
rect 19852 8614 19908 8652
rect 20188 8596 20244 9436
rect 20300 9604 20356 9614
rect 20300 8706 20356 9548
rect 20524 8820 20580 13470
rect 20636 12514 20692 12526
rect 20636 12462 20638 12514
rect 20690 12462 20692 12514
rect 20636 11508 20692 12462
rect 20636 11442 20692 11452
rect 20636 10836 20692 10846
rect 20636 10722 20692 10780
rect 20636 10670 20638 10722
rect 20690 10670 20692 10722
rect 20636 9604 20692 10670
rect 20636 9538 20692 9548
rect 20524 8754 20580 8764
rect 20300 8654 20302 8706
rect 20354 8654 20356 8706
rect 20300 8642 20356 8654
rect 20860 8708 20916 14364
rect 20972 14756 21028 14766
rect 20972 13860 21028 14700
rect 21420 14308 21476 16606
rect 21756 17666 21924 17668
rect 21756 17614 21870 17666
rect 21922 17614 21924 17666
rect 21756 17612 21924 17614
rect 21756 16434 21812 17612
rect 21868 17602 21924 17612
rect 21980 16772 22036 16782
rect 21756 16382 21758 16434
rect 21810 16382 21812 16434
rect 21756 16370 21812 16382
rect 21868 16658 21924 16670
rect 21868 16606 21870 16658
rect 21922 16606 21924 16658
rect 21868 16436 21924 16606
rect 21868 16370 21924 16380
rect 21644 15876 21700 15886
rect 21700 15820 21812 15876
rect 21644 15810 21700 15820
rect 21756 15762 21812 15820
rect 21756 15710 21758 15762
rect 21810 15710 21812 15762
rect 21756 15698 21812 15710
rect 21420 13860 21476 14252
rect 21980 13970 22036 16716
rect 22204 16660 22260 18732
rect 22316 18722 22372 18732
rect 22540 19346 22820 19348
rect 22540 19294 22766 19346
rect 22818 19294 22820 19346
rect 22540 19292 22820 19294
rect 22540 17890 22596 19292
rect 22764 19282 22820 19292
rect 23212 18900 23268 18910
rect 23212 18674 23268 18844
rect 23212 18622 23214 18674
rect 23266 18622 23268 18674
rect 23212 18610 23268 18622
rect 23884 18674 23940 24332
rect 24108 24164 24164 24670
rect 23996 24108 24164 24164
rect 24332 24610 24388 24622
rect 24332 24558 24334 24610
rect 24386 24558 24388 24610
rect 23996 23940 24052 24108
rect 23996 23874 24052 23884
rect 24108 23940 24164 23950
rect 24332 23940 24388 24558
rect 24108 23938 24388 23940
rect 24108 23886 24110 23938
rect 24162 23886 24388 23938
rect 24108 23884 24388 23886
rect 24108 23874 24164 23884
rect 24332 23828 24388 23884
rect 24332 23762 24388 23772
rect 23884 18622 23886 18674
rect 23938 18622 23940 18674
rect 23884 18610 23940 18622
rect 23996 23716 24052 23726
rect 22876 18564 22932 18574
rect 22876 18470 22932 18508
rect 23548 18562 23604 18574
rect 23548 18510 23550 18562
rect 23602 18510 23604 18562
rect 22540 17838 22542 17890
rect 22594 17838 22596 17890
rect 22540 17826 22596 17838
rect 23548 17892 23604 18510
rect 23996 18564 24052 23660
rect 24444 23716 24500 25790
rect 24556 25844 24612 26572
rect 25004 26626 25060 26684
rect 25004 26574 25006 26626
rect 25058 26574 25060 26626
rect 25004 26562 25060 26574
rect 25228 26626 25284 27020
rect 25228 26574 25230 26626
rect 25282 26574 25284 26626
rect 25228 26562 25284 26574
rect 25116 26068 25172 26078
rect 25172 26012 25284 26068
rect 25116 26002 25172 26012
rect 25228 25954 25284 26012
rect 25228 25902 25230 25954
rect 25282 25902 25284 25954
rect 25228 25890 25284 25902
rect 24556 25788 24836 25844
rect 24556 25620 24612 25630
rect 24556 25526 24612 25564
rect 24668 24724 24724 24734
rect 24556 24612 24612 24622
rect 24556 24518 24612 24556
rect 24444 23650 24500 23660
rect 24556 23940 24612 23950
rect 24668 23940 24724 24668
rect 24556 23938 24724 23940
rect 24556 23886 24558 23938
rect 24610 23886 24724 23938
rect 24556 23884 24724 23886
rect 24332 22596 24388 22606
rect 24556 22596 24612 23884
rect 24668 23492 24724 23502
rect 24668 23398 24724 23436
rect 24332 22594 24612 22596
rect 24332 22542 24334 22594
rect 24386 22542 24612 22594
rect 24332 22540 24612 22542
rect 24668 22706 24724 22718
rect 24668 22654 24670 22706
rect 24722 22654 24724 22706
rect 24668 22596 24724 22654
rect 24332 22530 24388 22540
rect 24668 22530 24724 22540
rect 24668 21588 24724 21598
rect 24668 21494 24724 21532
rect 24220 21252 24276 21262
rect 24220 21026 24276 21196
rect 24220 20974 24222 21026
rect 24274 20974 24276 21026
rect 24220 20802 24276 20974
rect 24220 20750 24222 20802
rect 24274 20750 24276 20802
rect 24220 20738 24276 20750
rect 24668 20804 24724 20814
rect 24668 20710 24724 20748
rect 24108 20244 24164 20254
rect 24108 19906 24164 20188
rect 24780 20188 24836 25788
rect 24892 25732 24948 25742
rect 24892 25058 24948 25676
rect 25340 25508 25396 28028
rect 25564 27858 25620 27870
rect 25564 27806 25566 27858
rect 25618 27806 25620 27858
rect 25564 27636 25620 27806
rect 26124 27858 26180 28364
rect 26124 27806 26126 27858
rect 26178 27806 26180 27858
rect 26124 27794 26180 27806
rect 26012 27636 26068 27646
rect 25564 27634 26068 27636
rect 25564 27582 26014 27634
rect 26066 27582 26068 27634
rect 25564 27580 26068 27582
rect 25564 26738 25620 26750
rect 25564 26686 25566 26738
rect 25618 26686 25620 26738
rect 25564 26516 25620 26686
rect 25676 26740 25732 27580
rect 26012 27570 26068 27580
rect 25676 26646 25732 26684
rect 26012 26964 26068 26974
rect 26236 26908 26292 28588
rect 26572 28532 26628 28542
rect 26572 27972 26628 28476
rect 26684 28308 26740 30268
rect 26796 28530 26852 30268
rect 27020 30100 27076 30606
rect 27020 30034 27076 30044
rect 27132 31444 27188 31454
rect 26908 29874 26964 29886
rect 26908 29822 26910 29874
rect 26962 29822 26964 29874
rect 26908 28980 26964 29822
rect 27020 29874 27076 29886
rect 27020 29822 27022 29874
rect 27074 29822 27076 29874
rect 27020 29540 27076 29822
rect 27132 29876 27188 31388
rect 27356 30770 27412 30782
rect 27356 30718 27358 30770
rect 27410 30718 27412 30770
rect 27356 30324 27412 30718
rect 27356 30258 27412 30268
rect 27132 29810 27188 29820
rect 27468 29874 27524 31724
rect 27580 31108 27636 31118
rect 27580 31014 27636 31052
rect 27916 30772 27972 30782
rect 27916 30678 27972 30716
rect 27692 30658 27748 30670
rect 27692 30606 27694 30658
rect 27746 30606 27748 30658
rect 27692 30548 27748 30606
rect 28028 30660 28084 31948
rect 28420 31948 28532 32004
rect 28364 31910 28420 31948
rect 29820 31780 29876 39676
rect 29932 39666 29988 39676
rect 30044 38948 30100 38958
rect 30268 38948 30324 39900
rect 30380 39890 30436 39900
rect 30100 38892 30324 38948
rect 30604 38948 30660 41692
rect 32508 41746 32564 41758
rect 32508 41694 32510 41746
rect 32562 41694 32564 41746
rect 31612 40962 31668 40974
rect 31612 40910 31614 40962
rect 31666 40910 31668 40962
rect 30716 40850 30772 40862
rect 30716 40798 30718 40850
rect 30770 40798 30772 40850
rect 30716 40516 30772 40798
rect 30716 40450 30772 40460
rect 31164 40740 31220 40750
rect 30044 38854 30100 38892
rect 30604 38882 30660 38892
rect 30716 36820 30772 36830
rect 30716 36726 30772 36764
rect 29932 36706 29988 36718
rect 29932 36654 29934 36706
rect 29986 36654 29988 36706
rect 29932 32900 29988 36654
rect 30380 36484 30436 36494
rect 30044 36482 30436 36484
rect 30044 36430 30382 36482
rect 30434 36430 30436 36482
rect 30044 36428 30436 36430
rect 30044 34690 30100 36428
rect 30380 36418 30436 36428
rect 30156 36036 30212 36046
rect 30156 35942 30212 35980
rect 30044 34638 30046 34690
rect 30098 34638 30100 34690
rect 30044 34626 30100 34638
rect 29932 32834 29988 32844
rect 30716 33684 30772 33694
rect 29820 31714 29876 31724
rect 28252 30884 28308 30894
rect 28252 30790 28308 30828
rect 28588 30770 28644 30782
rect 28588 30718 28590 30770
rect 28642 30718 28644 30770
rect 28364 30660 28420 30670
rect 28028 30658 28420 30660
rect 28028 30606 28366 30658
rect 28418 30606 28420 30658
rect 28028 30604 28420 30606
rect 28028 30548 28084 30604
rect 28364 30594 28420 30604
rect 27692 30492 28084 30548
rect 28588 30436 28644 30718
rect 29708 30772 29764 30782
rect 30716 30772 30772 33628
rect 30940 31892 30996 31902
rect 31164 31892 31220 40684
rect 31612 40292 31668 40910
rect 32508 40740 32564 41694
rect 32732 41188 32788 42590
rect 34412 42308 34468 43932
rect 35084 43986 35140 43998
rect 35084 43934 35086 43986
rect 35138 43934 35140 43986
rect 35084 43708 35140 43934
rect 34524 43652 35140 43708
rect 34524 42754 34580 43652
rect 35196 43540 35252 45164
rect 35532 44660 35588 45726
rect 35868 45780 35924 45838
rect 35868 45714 35924 45724
rect 35980 45892 36036 47740
rect 36372 47740 36484 47796
rect 36652 47906 36820 47908
rect 36652 47854 36766 47906
rect 36818 47854 36820 47906
rect 36652 47852 36820 47854
rect 36316 45892 36372 47740
rect 36652 47570 36708 47852
rect 36764 47842 36820 47852
rect 37100 48018 37156 48030
rect 37100 47966 37102 48018
rect 37154 47966 37156 48018
rect 37100 47796 37156 47966
rect 37100 47730 37156 47740
rect 38108 47796 38164 48638
rect 40012 48692 40068 48702
rect 38108 47730 38164 47740
rect 39340 48018 39396 48030
rect 39340 47966 39342 48018
rect 39394 47966 39396 48018
rect 36652 47518 36654 47570
rect 36706 47518 36708 47570
rect 36652 47506 36708 47518
rect 38668 47122 38724 47134
rect 38668 47070 38670 47122
rect 38722 47070 38724 47122
rect 36428 45892 36484 45902
rect 36316 45890 36484 45892
rect 36316 45838 36430 45890
rect 36482 45838 36484 45890
rect 36316 45836 36484 45838
rect 35980 44996 36036 45836
rect 35756 44940 35980 44996
rect 35644 44660 35700 44670
rect 35532 44604 35644 44660
rect 35532 43876 35588 44604
rect 35644 44566 35700 44604
rect 35644 44100 35700 44110
rect 35756 44100 35812 44940
rect 35980 44930 36036 44940
rect 36092 45780 36148 45790
rect 35700 44044 35812 44100
rect 35644 44006 35700 44044
rect 35532 43810 35588 43820
rect 36092 43876 36148 45724
rect 36428 44660 36484 45836
rect 38556 45892 38612 45902
rect 38668 45892 38724 47070
rect 39340 47124 39396 47966
rect 39452 47124 39508 47134
rect 39340 47122 39508 47124
rect 39340 47070 39454 47122
rect 39506 47070 39508 47122
rect 39340 47068 39508 47070
rect 39452 47010 39508 47068
rect 40012 47122 40068 48636
rect 40012 47070 40014 47122
rect 40066 47070 40068 47122
rect 40012 47058 40068 47070
rect 40124 48690 40180 48702
rect 40124 48638 40126 48690
rect 40178 48638 40180 48690
rect 39452 46958 39454 47010
rect 39506 46958 39508 47010
rect 39452 46946 39508 46958
rect 39004 46900 39060 46910
rect 38892 46562 38948 46574
rect 38892 46510 38894 46562
rect 38946 46510 38948 46562
rect 38556 45890 38836 45892
rect 38556 45838 38558 45890
rect 38610 45838 38836 45890
rect 38556 45836 38836 45838
rect 38556 45826 38612 45836
rect 38332 45332 38388 45342
rect 37660 44996 37716 45006
rect 37660 44902 37716 44940
rect 38332 44770 38388 45276
rect 38332 44718 38334 44770
rect 38386 44718 38388 44770
rect 37212 44660 37268 44670
rect 36484 44604 36820 44660
rect 36428 44566 36484 44604
rect 36204 43876 36260 43886
rect 36092 43874 36260 43876
rect 36092 43822 36206 43874
rect 36258 43822 36260 43874
rect 36092 43820 36260 43822
rect 36092 43764 36148 43820
rect 36204 43810 36260 43820
rect 36764 43876 36820 44604
rect 36764 43782 36820 43820
rect 34524 42702 34526 42754
rect 34578 42702 34580 42754
rect 34524 42690 34580 42702
rect 35084 43484 35252 43540
rect 35868 43652 36148 43708
rect 37100 43764 37156 43774
rect 34412 42252 34804 42308
rect 33404 41972 33460 41982
rect 33404 41878 33460 41916
rect 34636 41972 34692 41982
rect 34636 41878 34692 41916
rect 32732 41122 32788 41132
rect 33068 41858 33124 41870
rect 33068 41806 33070 41858
rect 33122 41806 33124 41858
rect 32508 40674 32564 40684
rect 33068 40516 33124 41806
rect 33740 41860 33796 41870
rect 33740 41858 34020 41860
rect 33740 41806 33742 41858
rect 33794 41806 34020 41858
rect 33740 41804 34020 41806
rect 33740 41794 33796 41804
rect 31612 40226 31668 40236
rect 32396 40460 33124 40516
rect 32284 40068 32340 40078
rect 32396 40068 32452 40460
rect 32284 40066 32452 40068
rect 32284 40014 32286 40066
rect 32338 40014 32452 40066
rect 32284 40012 32452 40014
rect 32508 40292 32564 40302
rect 32284 40002 32340 40012
rect 32508 38946 32564 40236
rect 33068 40292 33124 40302
rect 33068 39954 33124 40236
rect 33964 40068 34020 41804
rect 34076 41858 34132 41870
rect 34076 41806 34078 41858
rect 34130 41806 34132 41858
rect 34076 40404 34132 41806
rect 34412 40962 34468 40974
rect 34412 40910 34414 40962
rect 34466 40910 34468 40962
rect 34412 40740 34468 40910
rect 34748 40962 34804 42252
rect 35084 41972 35140 43484
rect 35196 43372 35460 43382
rect 35252 43316 35300 43372
rect 35356 43316 35404 43372
rect 35196 43306 35460 43316
rect 35868 42978 35924 43652
rect 35868 42926 35870 42978
rect 35922 42926 35924 42978
rect 35868 42914 35924 42926
rect 37100 42978 37156 43708
rect 37100 42926 37102 42978
rect 37154 42926 37156 42978
rect 37100 42914 37156 42926
rect 35308 42756 35364 42766
rect 35308 42662 35364 42700
rect 35196 41972 35252 41982
rect 35084 41970 35252 41972
rect 35084 41918 35198 41970
rect 35250 41918 35252 41970
rect 35084 41916 35252 41918
rect 35196 41906 35252 41916
rect 35868 41970 35924 41982
rect 35868 41918 35870 41970
rect 35922 41918 35924 41970
rect 35196 41356 35460 41366
rect 35252 41300 35300 41356
rect 35356 41300 35404 41356
rect 35196 41290 35460 41300
rect 34748 40910 34750 40962
rect 34802 40910 34804 40962
rect 34748 40898 34804 40910
rect 34972 41188 35028 41198
rect 34412 40674 34468 40684
rect 34076 40338 34132 40348
rect 34076 40068 34132 40078
rect 33964 40066 34132 40068
rect 33964 40014 34078 40066
rect 34130 40014 34132 40066
rect 33964 40012 34132 40014
rect 34076 40002 34132 40012
rect 33068 39902 33070 39954
rect 33122 39902 33124 39954
rect 33068 39890 33124 39902
rect 34972 39954 35028 41132
rect 35868 40962 35924 41918
rect 35868 40910 35870 40962
rect 35922 40910 35924 40962
rect 35868 40898 35924 40910
rect 36764 41746 36820 41758
rect 36764 41694 36766 41746
rect 36818 41694 36820 41746
rect 36764 40740 36820 41694
rect 37100 41748 37156 41758
rect 37212 41748 37268 44604
rect 38332 44100 38388 44718
rect 37884 44044 38388 44100
rect 38780 44996 38836 45836
rect 38780 44100 38836 44940
rect 38892 44660 38948 46510
rect 39004 45444 39060 46844
rect 39900 46676 39956 46686
rect 39900 46562 39956 46620
rect 39900 46510 39902 46562
rect 39954 46510 39956 46562
rect 39900 46498 39956 46510
rect 40124 46228 40180 48638
rect 40348 48132 40404 48972
rect 41244 48916 41300 48926
rect 40796 48804 40852 48814
rect 40796 48710 40852 48748
rect 41244 48802 41300 48860
rect 41244 48750 41246 48802
rect 41298 48750 41300 48802
rect 40236 48076 40404 48132
rect 40236 46900 40292 48076
rect 40348 47908 40404 47918
rect 40796 47908 40852 47918
rect 40348 47906 40852 47908
rect 40348 47854 40350 47906
rect 40402 47854 40798 47906
rect 40850 47854 40852 47906
rect 40348 47852 40852 47854
rect 40348 47842 40404 47852
rect 40796 47842 40852 47852
rect 40236 46806 40292 46844
rect 40684 46898 40740 46910
rect 40684 46846 40686 46898
rect 40738 46846 40740 46898
rect 40684 46676 40740 46846
rect 40684 46610 40740 46620
rect 41132 46900 41188 46910
rect 40124 46162 40180 46172
rect 40908 46228 40964 46238
rect 40012 45668 40068 45678
rect 40012 45666 40180 45668
rect 40012 45614 40014 45666
rect 40066 45614 40180 45666
rect 40012 45612 40180 45614
rect 40012 45602 40068 45612
rect 39004 45378 39060 45388
rect 38892 44658 39060 44660
rect 38892 44606 38894 44658
rect 38946 44606 39060 44658
rect 38892 44604 39060 44606
rect 38892 44594 38948 44604
rect 38892 44100 38948 44110
rect 38780 44098 38948 44100
rect 38780 44046 38894 44098
rect 38946 44046 38948 44098
rect 38780 44044 38948 44046
rect 37884 42978 37940 44044
rect 37884 42926 37886 42978
rect 37938 42926 37940 42978
rect 37884 42914 37940 42926
rect 37996 43876 38052 43886
rect 37996 41972 38052 43820
rect 38332 42084 38388 44044
rect 38332 42028 38724 42084
rect 37884 41970 38052 41972
rect 37884 41918 37998 41970
rect 38050 41918 38052 41970
rect 37884 41916 38052 41918
rect 37100 41746 37268 41748
rect 37100 41694 37102 41746
rect 37154 41694 37268 41746
rect 37100 41692 37268 41694
rect 37436 41860 37492 41870
rect 37100 40964 37156 41692
rect 37324 40964 37380 40974
rect 37100 40908 37324 40964
rect 36764 40674 36820 40684
rect 37324 40850 37380 40908
rect 37324 40798 37326 40850
rect 37378 40798 37380 40850
rect 37100 40626 37156 40638
rect 37100 40574 37102 40626
rect 37154 40574 37156 40626
rect 37100 40516 37156 40574
rect 37100 40450 37156 40460
rect 34972 39902 34974 39954
rect 35026 39902 35028 39954
rect 34972 39890 35028 39902
rect 35532 39954 35588 39966
rect 35532 39902 35534 39954
rect 35586 39902 35588 39954
rect 35532 39844 35588 39902
rect 35532 39778 35588 39788
rect 36428 39842 36484 39854
rect 36428 39790 36430 39842
rect 36482 39790 36484 39842
rect 35644 39730 35700 39742
rect 35644 39678 35646 39730
rect 35698 39678 35700 39730
rect 35644 39620 35700 39678
rect 36428 39732 36484 39790
rect 35644 39554 35700 39564
rect 36092 39618 36148 39630
rect 36092 39566 36094 39618
rect 36146 39566 36148 39618
rect 34524 39506 34580 39518
rect 34524 39454 34526 39506
rect 34578 39454 34580 39506
rect 32508 38894 32510 38946
rect 32562 38894 32564 38946
rect 32508 37716 32564 38894
rect 33628 38948 33684 38958
rect 33628 38834 33684 38892
rect 34412 38948 34468 38958
rect 34412 38854 34468 38892
rect 33628 38782 33630 38834
rect 33682 38782 33684 38834
rect 33628 38770 33684 38782
rect 33180 38722 33236 38734
rect 33180 38670 33182 38722
rect 33234 38670 33236 38722
rect 33180 38668 33236 38670
rect 33068 38612 33236 38668
rect 33740 38722 33796 38734
rect 33740 38670 33742 38722
rect 33794 38670 33796 38722
rect 32732 38500 32788 38510
rect 32508 36818 32564 37660
rect 32508 36766 32510 36818
rect 32562 36766 32564 36818
rect 32172 36596 32228 36606
rect 32508 36596 32564 36766
rect 32172 36594 32564 36596
rect 32172 36542 32174 36594
rect 32226 36542 32564 36594
rect 32172 36540 32564 36542
rect 32172 36530 32228 36540
rect 32172 35812 32228 35822
rect 32172 35718 32228 35756
rect 32060 34804 32116 34814
rect 32116 34748 32340 34804
rect 32060 34710 32116 34748
rect 32060 33796 32116 33806
rect 32060 33684 32116 33740
rect 31836 33682 32116 33684
rect 31836 33630 32062 33682
rect 32114 33630 32116 33682
rect 31836 33628 32116 33630
rect 31500 33572 31556 33582
rect 31500 33570 31780 33572
rect 31500 33518 31502 33570
rect 31554 33518 31780 33570
rect 31500 33516 31780 33518
rect 31500 33506 31556 33516
rect 31612 32900 31668 32910
rect 31276 31892 31332 31902
rect 31164 31890 31332 31892
rect 31164 31838 31278 31890
rect 31330 31838 31332 31890
rect 31164 31836 31332 31838
rect 30828 31668 30884 31678
rect 30940 31668 30996 31836
rect 31276 31826 31332 31836
rect 31612 31780 31668 32844
rect 30828 31666 30996 31668
rect 30828 31614 30830 31666
rect 30882 31614 30996 31666
rect 30828 31612 30996 31614
rect 30828 31602 30884 31612
rect 28588 30370 28644 30380
rect 29148 30660 29204 30670
rect 29036 30324 29092 30334
rect 28140 30100 28196 30110
rect 28140 30006 28196 30044
rect 27804 29988 27860 29998
rect 27468 29822 27470 29874
rect 27522 29822 27524 29874
rect 27468 29810 27524 29822
rect 27692 29986 27860 29988
rect 27692 29934 27806 29986
rect 27858 29934 27860 29986
rect 27692 29932 27860 29934
rect 27692 29764 27748 29932
rect 27804 29922 27860 29932
rect 27020 29474 27076 29484
rect 27468 29652 27524 29662
rect 26908 28914 26964 28924
rect 27132 29090 27188 29102
rect 27132 29038 27134 29090
rect 27186 29038 27188 29090
rect 27132 28642 27188 29038
rect 27132 28590 27134 28642
rect 27186 28590 27188 28642
rect 27132 28578 27188 28590
rect 26796 28478 26798 28530
rect 26850 28478 26852 28530
rect 26796 28466 26852 28478
rect 27020 28420 27076 28430
rect 26908 28364 27020 28420
rect 26684 28252 26852 28308
rect 26684 27972 26740 27982
rect 26572 27970 26740 27972
rect 26572 27918 26686 27970
rect 26738 27918 26740 27970
rect 26572 27916 26740 27918
rect 26348 27748 26404 27758
rect 26348 27654 26404 27692
rect 25900 26516 25956 26526
rect 25564 26450 25620 26460
rect 25788 26514 25956 26516
rect 25788 26462 25902 26514
rect 25954 26462 25956 26514
rect 25788 26460 25956 26462
rect 25340 25442 25396 25452
rect 25564 25842 25620 25854
rect 25564 25790 25566 25842
rect 25618 25790 25620 25842
rect 25564 25620 25620 25790
rect 24892 25006 24894 25058
rect 24946 25006 24948 25058
rect 24892 24994 24948 25006
rect 25228 25396 25284 25406
rect 25228 23940 25284 25340
rect 25452 24724 25508 24734
rect 25340 24612 25396 24622
rect 25340 24518 25396 24556
rect 25116 23884 25284 23940
rect 25116 23548 25172 23884
rect 25452 23826 25508 24668
rect 25564 24722 25620 25564
rect 25788 25284 25844 26460
rect 25900 26450 25956 26460
rect 26012 25954 26068 26908
rect 26124 26852 26292 26908
rect 26348 27076 26404 27086
rect 26348 26908 26404 27020
rect 26572 26908 26628 27916
rect 26684 27906 26740 27916
rect 26348 26852 26628 26908
rect 26124 26850 26180 26852
rect 26124 26798 26126 26850
rect 26178 26798 26180 26850
rect 26124 26786 26180 26798
rect 26348 26626 26404 26852
rect 26572 26740 26628 26750
rect 26348 26574 26350 26626
rect 26402 26574 26404 26626
rect 26348 26562 26404 26574
rect 26460 26738 26628 26740
rect 26460 26686 26574 26738
rect 26626 26686 26628 26738
rect 26460 26684 26628 26686
rect 26460 26068 26516 26684
rect 26572 26674 26628 26684
rect 26796 26628 26852 28252
rect 26908 26852 26964 28364
rect 27020 28354 27076 28364
rect 27468 27972 27524 29596
rect 27692 29090 27748 29708
rect 28476 29762 28532 29774
rect 28476 29710 28478 29762
rect 28530 29710 28532 29762
rect 28476 29652 28532 29710
rect 28476 29586 28532 29596
rect 28924 29652 28980 29662
rect 28924 29558 28980 29596
rect 29036 29428 29092 30268
rect 29036 29362 29092 29372
rect 27692 29038 27694 29090
rect 27746 29038 27748 29090
rect 27692 29026 27748 29038
rect 27020 27970 27524 27972
rect 27020 27918 27470 27970
rect 27522 27918 27524 27970
rect 27020 27916 27524 27918
rect 27020 27858 27076 27916
rect 27468 27906 27524 27916
rect 27580 28868 27636 28878
rect 27020 27806 27022 27858
rect 27074 27806 27076 27858
rect 27020 27794 27076 27806
rect 27580 26908 27636 28812
rect 29148 28756 29204 30604
rect 29260 30546 29316 30558
rect 29260 30494 29262 30546
rect 29314 30494 29316 30546
rect 29260 30436 29316 30494
rect 29260 30370 29316 30380
rect 29708 30546 29764 30716
rect 29708 30494 29710 30546
rect 29762 30494 29764 30546
rect 29596 30212 29652 30222
rect 29596 29874 29652 30156
rect 29596 29822 29598 29874
rect 29650 29822 29652 29874
rect 29596 29810 29652 29822
rect 29260 29764 29316 29774
rect 29316 29708 29540 29764
rect 29260 29670 29316 29708
rect 29148 28690 29204 28700
rect 29484 28868 29540 29708
rect 29484 28754 29540 28812
rect 29484 28702 29486 28754
rect 29538 28702 29540 28754
rect 29484 28690 29540 28702
rect 29596 29650 29652 29662
rect 29596 29598 29598 29650
rect 29650 29598 29652 29650
rect 29596 27972 29652 29598
rect 29708 29428 29764 30494
rect 30492 30770 30772 30772
rect 30492 30718 30718 30770
rect 30770 30718 30772 30770
rect 30492 30716 30772 30718
rect 30156 29988 30212 29998
rect 30044 29986 30212 29988
rect 30044 29934 30158 29986
rect 30210 29934 30212 29986
rect 30044 29932 30212 29934
rect 29932 29764 29988 29774
rect 29932 29670 29988 29708
rect 29708 29372 29988 29428
rect 29820 29204 29876 29214
rect 29708 28754 29764 28766
rect 29708 28702 29710 28754
rect 29762 28702 29764 28754
rect 29708 28196 29764 28702
rect 29820 28642 29876 29148
rect 29820 28590 29822 28642
rect 29874 28590 29876 28642
rect 29820 28578 29876 28590
rect 29708 28140 29876 28196
rect 29708 27972 29764 27982
rect 29596 27970 29764 27972
rect 29596 27918 29710 27970
rect 29762 27918 29764 27970
rect 29596 27916 29764 27918
rect 29708 27906 29764 27916
rect 29820 27972 29876 28140
rect 29820 27906 29876 27916
rect 29596 27746 29652 27758
rect 29596 27694 29598 27746
rect 29650 27694 29652 27746
rect 29596 26964 29652 27694
rect 29820 27746 29876 27758
rect 29820 27694 29822 27746
rect 29874 27694 29876 27746
rect 27020 26852 27076 26862
rect 27580 26852 27860 26908
rect 29596 26898 29652 26908
rect 29708 27636 29764 27646
rect 26908 26850 27076 26852
rect 26908 26798 27022 26850
rect 27074 26798 27076 26850
rect 26908 26796 27076 26798
rect 27020 26786 27076 26796
rect 26796 26572 27076 26628
rect 26236 26012 26516 26068
rect 26908 26068 26964 26078
rect 26012 25902 26014 25954
rect 26066 25902 26068 25954
rect 26012 25890 26068 25902
rect 26124 25956 26180 25966
rect 26124 25842 26180 25900
rect 26124 25790 26126 25842
rect 26178 25790 26180 25842
rect 26124 25778 26180 25790
rect 25900 25732 25956 25742
rect 25900 25638 25956 25676
rect 25788 25218 25844 25228
rect 26124 24724 26180 24734
rect 25564 24670 25566 24722
rect 25618 24670 25620 24722
rect 25564 24658 25620 24670
rect 25900 24668 26124 24724
rect 25788 24610 25844 24622
rect 25788 24558 25790 24610
rect 25842 24558 25844 24610
rect 25452 23774 25454 23826
rect 25506 23774 25508 23826
rect 25452 23762 25508 23774
rect 25676 24500 25732 24510
rect 25228 23716 25284 23726
rect 25284 23660 25396 23716
rect 25228 23650 25284 23660
rect 25116 23492 25284 23548
rect 25116 22596 25172 22606
rect 25116 21698 25172 22540
rect 25116 21646 25118 21698
rect 25170 21646 25172 21698
rect 25116 21252 25172 21646
rect 25116 21186 25172 21196
rect 24780 20132 25172 20188
rect 24108 19854 24110 19906
rect 24162 19854 24164 19906
rect 24108 19842 24164 19854
rect 24556 19572 24612 19582
rect 24556 19478 24612 19516
rect 24444 18564 24500 18574
rect 25004 18564 25060 18574
rect 23996 18562 24500 18564
rect 23996 18510 24446 18562
rect 24498 18510 24500 18562
rect 23996 18508 24500 18510
rect 23548 17826 23604 17836
rect 24444 17892 24500 18508
rect 24444 17826 24500 17836
rect 24556 18562 25060 18564
rect 24556 18510 25006 18562
rect 25058 18510 25060 18562
rect 24556 18508 25060 18510
rect 24220 17554 24276 17566
rect 24220 17502 24222 17554
rect 24274 17502 24276 17554
rect 23772 16772 23828 16782
rect 22204 16658 22708 16660
rect 22204 16606 22206 16658
rect 22258 16606 22708 16658
rect 22204 16604 22708 16606
rect 22204 16594 22260 16604
rect 22652 15876 22708 16604
rect 23772 16658 23828 16716
rect 23772 16606 23774 16658
rect 23826 16606 23828 16658
rect 23772 16594 23828 16606
rect 23436 16548 23492 16558
rect 23100 16546 23492 16548
rect 23100 16494 23438 16546
rect 23490 16494 23492 16546
rect 23100 16492 23492 16494
rect 22428 15874 22708 15876
rect 22428 15822 22654 15874
rect 22706 15822 22708 15874
rect 22428 15820 22708 15822
rect 22428 14756 22484 15820
rect 22652 15810 22708 15820
rect 22988 16436 23044 16446
rect 22988 15876 23044 16380
rect 22988 15810 23044 15820
rect 22988 15652 23044 15662
rect 22988 15558 23044 15596
rect 23100 15316 23156 16492
rect 23436 16482 23492 16492
rect 24108 16546 24164 16558
rect 24108 16494 24110 16546
rect 24162 16494 24164 16546
rect 24108 15874 24164 16494
rect 24108 15822 24110 15874
rect 24162 15822 24164 15874
rect 24108 15810 24164 15822
rect 24220 15876 24276 17502
rect 24444 16660 24500 16670
rect 24556 16660 24612 18508
rect 25004 18498 25060 18508
rect 24444 16658 24612 16660
rect 24444 16606 24446 16658
rect 24498 16606 24612 16658
rect 24444 16604 24612 16606
rect 24668 17554 24724 17566
rect 24668 17502 24670 17554
rect 24722 17502 24724 17554
rect 24444 16594 24500 16604
rect 23884 15764 23940 15774
rect 22428 14644 22484 14700
rect 22652 15260 23156 15316
rect 23436 15650 23492 15662
rect 23436 15598 23438 15650
rect 23490 15598 23492 15650
rect 22652 14754 22708 15260
rect 22652 14702 22654 14754
rect 22706 14702 22708 14754
rect 22652 14690 22708 14702
rect 22428 14642 22596 14644
rect 22428 14590 22430 14642
rect 22482 14590 22596 14642
rect 22428 14588 22596 14590
rect 21980 13918 21982 13970
rect 22034 13918 22036 13970
rect 21980 13906 22036 13918
rect 22092 14530 22148 14542
rect 22092 14478 22094 14530
rect 22146 14478 22148 14530
rect 20972 13858 21364 13860
rect 20972 13806 20974 13858
rect 21026 13806 21364 13858
rect 20972 13804 21364 13806
rect 20972 13794 21028 13804
rect 21308 12740 21364 13804
rect 21420 13766 21476 13804
rect 21644 13748 21700 13758
rect 21420 12740 21476 12750
rect 21308 12738 21476 12740
rect 21308 12686 21422 12738
rect 21474 12686 21476 12738
rect 21308 12684 21476 12686
rect 21308 12292 21364 12684
rect 21420 12674 21476 12684
rect 21308 12226 21364 12236
rect 21084 11506 21140 11518
rect 21084 11454 21086 11506
rect 21138 11454 21140 11506
rect 21084 10612 21140 11454
rect 21084 10546 21140 10556
rect 21644 10612 21700 13692
rect 22092 12852 22148 14478
rect 22316 14308 22372 14318
rect 22316 13748 22372 14252
rect 22316 13654 22372 13692
rect 21868 12796 22148 12852
rect 21868 12738 21924 12796
rect 21868 12686 21870 12738
rect 21922 12686 21924 12738
rect 21868 12674 21924 12686
rect 22092 11954 22148 12796
rect 22092 11902 22094 11954
rect 22146 11902 22148 11954
rect 22092 11890 22148 11902
rect 22428 11730 22484 14588
rect 22540 14532 22596 14588
rect 22540 14476 22820 14532
rect 22764 13858 22820 14476
rect 22764 13806 22766 13858
rect 22818 13806 22820 13858
rect 22764 13794 22820 13806
rect 23212 13860 23268 13870
rect 23436 13860 23492 15598
rect 23884 15650 23940 15708
rect 23884 15598 23886 15650
rect 23938 15598 23940 15650
rect 23884 15586 23940 15598
rect 24220 14756 24276 15820
rect 24668 15764 24724 17502
rect 25004 16772 25060 16782
rect 25004 16658 25060 16716
rect 25004 16606 25006 16658
rect 25058 16606 25060 16658
rect 25004 16594 25060 16606
rect 24668 15698 24724 15708
rect 23996 14700 24276 14756
rect 24332 15652 24388 15662
rect 23996 14530 24052 14700
rect 23996 14478 23998 14530
rect 24050 14478 24052 14530
rect 23996 14466 24052 14478
rect 23268 13804 23492 13860
rect 24220 13860 24276 13870
rect 23212 13766 23268 13804
rect 23324 12738 23380 13804
rect 24220 13766 24276 13804
rect 23324 12686 23326 12738
rect 23378 12686 23380 12738
rect 22876 11956 22932 11966
rect 22876 11844 22932 11900
rect 22428 11678 22430 11730
rect 22482 11678 22484 11730
rect 22428 11666 22484 11678
rect 22764 11842 22932 11844
rect 22764 11790 22878 11842
rect 22930 11790 22932 11842
rect 22764 11788 22932 11790
rect 22316 11620 22372 11630
rect 21980 11506 22036 11518
rect 21980 11454 21982 11506
rect 22034 11454 22036 11506
rect 21980 11396 22036 11454
rect 21980 10836 22036 11340
rect 21980 10770 22036 10780
rect 21980 10612 22036 10622
rect 21644 10610 21812 10612
rect 21644 10558 21646 10610
rect 21698 10558 21812 10610
rect 21644 10556 21812 10558
rect 21644 10546 21700 10556
rect 21308 10500 21364 10510
rect 21308 10406 21364 10444
rect 20860 8642 20916 8652
rect 21308 8930 21364 8942
rect 21308 8878 21310 8930
rect 21362 8878 21364 8930
rect 19852 8484 19908 8494
rect 19740 8428 19852 8484
rect 19852 8418 19908 8428
rect 19836 8092 20100 8102
rect 19892 8036 19940 8092
rect 19996 8036 20044 8092
rect 19836 8026 20100 8036
rect 20188 7924 20244 8540
rect 20748 8596 20804 8606
rect 20076 7868 20244 7924
rect 20636 8484 20692 8494
rect 19516 7534 19518 7586
rect 19570 7534 19572 7586
rect 19516 7522 19572 7534
rect 19964 7588 20020 7598
rect 20076 7588 20132 7868
rect 19964 7586 20132 7588
rect 19964 7534 19966 7586
rect 20018 7534 20132 7586
rect 19964 7532 20132 7534
rect 19964 7522 20020 7532
rect 20076 6804 20132 7532
rect 20636 7586 20692 8428
rect 20748 8482 20804 8540
rect 20748 8430 20750 8482
rect 20802 8430 20804 8482
rect 20748 8418 20804 8430
rect 21308 8428 21364 8878
rect 21532 8708 21588 8718
rect 21308 8372 21476 8428
rect 20636 7534 20638 7586
rect 20690 7534 20692 7586
rect 20076 6748 20244 6804
rect 20188 6692 20244 6748
rect 20412 6692 20468 6702
rect 20188 6636 20412 6692
rect 19404 6514 19460 6524
rect 20076 6580 20132 6590
rect 20132 6524 20244 6580
rect 20076 6514 20132 6524
rect 4620 6302 4622 6354
rect 4674 6302 4676 6354
rect 4620 6290 4676 6302
rect 18172 6356 18228 6366
rect 18172 6262 18228 6300
rect 19836 6076 20100 6086
rect 19892 6020 19940 6076
rect 19996 6020 20044 6076
rect 19836 6010 20100 6020
rect 20076 5796 20132 5806
rect 20188 5796 20244 6524
rect 20076 5794 20244 5796
rect 20076 5742 20078 5794
rect 20130 5742 20244 5794
rect 20076 5740 20244 5742
rect 20412 5796 20468 6636
rect 20636 6468 20692 7534
rect 21196 6580 21252 6590
rect 21196 6486 21252 6524
rect 20524 6356 20580 6366
rect 20524 6262 20580 6300
rect 20524 5796 20580 5806
rect 20412 5794 20580 5796
rect 20412 5742 20526 5794
rect 20578 5742 20580 5794
rect 20412 5740 20580 5742
rect 20636 5796 20692 6412
rect 20972 5796 21028 5806
rect 20636 5794 21028 5796
rect 20636 5742 20974 5794
rect 21026 5742 21028 5794
rect 20636 5740 21028 5742
rect 20076 5730 20132 5740
rect 20524 5730 20580 5740
rect 20972 5730 21028 5740
rect 21420 5684 21476 8372
rect 21532 7588 21588 8652
rect 21756 8428 21812 10556
rect 21980 10518 22036 10556
rect 22316 10610 22372 11564
rect 22316 10558 22318 10610
rect 22370 10558 22372 10610
rect 22316 10546 22372 10558
rect 22428 10388 22484 10398
rect 22428 9938 22484 10332
rect 22428 9886 22430 9938
rect 22482 9886 22484 9938
rect 22428 9874 22484 9886
rect 22764 8706 22820 11788
rect 22876 11778 22932 11788
rect 23100 11732 23156 11742
rect 23100 11638 23156 11676
rect 23324 11396 23380 12686
rect 24220 12740 24276 12750
rect 24332 12740 24388 15596
rect 24668 14644 24724 14654
rect 24444 14532 24500 14542
rect 24444 13860 24500 14476
rect 24444 13794 24500 13804
rect 24668 13858 24724 14588
rect 24668 13806 24670 13858
rect 24722 13806 24724 13858
rect 24668 13794 24724 13806
rect 24220 12738 24388 12740
rect 24220 12686 24222 12738
rect 24274 12686 24388 12738
rect 24220 12684 24388 12686
rect 23772 12404 23828 12414
rect 24220 12404 24276 12684
rect 23772 12402 24276 12404
rect 23772 12350 23774 12402
rect 23826 12350 24276 12402
rect 23772 12348 24276 12350
rect 24332 12514 24388 12526
rect 24332 12462 24334 12514
rect 24386 12462 24388 12514
rect 23548 11620 23604 11630
rect 23548 11526 23604 11564
rect 23212 11340 23324 11396
rect 22764 8654 22766 8706
rect 22818 8654 22820 8706
rect 22204 8484 22260 8522
rect 22764 8428 22820 8654
rect 21756 8372 21924 8428
rect 22204 8372 22820 8428
rect 22876 10498 22932 10510
rect 22876 10446 22878 10498
rect 22930 10446 22932 10498
rect 22876 10164 22932 10446
rect 21532 6578 21588 7532
rect 21532 6526 21534 6578
rect 21586 6526 21588 6578
rect 21532 6514 21588 6526
rect 21532 5684 21588 5694
rect 21420 5682 21588 5684
rect 21420 5630 21534 5682
rect 21586 5630 21588 5682
rect 21420 5628 21588 5630
rect 21532 5618 21588 5628
rect 21868 5682 21924 8372
rect 22540 7700 22596 7710
rect 21980 6692 22036 6702
rect 21980 6578 22036 6636
rect 21980 6526 21982 6578
rect 22034 6526 22036 6578
rect 21980 6514 22036 6526
rect 21868 5630 21870 5682
rect 21922 5630 21924 5682
rect 21868 5618 21924 5630
rect 22204 6356 22260 6366
rect 22204 5682 22260 6300
rect 22540 5794 22596 7644
rect 22652 6578 22708 8372
rect 22652 6526 22654 6578
rect 22706 6526 22708 6578
rect 22652 6514 22708 6526
rect 22540 5742 22542 5794
rect 22594 5742 22596 5794
rect 22540 5730 22596 5742
rect 22204 5630 22206 5682
rect 22258 5630 22260 5682
rect 22204 5618 22260 5630
rect 22876 5684 22932 10108
rect 23212 9938 23268 11340
rect 23324 11330 23380 11340
rect 23436 11508 23492 11518
rect 23436 10610 23492 11452
rect 23436 10558 23438 10610
rect 23490 10558 23492 10610
rect 23436 10546 23492 10558
rect 23212 9886 23214 9938
rect 23266 9886 23268 9938
rect 23212 9828 23268 9886
rect 23212 9826 23380 9828
rect 23212 9774 23214 9826
rect 23266 9774 23380 9826
rect 23212 9772 23380 9774
rect 23212 9762 23268 9772
rect 23324 8708 23380 9772
rect 23660 9492 23716 9502
rect 23772 9492 23828 12348
rect 24332 11956 24388 12462
rect 24332 11890 24388 11900
rect 25004 11956 25060 11966
rect 23660 9490 23828 9492
rect 23660 9438 23662 9490
rect 23714 9438 23828 9490
rect 23660 9436 23828 9438
rect 23996 11730 24052 11742
rect 23996 11678 23998 11730
rect 24050 11678 24052 11730
rect 23660 9378 23716 9436
rect 23660 9326 23662 9378
rect 23714 9326 23716 9378
rect 23660 9314 23716 9326
rect 23884 8820 23940 8830
rect 23324 8706 23716 8708
rect 23324 8654 23326 8706
rect 23378 8654 23716 8706
rect 23324 8652 23716 8654
rect 23324 8642 23380 8652
rect 23660 8596 23716 8652
rect 23660 8502 23716 8540
rect 23884 8594 23940 8764
rect 23884 8542 23886 8594
rect 23938 8542 23940 8594
rect 23884 8530 23940 8542
rect 23996 7700 24052 11678
rect 24220 11620 24276 11630
rect 24220 11526 24276 11564
rect 25004 11508 25060 11900
rect 25116 11732 25172 20132
rect 25228 18900 25284 23492
rect 25340 21810 25396 23660
rect 25676 22706 25732 24444
rect 25788 24052 25844 24558
rect 25788 23986 25844 23996
rect 25788 23828 25844 23838
rect 25788 23734 25844 23772
rect 25788 23604 25844 23614
rect 25788 22820 25844 23548
rect 25900 23042 25956 24668
rect 26124 24658 26180 24668
rect 25900 22990 25902 23042
rect 25954 22990 25956 23042
rect 25900 22978 25956 22990
rect 25788 22764 26180 22820
rect 25676 22654 25678 22706
rect 25730 22654 25732 22706
rect 25564 22596 25620 22606
rect 25564 22502 25620 22540
rect 25340 21758 25342 21810
rect 25394 21758 25396 21810
rect 25340 21746 25396 21758
rect 25676 21812 25732 22654
rect 26124 22034 26180 22764
rect 26124 21982 26126 22034
rect 26178 21982 26180 22034
rect 26124 21970 26180 21982
rect 25676 21718 25732 21756
rect 25452 21588 25508 21598
rect 25452 20466 25508 21532
rect 26236 21028 26292 26012
rect 26572 25956 26628 25966
rect 26460 25900 26572 25956
rect 26348 25730 26404 25742
rect 26348 25678 26350 25730
rect 26402 25678 26404 25730
rect 26348 25396 26404 25678
rect 26348 25330 26404 25340
rect 26460 24948 26516 25900
rect 26572 25890 26628 25900
rect 26908 25954 26964 26012
rect 26908 25902 26910 25954
rect 26962 25902 26964 25954
rect 26908 25890 26964 25902
rect 26684 25844 26740 25854
rect 27020 25844 27076 26572
rect 26740 25788 26852 25844
rect 26684 25778 26740 25788
rect 26796 25730 26852 25788
rect 27020 25750 27076 25788
rect 27356 26516 27412 26526
rect 26796 25678 26798 25730
rect 26850 25678 26852 25730
rect 26796 25666 26852 25678
rect 27244 25730 27300 25742
rect 27244 25678 27246 25730
rect 27298 25678 27300 25730
rect 26572 25620 26628 25630
rect 26628 25564 26740 25620
rect 26572 25554 26628 25564
rect 26460 24892 26628 24948
rect 26460 24724 26516 24734
rect 26460 24630 26516 24668
rect 26572 24612 26628 24892
rect 26684 24836 26740 25564
rect 26908 25396 26964 25406
rect 26796 25060 26852 25070
rect 26796 24966 26852 25004
rect 26684 24780 26852 24836
rect 26684 24612 26740 24622
rect 26572 24610 26740 24612
rect 26572 24558 26686 24610
rect 26738 24558 26740 24610
rect 26572 24556 26740 24558
rect 26684 24546 26740 24556
rect 26460 24500 26516 24510
rect 26348 24052 26404 24062
rect 26348 23958 26404 23996
rect 26460 23938 26516 24444
rect 26460 23886 26462 23938
rect 26514 23886 26516 23938
rect 26460 23874 26516 23886
rect 26684 23940 26740 23950
rect 26684 23714 26740 23884
rect 26684 23662 26686 23714
rect 26738 23662 26740 23714
rect 26684 23604 26740 23662
rect 26684 23538 26740 23548
rect 26348 23492 26404 23502
rect 26348 22706 26404 23436
rect 26348 22654 26350 22706
rect 26402 22654 26404 22706
rect 26348 22642 26404 22654
rect 26796 22932 26852 24780
rect 26908 24722 26964 25340
rect 27244 25396 27300 25678
rect 27244 25330 27300 25340
rect 26908 24670 26910 24722
rect 26962 24670 26964 24722
rect 26908 24658 26964 24670
rect 27244 23940 27300 23950
rect 27244 23846 27300 23884
rect 26796 22706 26852 22876
rect 26796 22654 26798 22706
rect 26850 22654 26852 22706
rect 26796 22642 26852 22654
rect 26908 22596 26964 22606
rect 26908 22502 26964 22540
rect 27356 22260 27412 26460
rect 27692 25620 27748 25630
rect 27580 25564 27692 25620
rect 27468 24612 27524 24622
rect 27468 24518 27524 24556
rect 27580 24500 27636 25564
rect 27692 25554 27748 25564
rect 27804 24612 27860 26852
rect 28588 26514 28644 26526
rect 28588 26462 28590 26514
rect 28642 26462 28644 26514
rect 27916 25956 27972 25966
rect 27916 24836 27972 25900
rect 28476 25956 28532 25966
rect 28588 25956 28644 26462
rect 29596 26514 29652 26526
rect 29596 26462 29598 26514
rect 29650 26462 29652 26514
rect 29484 26292 29540 26302
rect 28476 25954 28588 25956
rect 28476 25902 28478 25954
rect 28530 25902 28588 25954
rect 28476 25900 28588 25902
rect 28476 25890 28532 25900
rect 28588 25890 28644 25900
rect 29372 25956 29428 25966
rect 29372 25862 29428 25900
rect 28028 25620 28084 25630
rect 28028 25526 28084 25564
rect 28588 25620 28644 25630
rect 27916 24834 28084 24836
rect 27916 24782 27918 24834
rect 27970 24782 28084 24834
rect 27916 24780 28084 24782
rect 27916 24770 27972 24780
rect 27804 24556 27972 24612
rect 27580 24276 27636 24444
rect 27468 24220 27636 24276
rect 27692 24388 27748 24398
rect 27468 23940 27524 24220
rect 27468 23826 27524 23884
rect 27468 23774 27470 23826
rect 27522 23774 27524 23826
rect 27468 23762 27524 23774
rect 27580 23828 27636 23838
rect 27580 23734 27636 23772
rect 27468 22932 27524 22942
rect 27468 22482 27524 22876
rect 27468 22430 27470 22482
rect 27522 22430 27524 22482
rect 27468 22418 27524 22430
rect 27356 22204 27524 22260
rect 26236 20962 26292 20972
rect 26348 21812 26404 21822
rect 26348 20802 26404 21756
rect 27356 21812 27412 21822
rect 27356 21718 27412 21756
rect 26460 21700 26516 21710
rect 26460 21606 26516 21644
rect 26908 21586 26964 21598
rect 26908 21534 26910 21586
rect 26962 21534 26964 21586
rect 26348 20750 26350 20802
rect 26402 20750 26404 20802
rect 26348 20738 26404 20750
rect 26796 21252 26852 21262
rect 26796 20802 26852 21196
rect 26796 20750 26798 20802
rect 26850 20750 26852 20802
rect 26796 20738 26852 20750
rect 25452 20414 25454 20466
rect 25506 20414 25508 20466
rect 25452 20354 25508 20414
rect 25452 20302 25454 20354
rect 25506 20302 25508 20354
rect 25340 20244 25396 20254
rect 25340 19908 25396 20188
rect 25452 19908 25508 20302
rect 25900 20466 25956 20478
rect 25900 20414 25902 20466
rect 25954 20414 25956 20466
rect 25900 20354 25956 20414
rect 25900 20302 25902 20354
rect 25954 20302 25956 20354
rect 25900 20290 25956 20302
rect 26908 20354 26964 21534
rect 27132 20468 27188 20478
rect 27244 20468 27300 20478
rect 27132 20466 27244 20468
rect 27132 20414 27134 20466
rect 27186 20414 27244 20466
rect 27132 20412 27244 20414
rect 27132 20402 27188 20412
rect 27244 20374 27300 20412
rect 26908 20302 26910 20354
rect 26962 20302 26964 20354
rect 26908 20290 26964 20302
rect 27356 20354 27412 20366
rect 27356 20302 27358 20354
rect 27410 20302 27412 20354
rect 26012 19908 26068 19918
rect 25340 19906 25508 19908
rect 25340 19854 25342 19906
rect 25394 19854 25508 19906
rect 25340 19852 25508 19854
rect 25788 19852 26012 19908
rect 25340 19842 25396 19852
rect 25228 18834 25284 18844
rect 25676 18452 25732 18462
rect 25676 18358 25732 18396
rect 25788 17892 25844 19852
rect 26012 19814 26068 19852
rect 27356 19796 27412 20302
rect 26460 19572 26516 19582
rect 26908 19572 26964 19582
rect 26460 19570 26628 19572
rect 26460 19518 26462 19570
rect 26514 19518 26628 19570
rect 26460 19516 26628 19518
rect 26460 19506 26516 19516
rect 26348 18564 26404 18574
rect 26348 18562 26516 18564
rect 26348 18510 26350 18562
rect 26402 18510 26516 18562
rect 26348 18508 26516 18510
rect 26348 18498 26404 18508
rect 26348 17892 26404 17902
rect 25788 17890 26180 17892
rect 25788 17838 25790 17890
rect 25842 17838 26180 17890
rect 25788 17836 26180 17838
rect 25788 17826 25844 17836
rect 25340 17556 25396 17566
rect 25340 17462 25396 17500
rect 25564 16546 25620 16558
rect 25564 16494 25566 16546
rect 25618 16494 25620 16546
rect 25564 15986 25620 16494
rect 25564 15934 25566 15986
rect 25618 15934 25620 15986
rect 25564 15922 25620 15934
rect 25340 15876 25396 15886
rect 25340 15762 25396 15820
rect 25340 15710 25342 15762
rect 25394 15710 25396 15762
rect 25340 13860 25396 15710
rect 25452 15762 25508 15774
rect 25452 15710 25454 15762
rect 25506 15710 25508 15762
rect 25452 14532 25508 15710
rect 25788 15764 25844 15774
rect 25844 15708 25956 15764
rect 25788 15670 25844 15708
rect 25452 14466 25508 14476
rect 25788 14420 25844 14430
rect 25452 13860 25508 13870
rect 25340 13804 25452 13860
rect 25452 13766 25508 13804
rect 25788 12626 25844 14364
rect 25900 13858 25956 15708
rect 26012 15652 26068 15662
rect 26012 15558 26068 15596
rect 26012 14644 26068 14654
rect 26124 14644 26180 17836
rect 26348 17798 26404 17836
rect 26460 17556 26516 18508
rect 26572 17780 26628 19516
rect 26684 18900 26740 18910
rect 26684 18806 26740 18844
rect 26908 18898 26964 19516
rect 26908 18846 26910 18898
rect 26962 18846 26964 18898
rect 26908 18834 26964 18846
rect 27244 18898 27300 18910
rect 27244 18846 27246 18898
rect 27298 18846 27300 18898
rect 27244 18786 27300 18846
rect 27244 18734 27246 18786
rect 27298 18734 27300 18786
rect 27244 18722 27300 18734
rect 26572 17714 26628 17724
rect 27356 17890 27412 19740
rect 27356 17838 27358 17890
rect 27410 17838 27412 17890
rect 26908 17556 26964 17566
rect 27356 17556 27412 17838
rect 26460 17554 27076 17556
rect 26460 17502 26910 17554
rect 26962 17502 27076 17554
rect 26460 17500 27076 17502
rect 26908 17462 26964 17500
rect 27020 17108 27076 17500
rect 27356 17490 27412 17500
rect 27020 17052 27412 17108
rect 27244 16772 27300 16782
rect 27244 16678 27300 16716
rect 26236 16436 26292 16446
rect 26236 16434 26516 16436
rect 26236 16382 26238 16434
rect 26290 16382 26516 16434
rect 26236 16380 26516 16382
rect 26236 16370 26292 16380
rect 26068 14588 26180 14644
rect 26012 14550 26068 14588
rect 26124 13970 26180 14588
rect 26236 14532 26292 14570
rect 26236 14466 26292 14476
rect 26348 14420 26404 14430
rect 26124 13918 26126 13970
rect 26178 13918 26180 13970
rect 26124 13906 26180 13918
rect 26236 14308 26292 14318
rect 25900 13806 25902 13858
rect 25954 13806 25956 13858
rect 25900 13794 25956 13806
rect 25788 12574 25790 12626
rect 25842 12574 25844 12626
rect 25788 12562 25844 12574
rect 25116 11666 25172 11676
rect 25340 11732 25396 11742
rect 25340 11638 25396 11676
rect 25004 10610 25060 11452
rect 25004 10558 25006 10610
rect 25058 10558 25060 10610
rect 24108 10388 24164 10398
rect 24108 10294 24164 10332
rect 24220 10052 24276 10062
rect 24220 9826 24276 9996
rect 24220 9774 24222 9826
rect 24274 9774 24276 9826
rect 24220 9762 24276 9774
rect 24668 9938 24724 9950
rect 24668 9886 24670 9938
rect 24722 9886 24724 9938
rect 24668 9826 24724 9886
rect 24668 9774 24670 9826
rect 24722 9774 24724 9826
rect 24668 9762 24724 9774
rect 24220 9378 24276 9390
rect 24220 9326 24222 9378
rect 24274 9326 24276 9378
rect 24220 8482 24276 9326
rect 24220 8430 24222 8482
rect 24274 8430 24276 8482
rect 24220 8428 24276 8430
rect 24668 8820 24724 8830
rect 24220 8372 24388 8428
rect 23996 7634 24052 7644
rect 22988 7588 23044 7598
rect 22988 7494 23044 7532
rect 23996 7364 24052 7374
rect 23660 7362 24052 7364
rect 23660 7310 23998 7362
rect 24050 7310 24052 7362
rect 23660 7308 24052 7310
rect 22988 5684 23044 5694
rect 22876 5682 23044 5684
rect 22876 5630 22990 5682
rect 23042 5630 23044 5682
rect 22876 5628 23044 5630
rect 22988 5618 23044 5628
rect 23660 5682 23716 7308
rect 23996 7298 24052 7308
rect 24332 6580 24388 8372
rect 24668 7924 24724 8764
rect 25004 8594 25060 10558
rect 25900 10722 25956 10734
rect 25900 10670 25902 10722
rect 25954 10670 25956 10722
rect 25340 10052 25396 10062
rect 25340 9828 25396 9996
rect 25228 9826 25396 9828
rect 25228 9774 25342 9826
rect 25394 9774 25396 9826
rect 25228 9772 25396 9774
rect 25004 8542 25006 8594
rect 25058 8542 25060 8594
rect 24892 7924 24948 7934
rect 24668 7868 24892 7924
rect 24668 7810 24724 7868
rect 24892 7858 24948 7868
rect 24668 7758 24670 7810
rect 24722 7758 24724 7810
rect 24668 7746 24724 7758
rect 25004 7588 25060 8542
rect 25004 7522 25060 7532
rect 25116 8596 25172 8606
rect 25116 7586 25172 8540
rect 25228 7698 25284 9772
rect 25340 9762 25396 9772
rect 25900 9714 25956 10670
rect 25900 9662 25902 9714
rect 25954 9662 25956 9714
rect 25900 9650 25956 9662
rect 26236 9714 26292 14252
rect 26348 13858 26404 14364
rect 26348 13806 26350 13858
rect 26402 13806 26404 13858
rect 26348 13794 26404 13806
rect 26460 12852 26516 16380
rect 26796 15540 26852 15550
rect 26684 15538 26852 15540
rect 26684 15486 26798 15538
rect 26850 15486 26852 15538
rect 26684 15484 26852 15486
rect 26572 14308 26628 14318
rect 26572 14214 26628 14252
rect 26684 13860 26740 15484
rect 26796 15474 26852 15484
rect 27020 15316 27076 15326
rect 26684 13794 26740 13804
rect 26796 14756 26852 14766
rect 26796 13860 26852 14700
rect 26908 14644 26964 14654
rect 26908 14550 26964 14588
rect 26796 13858 26908 13860
rect 26796 13806 26798 13858
rect 26850 13806 26908 13858
rect 26796 13794 26908 13806
rect 26852 13748 26908 13794
rect 26852 13692 26964 13748
rect 26908 12962 26964 13692
rect 27020 13636 27076 15260
rect 27244 13636 27300 13646
rect 27020 13634 27300 13636
rect 27020 13582 27246 13634
rect 27298 13582 27300 13634
rect 27020 13580 27300 13582
rect 26908 12910 26910 12962
rect 26962 12910 26964 12962
rect 26908 12898 26964 12910
rect 26572 12852 26628 12862
rect 26460 12850 26628 12852
rect 26460 12798 26574 12850
rect 26626 12798 26628 12850
rect 26460 12796 26628 12798
rect 26572 12786 26628 12796
rect 27132 11844 27188 11854
rect 26348 11508 26404 11518
rect 26348 11414 26404 11452
rect 27132 10610 27188 11788
rect 27244 11506 27300 13580
rect 27356 13412 27412 17052
rect 27468 15428 27524 22204
rect 27692 20802 27748 24332
rect 27692 20750 27694 20802
rect 27746 20750 27748 20802
rect 27692 20354 27748 20750
rect 27692 20302 27694 20354
rect 27746 20302 27748 20354
rect 27692 20290 27748 20302
rect 27804 22594 27860 22606
rect 27804 22542 27806 22594
rect 27858 22542 27860 22594
rect 27804 21588 27860 22542
rect 27804 20244 27860 21532
rect 27804 20178 27860 20188
rect 27580 19570 27636 19582
rect 27580 19518 27582 19570
rect 27634 19518 27636 19570
rect 27580 19012 27636 19518
rect 27692 19012 27748 19022
rect 27580 19010 27748 19012
rect 27580 18958 27694 19010
rect 27746 18958 27748 19010
rect 27580 18956 27748 18958
rect 27692 18786 27748 18956
rect 27692 18734 27694 18786
rect 27746 18734 27748 18786
rect 27692 18722 27748 18734
rect 27692 17556 27748 17566
rect 27468 15362 27524 15372
rect 27580 16546 27636 16558
rect 27580 16494 27582 16546
rect 27634 16494 27636 16546
rect 27580 16324 27636 16494
rect 27468 15204 27524 15214
rect 27468 14644 27524 15148
rect 27468 14578 27524 14588
rect 27356 13346 27412 13356
rect 27356 12962 27412 12974
rect 27580 12964 27636 16268
rect 27692 15204 27748 17500
rect 27692 15148 27860 15204
rect 27804 15092 27860 15148
rect 27692 14420 27748 14430
rect 27804 14420 27860 15036
rect 27748 14364 27860 14420
rect 27692 14306 27748 14364
rect 27692 14254 27694 14306
rect 27746 14254 27748 14306
rect 27692 14242 27748 14254
rect 27692 13970 27748 13982
rect 27692 13918 27694 13970
rect 27746 13918 27748 13970
rect 27692 13858 27748 13918
rect 27692 13806 27694 13858
rect 27746 13806 27748 13858
rect 27692 13794 27748 13806
rect 27356 12910 27358 12962
rect 27410 12910 27412 12962
rect 27356 12738 27412 12910
rect 27356 12686 27358 12738
rect 27410 12686 27412 12738
rect 27356 12674 27412 12686
rect 27468 12908 27636 12964
rect 27804 12962 27860 12974
rect 27804 12910 27806 12962
rect 27858 12910 27860 12962
rect 27244 11454 27246 11506
rect 27298 11454 27300 11506
rect 27244 11442 27300 11454
rect 27132 10558 27134 10610
rect 27186 10558 27188 10610
rect 27132 10546 27188 10558
rect 26908 10498 26964 10510
rect 26908 10446 26910 10498
rect 26962 10446 26964 10498
rect 26908 9826 26964 10446
rect 27356 10498 27412 10510
rect 27356 10446 27358 10498
rect 27410 10446 27412 10498
rect 26908 9774 26910 9826
rect 26962 9774 26964 9826
rect 26908 9762 26964 9774
rect 27020 10052 27076 10062
rect 26236 9662 26238 9714
rect 26290 9662 26292 9714
rect 26236 9650 26292 9662
rect 26572 9602 26628 9614
rect 26572 9550 26574 9602
rect 26626 9550 26628 9602
rect 26572 8428 26628 9550
rect 27020 8484 27076 9996
rect 27244 8596 27300 8606
rect 27244 8484 27300 8540
rect 26908 8482 27300 8484
rect 26908 8430 27246 8482
rect 27298 8430 27300 8482
rect 26908 8428 27300 8430
rect 25228 7646 25230 7698
rect 25282 7646 25284 7698
rect 25228 7634 25284 7646
rect 25676 8372 26628 8428
rect 26684 8372 26964 8428
rect 27244 8418 27300 8428
rect 25116 7534 25118 7586
rect 25170 7534 25172 7586
rect 25116 6692 25172 7534
rect 25116 6626 25172 6636
rect 25676 6690 25732 8372
rect 25676 6638 25678 6690
rect 25730 6638 25732 6690
rect 25676 6626 25732 6638
rect 25900 7586 25956 7598
rect 25900 7534 25902 7586
rect 25954 7534 25956 7586
rect 24332 6514 24388 6524
rect 24668 6580 24724 6590
rect 24332 6356 24388 6366
rect 24332 5794 24388 6300
rect 24332 5742 24334 5794
rect 24386 5742 24388 5794
rect 24332 5730 24388 5742
rect 23660 5630 23662 5682
rect 23714 5630 23716 5682
rect 23660 5618 23716 5630
rect 4476 5068 4740 5078
rect 4532 5012 4580 5068
rect 4636 5012 4684 5068
rect 4476 5002 4740 5012
rect 23996 4676 24052 4686
rect 23996 4582 24052 4620
rect 24668 4674 24724 6524
rect 25228 6580 25284 6590
rect 25228 5796 25284 6524
rect 25900 6580 25956 7534
rect 25900 6514 25956 6524
rect 26124 7588 26180 7598
rect 25340 6356 25396 6366
rect 25340 6262 25396 6300
rect 25340 5796 25396 5806
rect 25228 5794 25396 5796
rect 25228 5742 25342 5794
rect 25394 5742 25396 5794
rect 25228 5740 25396 5742
rect 25340 5730 25396 5740
rect 25900 5458 25956 5470
rect 25900 5406 25902 5458
rect 25954 5406 25956 5458
rect 24668 4622 24670 4674
rect 24722 4622 24724 4674
rect 24668 4610 24724 4622
rect 25452 5346 25508 5358
rect 25452 5294 25454 5346
rect 25506 5294 25508 5346
rect 25452 4676 25508 5294
rect 25452 4582 25508 4620
rect 25900 4676 25956 5406
rect 26124 5346 26180 7532
rect 26124 5294 26126 5346
rect 26178 5294 26180 5346
rect 26124 5282 26180 5294
rect 26348 5460 26404 5470
rect 26348 5346 26404 5404
rect 26348 5294 26350 5346
rect 26402 5294 26404 5346
rect 26348 5282 26404 5294
rect 25900 4610 25956 4620
rect 26684 4676 26740 8372
rect 27356 7812 27412 10446
rect 27468 10164 27524 12908
rect 27804 12738 27860 12910
rect 27804 12686 27806 12738
rect 27858 12686 27860 12738
rect 27804 12674 27860 12686
rect 27804 11844 27860 11854
rect 27804 11730 27860 11788
rect 27804 11678 27806 11730
rect 27858 11678 27860 11730
rect 27804 11666 27860 11678
rect 27804 10948 27860 10958
rect 27916 10948 27972 24556
rect 28028 23828 28084 24780
rect 28588 24834 28644 25564
rect 28588 24782 28590 24834
rect 28642 24782 28644 24834
rect 28588 24770 28644 24782
rect 28924 25618 28980 25630
rect 28924 25566 28926 25618
rect 28978 25566 28980 25618
rect 28924 24612 28980 25566
rect 29372 24722 29428 24734
rect 29372 24670 29374 24722
rect 29426 24670 29428 24722
rect 28924 24546 28980 24556
rect 29260 24612 29316 24622
rect 28028 23762 28084 23772
rect 29260 23716 29316 24556
rect 29372 24052 29428 24670
rect 29484 24276 29540 26236
rect 29596 25620 29652 26462
rect 29708 25842 29764 27580
rect 29708 25790 29710 25842
rect 29762 25790 29764 25842
rect 29708 25778 29764 25790
rect 29596 25554 29652 25564
rect 29820 24724 29876 27694
rect 29932 27412 29988 29372
rect 30044 29092 30100 29932
rect 30156 29922 30212 29932
rect 30492 29874 30548 30716
rect 30716 30706 30772 30716
rect 30828 30660 30884 30670
rect 30940 30660 30996 31612
rect 31388 31778 31668 31780
rect 31388 31726 31614 31778
rect 31666 31726 31668 31778
rect 31388 31724 31668 31726
rect 31164 30884 31220 30894
rect 31388 30884 31444 31724
rect 31612 31714 31668 31724
rect 31164 30882 31444 30884
rect 31164 30830 31166 30882
rect 31218 30830 31444 30882
rect 31164 30828 31444 30830
rect 31500 31554 31556 31566
rect 31500 31502 31502 31554
rect 31554 31502 31556 31554
rect 31164 30818 31220 30828
rect 30940 30604 31220 30660
rect 30828 30566 30884 30604
rect 31052 30436 31108 30446
rect 30492 29822 30494 29874
rect 30546 29822 30548 29874
rect 30492 29810 30548 29822
rect 30604 30434 31108 30436
rect 30604 30382 31054 30434
rect 31106 30382 31108 30434
rect 30604 30380 31108 30382
rect 30604 29092 30660 30380
rect 31052 30370 31108 30380
rect 31164 30212 31220 30604
rect 30044 27748 30100 29036
rect 30268 29036 30660 29092
rect 30940 30156 31220 30212
rect 31388 30658 31444 30670
rect 31388 30606 31390 30658
rect 31442 30606 31444 30658
rect 31388 30212 31444 30606
rect 30156 28756 30212 28766
rect 30156 28662 30212 28700
rect 30044 27746 30212 27748
rect 30044 27694 30046 27746
rect 30098 27694 30212 27746
rect 30044 27692 30212 27694
rect 30044 27682 30100 27692
rect 30156 27524 30212 27692
rect 30268 27746 30324 29036
rect 30716 28980 30772 28990
rect 30380 28868 30436 28878
rect 30380 28754 30436 28812
rect 30380 28702 30382 28754
rect 30434 28702 30436 28754
rect 30380 28690 30436 28702
rect 30604 28754 30660 28766
rect 30604 28702 30606 28754
rect 30658 28702 30660 28754
rect 30268 27694 30270 27746
rect 30322 27694 30324 27746
rect 30268 27682 30324 27694
rect 30156 27468 30436 27524
rect 29932 27356 30212 27412
rect 30156 26964 30212 27356
rect 30156 26908 30324 26964
rect 29932 26738 29988 26750
rect 30156 26740 30212 26750
rect 29932 26686 29934 26738
rect 29986 26686 29988 26738
rect 29932 26068 29988 26686
rect 29932 26002 29988 26012
rect 30044 26738 30212 26740
rect 30044 26686 30158 26738
rect 30210 26686 30212 26738
rect 30044 26684 30212 26686
rect 29932 25618 29988 25630
rect 29932 25566 29934 25618
rect 29986 25566 29988 25618
rect 29932 24946 29988 25566
rect 29932 24894 29934 24946
rect 29986 24894 29988 24946
rect 29932 24882 29988 24894
rect 30044 24948 30100 26684
rect 30156 26674 30212 26684
rect 30268 26516 30324 26908
rect 30380 26738 30436 27468
rect 30604 27076 30660 28702
rect 30716 28642 30772 28924
rect 30716 28590 30718 28642
rect 30770 28590 30772 28642
rect 30716 28578 30772 28590
rect 30940 28084 30996 30156
rect 31388 30146 31444 30156
rect 31052 29876 31108 29886
rect 31388 29876 31444 29886
rect 31052 29874 31444 29876
rect 31052 29822 31054 29874
rect 31106 29822 31390 29874
rect 31442 29822 31444 29874
rect 31052 29820 31444 29822
rect 31052 29810 31108 29820
rect 31276 29540 31332 29820
rect 31388 29810 31444 29820
rect 31500 29652 31556 31502
rect 31724 30772 31780 33516
rect 31836 32116 31892 33628
rect 32060 33618 32116 33628
rect 32172 33572 32228 33582
rect 31948 32900 32004 32910
rect 32004 32844 32116 32900
rect 31948 32806 32004 32844
rect 31836 32050 31892 32060
rect 31948 32562 32004 32574
rect 31948 32510 31950 32562
rect 32002 32510 32004 32562
rect 31836 31892 31892 31902
rect 31836 31798 31892 31836
rect 31724 30716 31892 30772
rect 31724 30548 31780 30558
rect 31276 29474 31332 29484
rect 31388 29596 31556 29652
rect 31612 30546 31780 30548
rect 31612 30494 31726 30546
rect 31778 30494 31780 30546
rect 31612 30492 31780 30494
rect 31612 29652 31668 30492
rect 31724 30482 31780 30492
rect 31276 29092 31332 29102
rect 31052 28754 31108 28766
rect 31052 28702 31054 28754
rect 31106 28702 31108 28754
rect 31052 28644 31108 28702
rect 31052 28578 31108 28588
rect 31276 28642 31332 29036
rect 31276 28590 31278 28642
rect 31330 28590 31332 28642
rect 30940 28028 31108 28084
rect 30828 27972 30884 27982
rect 30828 27878 30884 27916
rect 30716 27748 30772 27758
rect 30716 27746 30884 27748
rect 30716 27694 30718 27746
rect 30770 27694 30884 27746
rect 30716 27692 30884 27694
rect 30716 27682 30772 27692
rect 30716 27076 30772 27086
rect 30604 27074 30772 27076
rect 30604 27022 30718 27074
rect 30770 27022 30772 27074
rect 30604 27020 30772 27022
rect 30716 27010 30772 27020
rect 30828 26908 30884 27692
rect 30716 26852 30884 26908
rect 30940 27746 30996 27758
rect 30940 27694 30942 27746
rect 30994 27694 30996 27746
rect 30380 26686 30382 26738
rect 30434 26686 30436 26738
rect 30380 26674 30436 26686
rect 30604 26740 30660 26750
rect 30604 26646 30660 26684
rect 30156 26460 30324 26516
rect 30156 26180 30212 26460
rect 30156 26114 30212 26124
rect 30604 26292 30660 26302
rect 30268 25732 30324 25742
rect 30492 25732 30548 25742
rect 30268 25730 30548 25732
rect 30268 25678 30270 25730
rect 30322 25678 30494 25730
rect 30546 25678 30548 25730
rect 30268 25676 30548 25678
rect 30268 25666 30324 25676
rect 30492 25666 30548 25676
rect 30604 25730 30660 26236
rect 30604 25678 30606 25730
rect 30658 25678 30660 25730
rect 30604 25666 30660 25678
rect 30156 25508 30212 25518
rect 30156 25414 30212 25452
rect 30716 25060 30772 26852
rect 30828 25844 30884 25854
rect 30828 25750 30884 25788
rect 30716 24994 30772 25004
rect 30044 24882 30100 24892
rect 30828 24948 30884 24958
rect 30940 24948 30996 27694
rect 31052 26908 31108 28028
rect 31164 27748 31220 27758
rect 31276 27748 31332 28590
rect 31164 27746 31332 27748
rect 31164 27694 31166 27746
rect 31218 27694 31332 27746
rect 31164 27692 31332 27694
rect 31388 27746 31444 29596
rect 31612 29092 31668 29596
rect 31724 29986 31780 29998
rect 31724 29934 31726 29986
rect 31778 29934 31780 29986
rect 31724 29316 31780 29934
rect 31836 29652 31892 30716
rect 31836 29586 31892 29596
rect 31724 29260 31892 29316
rect 31724 29092 31780 29102
rect 31612 29036 31724 29092
rect 31724 29026 31780 29036
rect 31500 28868 31556 28878
rect 31500 28774 31556 28812
rect 31388 27694 31390 27746
rect 31442 27694 31444 27746
rect 31164 27682 31220 27692
rect 31388 27682 31444 27694
rect 31500 28530 31556 28542
rect 31500 28478 31502 28530
rect 31554 28478 31556 28530
rect 31500 27636 31556 28478
rect 31836 28420 31892 29260
rect 31836 28354 31892 28364
rect 31500 27570 31556 27580
rect 31836 27970 31892 27982
rect 31836 27918 31838 27970
rect 31890 27918 31892 27970
rect 31052 26852 31668 26908
rect 31164 26740 31220 26750
rect 31500 26740 31556 26750
rect 31612 26740 31668 26796
rect 31164 26738 31668 26740
rect 31164 26686 31166 26738
rect 31218 26686 31502 26738
rect 31554 26686 31668 26738
rect 31164 26684 31668 26686
rect 31164 26674 31220 26684
rect 31500 26674 31556 26684
rect 31388 26516 31444 26526
rect 31388 25956 31444 26460
rect 31388 25842 31444 25900
rect 31388 25790 31390 25842
rect 31442 25790 31444 25842
rect 31388 25778 31444 25790
rect 31612 25842 31668 26684
rect 31724 26738 31780 26750
rect 31724 26686 31726 26738
rect 31778 26686 31780 26738
rect 31724 26628 31780 26686
rect 31724 26562 31780 26572
rect 31724 26292 31780 26302
rect 31836 26292 31892 27918
rect 31948 26740 32004 32510
rect 32060 32004 32116 32844
rect 32172 32786 32228 33516
rect 32172 32734 32174 32786
rect 32226 32734 32228 32786
rect 32172 32722 32228 32734
rect 32284 32676 32340 34748
rect 32508 34580 32564 36540
rect 32508 34514 32564 34524
rect 32620 38498 32788 38500
rect 32620 38446 32734 38498
rect 32786 38446 32788 38498
rect 32620 38444 32788 38446
rect 32396 33796 32452 33806
rect 32396 33702 32452 33740
rect 32508 33460 32564 33470
rect 32508 33366 32564 33404
rect 32508 32676 32564 32686
rect 32284 32674 32564 32676
rect 32284 32622 32510 32674
rect 32562 32622 32564 32674
rect 32284 32620 32564 32622
rect 32508 32610 32564 32620
rect 32620 32228 32676 38444
rect 32732 38434 32788 38444
rect 33068 37154 33124 38612
rect 33740 38162 33796 38670
rect 34524 38500 34580 39454
rect 35196 39340 35460 39350
rect 35252 39284 35300 39340
rect 35356 39284 35404 39340
rect 35196 39274 35460 39284
rect 34524 38434 34580 38444
rect 34748 38948 34804 38958
rect 33740 38110 33742 38162
rect 33794 38110 33796 38162
rect 33740 38098 33796 38110
rect 33068 37102 33070 37154
rect 33122 37102 33124 37154
rect 33068 37090 33124 37102
rect 34636 35588 34692 35598
rect 34300 35532 34636 35588
rect 32732 34804 32788 34814
rect 33068 34804 33124 34814
rect 32788 34802 33124 34804
rect 32788 34750 33070 34802
rect 33122 34750 33124 34802
rect 32788 34748 33124 34750
rect 32732 34738 32788 34748
rect 33068 34738 33124 34748
rect 33404 34690 33460 34702
rect 33404 34638 33406 34690
rect 33458 34638 33460 34690
rect 32732 34580 32788 34590
rect 32732 33796 32788 34524
rect 33180 34578 33236 34590
rect 33180 34526 33182 34578
rect 33234 34526 33236 34578
rect 33180 33908 33236 34526
rect 33404 34580 33460 34638
rect 33404 34514 33460 34524
rect 34076 34690 34132 34702
rect 34076 34638 34078 34690
rect 34130 34638 34132 34690
rect 33180 33842 33236 33852
rect 34076 33906 34132 34638
rect 34076 33854 34078 33906
rect 34130 33854 34132 33906
rect 34076 33842 34132 33854
rect 32732 33730 32788 33740
rect 33516 33796 33572 33806
rect 33516 33702 33572 33740
rect 34076 33684 34132 33694
rect 33068 33460 33124 33470
rect 33292 33460 33348 33470
rect 33068 33458 33236 33460
rect 33068 33406 33070 33458
rect 33122 33406 33236 33458
rect 33068 33404 33236 33406
rect 33068 33394 33124 33404
rect 32620 32162 32676 32172
rect 32844 32562 32900 32574
rect 32844 32510 32846 32562
rect 32898 32510 32900 32562
rect 32172 32004 32228 32014
rect 32060 32002 32228 32004
rect 32060 31950 32174 32002
rect 32226 31950 32228 32002
rect 32060 31948 32228 31950
rect 32172 31938 32228 31948
rect 32508 31892 32564 31902
rect 32844 31892 32900 32510
rect 33068 32452 33124 32462
rect 32508 31890 32900 31892
rect 32508 31838 32510 31890
rect 32562 31838 32900 31890
rect 32508 31836 32900 31838
rect 32956 32450 33124 32452
rect 32956 32398 33070 32450
rect 33122 32398 33124 32450
rect 32956 32396 33124 32398
rect 32508 31826 32564 31836
rect 32284 30882 32340 30894
rect 32284 30830 32286 30882
rect 32338 30830 32340 30882
rect 32060 30660 32116 30670
rect 32060 30566 32116 30604
rect 32172 29988 32228 29998
rect 32284 29988 32340 30830
rect 32620 30100 32676 31836
rect 32732 31668 32788 31678
rect 32732 30882 32788 31612
rect 32956 31106 33012 32396
rect 33068 32386 33124 32396
rect 33068 32228 33124 32238
rect 33068 31778 33124 32172
rect 33068 31726 33070 31778
rect 33122 31726 33124 31778
rect 33068 31714 33124 31726
rect 32956 31054 32958 31106
rect 33010 31054 33012 31106
rect 32956 31042 33012 31054
rect 32732 30830 32734 30882
rect 32786 30830 32788 30882
rect 32732 30770 32788 30830
rect 32732 30718 32734 30770
rect 32786 30718 32788 30770
rect 32732 30706 32788 30718
rect 32844 30882 32900 30894
rect 32844 30830 32846 30882
rect 32898 30830 32900 30882
rect 32620 30034 32676 30044
rect 32172 29986 32340 29988
rect 32172 29934 32174 29986
rect 32226 29934 32340 29986
rect 32172 29932 32340 29934
rect 32172 29922 32228 29932
rect 32508 29876 32564 29886
rect 32508 29874 32676 29876
rect 32508 29822 32510 29874
rect 32562 29822 32676 29874
rect 32508 29820 32676 29822
rect 32508 29810 32564 29820
rect 32172 29652 32228 29662
rect 32172 29316 32228 29596
rect 32060 28756 32116 28766
rect 32172 28756 32228 29260
rect 32620 28868 32676 29820
rect 32508 28756 32564 28766
rect 32060 28754 32564 28756
rect 32060 28702 32062 28754
rect 32114 28702 32510 28754
rect 32562 28702 32564 28754
rect 32060 28700 32564 28702
rect 32060 28690 32116 28700
rect 32508 28690 32564 28700
rect 32396 28532 32452 28542
rect 32172 28530 32452 28532
rect 32172 28478 32398 28530
rect 32450 28478 32452 28530
rect 32172 28476 32452 28478
rect 32172 27858 32228 28476
rect 32396 28466 32452 28476
rect 32620 28532 32676 28812
rect 32844 28754 32900 30830
rect 33180 30770 33236 33404
rect 33348 33404 33572 33460
rect 33292 33394 33348 33404
rect 33516 32786 33572 33404
rect 33516 32734 33518 32786
rect 33570 32734 33572 32786
rect 33516 32722 33572 32734
rect 34076 32674 34132 33628
rect 34188 33682 34244 33694
rect 34188 33630 34190 33682
rect 34242 33630 34244 33682
rect 34188 33460 34244 33630
rect 34188 32898 34244 33404
rect 34188 32846 34190 32898
rect 34242 32846 34244 32898
rect 34188 32834 34244 32846
rect 34076 32622 34078 32674
rect 34130 32622 34132 32674
rect 34076 32610 34132 32622
rect 33292 31890 33348 31902
rect 33292 31838 33294 31890
rect 33346 31838 33348 31890
rect 33292 31668 33348 31838
rect 33516 31790 33572 31802
rect 33516 31738 33518 31790
rect 33570 31780 33572 31790
rect 33628 31780 33684 31790
rect 33570 31738 33628 31780
rect 33516 31724 33628 31738
rect 33684 31724 34020 31780
rect 33628 31714 33684 31724
rect 33292 31612 33572 31668
rect 33516 31556 33572 31612
rect 33516 31500 33684 31556
rect 33404 31444 33460 31454
rect 33180 30718 33182 30770
rect 33234 30718 33236 30770
rect 33180 30706 33236 30718
rect 33292 31442 33460 31444
rect 33292 31390 33406 31442
rect 33458 31390 33460 31442
rect 33292 31388 33460 31390
rect 32956 30658 33012 30670
rect 32956 30606 32958 30658
rect 33010 30606 33012 30658
rect 32956 30548 33012 30606
rect 33292 30548 33348 31388
rect 33404 31378 33460 31388
rect 33516 30882 33572 30894
rect 33516 30830 33518 30882
rect 33570 30830 33572 30882
rect 33516 30770 33572 30830
rect 33516 30718 33518 30770
rect 33570 30718 33572 30770
rect 33516 30706 33572 30718
rect 32956 30482 33012 30492
rect 33068 30492 33348 30548
rect 33628 30660 33684 31500
rect 33852 30882 33908 30894
rect 33852 30830 33854 30882
rect 33906 30830 33908 30882
rect 33740 30660 33796 30670
rect 33628 30658 33796 30660
rect 33628 30606 33742 30658
rect 33794 30606 33796 30658
rect 33628 30604 33796 30606
rect 33628 30548 33684 30604
rect 33740 30594 33796 30604
rect 33068 29762 33124 30492
rect 33516 29876 33572 29886
rect 33068 29710 33070 29762
rect 33122 29710 33124 29762
rect 33068 29698 33124 29710
rect 33180 29764 33236 29774
rect 33180 29670 33236 29708
rect 33292 29764 33348 29774
rect 33292 29762 33460 29764
rect 33292 29710 33294 29762
rect 33346 29710 33460 29762
rect 33292 29708 33460 29710
rect 33292 29698 33348 29708
rect 33292 28980 33348 28990
rect 32844 28702 32846 28754
rect 32898 28702 32900 28754
rect 32844 28690 32900 28702
rect 32956 28756 33012 28766
rect 32956 28662 33012 28700
rect 33068 28756 33124 28766
rect 33068 28754 33236 28756
rect 33068 28702 33070 28754
rect 33122 28702 33236 28754
rect 33068 28700 33236 28702
rect 33068 28690 33124 28700
rect 32620 28466 32676 28476
rect 32172 27806 32174 27858
rect 32226 27806 32228 27858
rect 32172 27748 32228 27806
rect 32172 27682 32228 27692
rect 32620 27860 32676 27870
rect 31948 26674 32004 26684
rect 32284 26852 32340 26862
rect 32284 26738 32340 26796
rect 32284 26686 32286 26738
rect 32338 26686 32340 26738
rect 32284 26674 32340 26686
rect 32508 26740 32564 26750
rect 32060 26516 32116 26526
rect 32060 26422 32116 26460
rect 31780 26236 31892 26292
rect 32508 26292 32564 26684
rect 31724 26226 31780 26236
rect 32508 26226 32564 26236
rect 32508 25956 32564 25966
rect 32620 25956 32676 27804
rect 33068 27746 33124 27758
rect 33068 27694 33070 27746
rect 33122 27694 33124 27746
rect 33068 26964 33124 27694
rect 33180 27524 33236 28700
rect 33180 27458 33236 27468
rect 33292 28754 33348 28924
rect 33292 28702 33294 28754
rect 33346 28702 33348 28754
rect 33180 26964 33236 26974
rect 33068 26962 33236 26964
rect 33068 26910 33182 26962
rect 33234 26910 33236 26962
rect 33068 26908 33236 26910
rect 33180 26898 33236 26908
rect 32508 25954 32676 25956
rect 32508 25902 32510 25954
rect 32562 25902 32676 25954
rect 32508 25900 32676 25902
rect 32844 26738 32900 26750
rect 32844 26686 32846 26738
rect 32898 26686 32900 26738
rect 32508 25890 32564 25900
rect 31612 25790 31614 25842
rect 31666 25790 31668 25842
rect 31164 25620 31220 25630
rect 31164 25526 31220 25564
rect 31388 24948 31444 24958
rect 30940 24946 31444 24948
rect 30940 24894 31390 24946
rect 31442 24894 31444 24946
rect 30940 24892 31444 24894
rect 30828 24854 30884 24892
rect 31388 24882 31444 24892
rect 29820 24668 29988 24724
rect 29596 24610 29652 24622
rect 29596 24558 29598 24610
rect 29650 24558 29652 24610
rect 29596 24500 29652 24558
rect 29596 24434 29652 24444
rect 29820 24498 29876 24510
rect 29820 24446 29822 24498
rect 29874 24446 29876 24498
rect 29820 24388 29876 24446
rect 29820 24322 29876 24332
rect 29484 24220 29652 24276
rect 29372 23986 29428 23996
rect 29484 23716 29540 23726
rect 29260 23714 29540 23716
rect 29260 23662 29486 23714
rect 29538 23662 29540 23714
rect 29260 23660 29540 23662
rect 29260 22708 29316 22718
rect 29484 22708 29540 23660
rect 29260 22706 29540 22708
rect 29260 22654 29262 22706
rect 29314 22654 29486 22706
rect 29538 22654 29540 22706
rect 29260 22652 29540 22654
rect 29260 22642 29316 22652
rect 29484 22642 29540 22652
rect 29596 22594 29652 24220
rect 29596 22542 29598 22594
rect 29650 22542 29652 22594
rect 29596 22530 29652 22542
rect 29820 22594 29876 22606
rect 29820 22542 29822 22594
rect 29874 22542 29876 22594
rect 28588 22482 28644 22494
rect 28588 22430 28590 22482
rect 28642 22430 28644 22482
rect 28140 21812 28196 21822
rect 28140 20802 28196 21756
rect 28588 21700 28644 22430
rect 28700 21812 28756 21822
rect 28700 21718 28756 21756
rect 28588 21252 28644 21644
rect 28588 21186 28644 21196
rect 29148 21698 29204 21710
rect 29148 21646 29150 21698
rect 29202 21646 29204 21698
rect 28140 20750 28142 20802
rect 28194 20750 28196 20802
rect 28028 19570 28084 19582
rect 28028 19518 28030 19570
rect 28082 19518 28084 19570
rect 28028 18788 28084 19518
rect 28140 19010 28196 20750
rect 28476 20468 28532 20478
rect 28476 19570 28532 20412
rect 28588 20466 28644 20478
rect 28588 20414 28590 20466
rect 28642 20414 28644 20466
rect 28588 20356 28644 20414
rect 29148 20356 29204 21646
rect 29820 20916 29876 22542
rect 29932 22370 29988 24668
rect 30492 24668 30884 24724
rect 30268 24612 30324 24622
rect 30268 24518 30324 24556
rect 30492 24610 30548 24668
rect 30492 24558 30494 24610
rect 30546 24558 30548 24610
rect 30492 24546 30548 24558
rect 30604 24500 30660 24510
rect 30604 24276 30660 24444
rect 30492 24220 30660 24276
rect 30492 24164 30548 24220
rect 30156 24108 30548 24164
rect 29932 22318 29934 22370
rect 29986 22318 29988 22370
rect 29932 22306 29988 22318
rect 30044 22706 30100 22718
rect 30044 22654 30046 22706
rect 30098 22654 30100 22706
rect 30044 22596 30100 22654
rect 29820 20850 29876 20860
rect 29932 21812 29988 21822
rect 30044 21812 30100 22540
rect 30156 22484 30212 24108
rect 30604 24052 30660 24062
rect 30604 23958 30660 23996
rect 30716 23492 30772 23502
rect 30716 22706 30772 23436
rect 30716 22654 30718 22706
rect 30770 22654 30772 22706
rect 30156 22390 30212 22428
rect 30492 22594 30548 22606
rect 30492 22542 30494 22594
rect 30546 22542 30548 22594
rect 30492 21924 30548 22542
rect 30716 22372 30772 22654
rect 30716 22306 30772 22316
rect 30604 21924 30660 21934
rect 30492 21922 30660 21924
rect 30492 21870 30606 21922
rect 30658 21870 30660 21922
rect 30492 21868 30660 21870
rect 30604 21858 30660 21868
rect 29932 21810 30100 21812
rect 29932 21758 29934 21810
rect 29986 21758 30100 21810
rect 29932 21756 30100 21758
rect 30828 21812 30884 24668
rect 31052 24610 31108 24622
rect 31052 24558 31054 24610
rect 31106 24558 31108 24610
rect 31052 23940 31108 24558
rect 31276 24610 31332 24622
rect 31276 24558 31278 24610
rect 31330 24558 31332 24610
rect 31164 23940 31220 23950
rect 31052 23884 31164 23940
rect 31164 23874 31220 23884
rect 31164 22820 31220 22830
rect 30940 22764 31164 22820
rect 30940 22706 30996 22764
rect 30940 22654 30942 22706
rect 30994 22654 30996 22706
rect 30940 22642 30996 22654
rect 30940 21812 30996 21822
rect 30828 21810 30996 21812
rect 30828 21758 30942 21810
rect 30994 21758 30996 21810
rect 30828 21756 30996 21758
rect 28588 20300 29148 20356
rect 28476 19518 28478 19570
rect 28530 19518 28532 19570
rect 28140 18958 28142 19010
rect 28194 18958 28196 19010
rect 28140 18946 28196 18958
rect 28252 19458 28308 19470
rect 28252 19406 28254 19458
rect 28306 19406 28308 19458
rect 28252 18898 28308 19406
rect 28476 19460 28532 19518
rect 28924 19906 28980 20300
rect 29148 20290 29204 20300
rect 29484 20468 29540 20478
rect 28924 19854 28926 19906
rect 28978 19854 28980 19906
rect 28476 19404 28756 19460
rect 28252 18846 28254 18898
rect 28306 18846 28308 18898
rect 28028 18722 28084 18732
rect 28140 18788 28196 18798
rect 28252 18788 28308 18846
rect 28140 18786 28308 18788
rect 28140 18734 28142 18786
rect 28194 18734 28308 18786
rect 28140 18732 28308 18734
rect 28588 18788 28644 18798
rect 28140 18722 28196 18732
rect 28588 18694 28644 18732
rect 28700 18564 28756 19404
rect 28924 19458 28980 19854
rect 29260 19908 29316 19918
rect 29260 19682 29316 19852
rect 29260 19630 29262 19682
rect 29314 19630 29316 19682
rect 29260 19618 29316 19630
rect 28924 19406 28926 19458
rect 28978 19406 28980 19458
rect 28924 19394 28980 19406
rect 29484 18788 29540 20412
rect 29932 20466 29988 21756
rect 30940 21746 30996 21756
rect 31052 21812 31108 22764
rect 31164 22754 31220 22764
rect 31276 22706 31332 24558
rect 31500 24500 31556 24510
rect 31500 24406 31556 24444
rect 31388 23940 31444 23950
rect 31388 23846 31444 23884
rect 31612 23716 31668 25790
rect 31724 25732 31780 25742
rect 31724 25638 31780 25676
rect 31948 25732 32004 25742
rect 32172 25732 32228 25742
rect 31948 25730 32116 25732
rect 31948 25678 31950 25730
rect 32002 25678 32116 25730
rect 31948 25676 32116 25678
rect 31948 25666 32004 25676
rect 32060 25508 32116 25676
rect 32172 25638 32228 25676
rect 32620 25732 32676 25742
rect 31836 24610 31892 24622
rect 31836 24558 31838 24610
rect 31890 24558 31892 24610
rect 31724 23828 31780 23838
rect 31724 23716 31780 23772
rect 31612 23714 31780 23716
rect 31612 23662 31726 23714
rect 31778 23662 31780 23714
rect 31612 23660 31780 23662
rect 31500 23604 31556 23614
rect 31276 22654 31278 22706
rect 31330 22654 31332 22706
rect 31276 22642 31332 22654
rect 31388 23548 31500 23604
rect 31388 22706 31444 23548
rect 31500 23538 31556 23548
rect 31388 22654 31390 22706
rect 31442 22654 31444 22706
rect 31388 22642 31444 22654
rect 31164 22596 31220 22606
rect 31164 22502 31220 22540
rect 31612 22596 31668 23660
rect 31724 23650 31780 23660
rect 31836 22708 31892 24558
rect 31948 24612 32004 24622
rect 31948 24518 32004 24556
rect 31948 23714 32004 23726
rect 31948 23662 31950 23714
rect 32002 23662 32004 23714
rect 31948 23604 32004 23662
rect 32060 23716 32116 25452
rect 32060 23650 32116 23660
rect 32396 23714 32452 23726
rect 32396 23662 32398 23714
rect 32450 23662 32452 23714
rect 31948 23538 32004 23548
rect 32396 23492 32452 23662
rect 32508 23492 32564 23502
rect 32396 23436 32508 23492
rect 32508 23426 32564 23436
rect 31836 22652 32564 22708
rect 31612 22530 31668 22540
rect 31948 22484 32004 22494
rect 31836 22482 32004 22484
rect 31836 22430 31950 22482
rect 32002 22430 32004 22482
rect 31836 22428 32004 22430
rect 31836 22372 31892 22428
rect 31948 22418 32004 22428
rect 32284 22484 32340 22494
rect 32284 22390 32340 22428
rect 30268 21700 30324 21710
rect 30324 21644 30436 21700
rect 30268 21606 30324 21644
rect 30268 20916 30324 20926
rect 30268 20822 30324 20860
rect 29932 20414 29934 20466
rect 29986 20414 29988 20466
rect 29820 20356 29876 20366
rect 29708 20300 29820 20356
rect 29596 19796 29652 19806
rect 29596 19702 29652 19740
rect 29708 19682 29764 20300
rect 29820 20290 29876 20300
rect 29708 19630 29710 19682
rect 29762 19630 29764 19682
rect 29708 19572 29764 19630
rect 29596 19516 29764 19572
rect 29932 19684 29988 20414
rect 30380 20468 30436 21644
rect 30380 20402 30436 20412
rect 30492 20692 30548 20702
rect 30380 19908 30436 19918
rect 30268 19684 30324 19694
rect 29932 19628 30268 19684
rect 29596 19236 29652 19516
rect 29932 19460 29988 19628
rect 30268 19618 30324 19628
rect 29596 19170 29652 19180
rect 29708 19404 29988 19460
rect 29484 18722 29540 18732
rect 29596 18564 29652 18574
rect 29708 18564 29764 19404
rect 28700 18562 29764 18564
rect 28700 18510 29598 18562
rect 29650 18510 29764 18562
rect 28700 18508 29764 18510
rect 29932 19236 29988 19246
rect 28812 18340 28868 18350
rect 28028 17778 28084 17790
rect 28028 17726 28030 17778
rect 28082 17726 28084 17778
rect 28028 16660 28084 17726
rect 28700 17668 28756 17678
rect 28028 16594 28084 16604
rect 28476 17666 28756 17668
rect 28476 17614 28702 17666
rect 28754 17614 28756 17666
rect 28476 17612 28756 17614
rect 28252 16434 28308 16446
rect 28252 16382 28254 16434
rect 28306 16382 28308 16434
rect 28028 16324 28084 16334
rect 28252 16324 28308 16382
rect 28084 16268 28308 16324
rect 28028 16258 28084 16268
rect 28476 15874 28532 17612
rect 28700 17602 28756 17612
rect 28812 16884 28868 18284
rect 28588 16548 28644 16558
rect 28812 16548 28868 16828
rect 28588 16546 28868 16548
rect 28588 16494 28590 16546
rect 28642 16494 28868 16546
rect 28588 16492 28868 16494
rect 28588 16482 28644 16492
rect 28476 15822 28478 15874
rect 28530 15822 28532 15874
rect 28476 15810 28532 15822
rect 28812 15764 28868 15774
rect 28924 15764 28980 18508
rect 29596 18498 29652 18508
rect 29820 18452 29876 18462
rect 29820 17890 29876 18396
rect 29820 17838 29822 17890
rect 29874 17838 29876 17890
rect 29820 17826 29876 17838
rect 29260 17666 29316 17678
rect 29260 17614 29262 17666
rect 29314 17614 29316 17666
rect 29260 16772 29316 17614
rect 29260 16706 29316 16716
rect 29372 16884 29428 16894
rect 28812 15762 28980 15764
rect 28812 15710 28814 15762
rect 28866 15710 28980 15762
rect 28812 15708 28980 15710
rect 29148 16546 29204 16558
rect 29148 16494 29150 16546
rect 29202 16494 29204 16546
rect 28252 15652 28308 15662
rect 28252 15650 28532 15652
rect 28252 15598 28254 15650
rect 28306 15598 28532 15650
rect 28252 15596 28532 15598
rect 28252 15586 28308 15596
rect 28364 15428 28420 15438
rect 28140 14420 28196 14430
rect 28140 14326 28196 14364
rect 28252 14306 28308 14318
rect 28252 14254 28254 14306
rect 28306 14254 28308 14306
rect 28140 13636 28196 13646
rect 28140 13542 28196 13580
rect 28028 13412 28084 13422
rect 28028 11844 28084 13356
rect 28028 11778 28084 11788
rect 28252 11506 28308 14254
rect 28364 12964 28420 15372
rect 28476 15316 28532 15596
rect 28476 15148 28532 15260
rect 28476 15092 28644 15148
rect 28588 14418 28644 15092
rect 28812 14868 28868 15708
rect 29036 15540 29092 15550
rect 29148 15540 29204 16494
rect 29036 15538 29204 15540
rect 29036 15486 29038 15538
rect 29090 15486 29204 15538
rect 29036 15484 29204 15486
rect 29036 15148 29092 15484
rect 29036 15092 29316 15148
rect 28812 14802 28868 14812
rect 28588 14366 28590 14418
rect 28642 14366 28644 14418
rect 28588 13524 28644 14366
rect 29260 14420 29316 15092
rect 29372 14754 29428 16828
rect 29820 16660 29876 16670
rect 29932 16660 29988 19180
rect 29820 16658 29988 16660
rect 29820 16606 29822 16658
rect 29874 16606 29988 16658
rect 29820 16604 29988 16606
rect 29820 16594 29876 16604
rect 29484 16546 29540 16558
rect 29484 16494 29486 16546
rect 29538 16494 29540 16546
rect 29484 15204 29540 16494
rect 29932 15764 29988 16604
rect 30156 17666 30212 17678
rect 30156 17614 30158 17666
rect 30210 17614 30212 17666
rect 30156 16658 30212 17614
rect 30380 17556 30436 19852
rect 30492 17778 30548 20636
rect 30604 20692 30660 20702
rect 30828 20692 30884 20702
rect 31052 20692 31108 21756
rect 31164 21812 31220 21822
rect 31724 21812 31780 21822
rect 31164 21810 31780 21812
rect 31164 21758 31166 21810
rect 31218 21758 31726 21810
rect 31778 21758 31780 21810
rect 31164 21756 31780 21758
rect 31164 21746 31220 21756
rect 31724 21746 31780 21756
rect 31164 20692 31220 20702
rect 30604 20690 30772 20692
rect 30604 20638 30606 20690
rect 30658 20638 30772 20690
rect 30604 20636 30772 20638
rect 30604 20626 30660 20636
rect 30716 19906 30772 20636
rect 30828 20598 30884 20636
rect 30940 20690 31220 20692
rect 30940 20638 31166 20690
rect 31218 20638 31220 20690
rect 30940 20636 31220 20638
rect 30716 19854 30718 19906
rect 30770 19854 30772 19906
rect 30716 19842 30772 19854
rect 30828 20468 30884 20478
rect 30828 19794 30884 20412
rect 30828 19742 30830 19794
rect 30882 19742 30884 19794
rect 30828 19730 30884 19742
rect 30604 19682 30660 19694
rect 30604 19630 30606 19682
rect 30658 19630 30660 19682
rect 30604 19572 30660 19630
rect 30940 19572 30996 20636
rect 31164 20626 31220 20636
rect 31388 20690 31444 20702
rect 31388 20638 31390 20690
rect 31442 20638 31444 20690
rect 31276 20468 31332 20478
rect 31388 20468 31444 20638
rect 31332 20412 31444 20468
rect 31276 20402 31332 20412
rect 31052 19684 31108 19694
rect 31052 19590 31108 19628
rect 30604 19516 30996 19572
rect 30940 19460 30996 19516
rect 30940 19404 31332 19460
rect 31276 18562 31332 19404
rect 31276 18510 31278 18562
rect 31330 18510 31332 18562
rect 31276 18498 31332 18510
rect 31388 18730 31444 20412
rect 31612 20690 31668 20702
rect 31612 20638 31614 20690
rect 31666 20638 31668 20690
rect 31612 19684 31668 20638
rect 31836 20578 31892 22316
rect 31948 21698 32004 21710
rect 31948 21646 31950 21698
rect 32002 21646 32004 21698
rect 31948 20690 32004 21646
rect 31948 20638 31950 20690
rect 32002 20638 32004 20690
rect 31948 20626 32004 20638
rect 32284 21698 32340 21710
rect 32284 21646 32286 21698
rect 32338 21646 32340 21698
rect 32284 20692 32340 21646
rect 32508 20914 32564 22652
rect 32620 22594 32676 25676
rect 32844 25620 32900 26686
rect 33292 26740 33348 28702
rect 33404 28082 33460 29708
rect 33516 29762 33572 29820
rect 33516 29710 33518 29762
rect 33570 29710 33572 29762
rect 33516 28980 33572 29710
rect 33516 28914 33572 28924
rect 33516 28754 33572 28766
rect 33516 28702 33518 28754
rect 33570 28702 33572 28754
rect 33516 28196 33572 28702
rect 33516 28130 33572 28140
rect 33404 28030 33406 28082
rect 33458 28030 33460 28082
rect 33404 28018 33460 28030
rect 33404 27858 33460 27870
rect 33404 27806 33406 27858
rect 33458 27806 33460 27858
rect 33404 26908 33460 27806
rect 33516 27860 33572 27870
rect 33516 27766 33572 27804
rect 33628 27188 33684 30492
rect 33740 29764 33796 29774
rect 33740 29670 33796 29708
rect 33852 28756 33908 30830
rect 33964 30770 34020 31724
rect 33964 30718 33966 30770
rect 34018 30718 34020 30770
rect 33964 30706 34020 30718
rect 34188 29986 34244 29998
rect 34188 29934 34190 29986
rect 34242 29934 34244 29986
rect 34188 29876 34244 29934
rect 34188 29810 34244 29820
rect 33964 28756 34020 28766
rect 33852 28754 34020 28756
rect 33852 28702 33966 28754
rect 34018 28702 34020 28754
rect 33852 28700 34020 28702
rect 33964 28690 34020 28700
rect 34188 28754 34244 28766
rect 34188 28702 34190 28754
rect 34242 28702 34244 28754
rect 34076 28644 34132 28654
rect 34076 28550 34132 28588
rect 34188 28084 34244 28702
rect 34300 28532 34356 35532
rect 34636 35494 34692 35532
rect 34748 34914 34804 38892
rect 36092 38948 36148 39566
rect 36092 38882 36148 38892
rect 36316 38164 36372 38174
rect 36428 38164 36484 39676
rect 36988 39730 37044 39742
rect 36988 39678 36990 39730
rect 37042 39678 37044 39730
rect 36988 39620 37044 39678
rect 36988 39058 37044 39564
rect 36988 39006 36990 39058
rect 37042 39006 37044 39058
rect 36988 38994 37044 39006
rect 37212 39170 37268 39182
rect 37212 39118 37214 39170
rect 37266 39118 37268 39170
rect 37212 38948 37268 39118
rect 37324 39172 37380 40798
rect 37436 40180 37492 41804
rect 37548 41746 37604 41758
rect 37548 41694 37550 41746
rect 37602 41694 37604 41746
rect 37548 41636 37604 41694
rect 37548 41570 37604 41580
rect 37884 40964 37940 41916
rect 37996 41906 38052 41916
rect 38668 41748 38724 42028
rect 38668 40964 38724 41692
rect 38892 41636 38948 44044
rect 39004 43876 39060 44604
rect 39004 43810 39060 43820
rect 40012 43876 40068 43886
rect 39340 43652 39396 43662
rect 39340 43650 39732 43652
rect 39340 43598 39342 43650
rect 39394 43598 39732 43650
rect 39340 43596 39732 43598
rect 39340 43586 39396 43596
rect 39676 42866 39732 43596
rect 39676 42814 39678 42866
rect 39730 42814 39732 42866
rect 39676 42802 39732 42814
rect 40012 42754 40068 43820
rect 40124 43708 40180 45612
rect 40908 43986 40964 46172
rect 41132 46114 41188 46844
rect 41244 46676 41300 48750
rect 41356 48804 41412 49758
rect 41804 49810 41860 49822
rect 41804 49758 41806 49810
rect 41858 49758 41860 49810
rect 41692 49028 41748 49038
rect 41692 48934 41748 48972
rect 41804 48916 41860 49758
rect 42252 49810 42308 49822
rect 42252 49758 42254 49810
rect 42306 49758 42308 49810
rect 42252 49028 42308 49758
rect 42364 49028 42420 49038
rect 42252 48972 42364 49028
rect 41804 48850 41860 48860
rect 42140 48916 42196 48926
rect 41356 48738 41412 48748
rect 42140 48802 42196 48860
rect 42140 48750 42142 48802
rect 42194 48750 42196 48802
rect 42140 48738 42196 48750
rect 42364 48802 42420 48972
rect 43484 48916 43540 48926
rect 42364 48750 42366 48802
rect 42418 48750 42420 48802
rect 42364 48738 42420 48750
rect 42812 48804 42868 48814
rect 42812 48692 42868 48748
rect 43372 48692 43428 48702
rect 42812 48690 43428 48692
rect 42812 48638 43374 48690
rect 43426 48638 43428 48690
rect 42812 48636 43428 48638
rect 41804 48132 41860 48142
rect 41804 48130 41972 48132
rect 41804 48078 41806 48130
rect 41858 48078 41972 48130
rect 41804 48076 41972 48078
rect 41804 48066 41860 48076
rect 41244 46610 41300 46620
rect 41468 47906 41524 47918
rect 41468 47854 41470 47906
rect 41522 47854 41524 47906
rect 41132 46062 41134 46114
rect 41186 46062 41188 46114
rect 41132 46050 41188 46062
rect 41468 45556 41524 47854
rect 41580 46676 41636 46686
rect 41580 46114 41636 46620
rect 41580 46062 41582 46114
rect 41634 46062 41636 46114
rect 41580 46050 41636 46062
rect 41916 45668 41972 48076
rect 42812 48020 42868 48636
rect 43372 48626 43428 48636
rect 42812 48018 42980 48020
rect 42812 47966 42814 48018
rect 42866 47966 42980 48018
rect 42812 47964 42980 47966
rect 42812 47954 42868 47964
rect 42924 46674 42980 47964
rect 43484 47906 43540 48860
rect 43708 48916 43764 48926
rect 43708 48130 43764 48860
rect 44156 48692 44212 48702
rect 43708 48078 43710 48130
rect 43762 48078 43764 48130
rect 43708 48066 43764 48078
rect 43820 48690 44212 48692
rect 43820 48638 44158 48690
rect 44210 48638 44212 48690
rect 43820 48636 44212 48638
rect 43484 47854 43486 47906
rect 43538 47854 43540 47906
rect 43484 47842 43540 47854
rect 42924 46622 42926 46674
rect 42978 46622 42980 46674
rect 41916 45612 42420 45668
rect 41468 45500 41636 45556
rect 41468 45332 41524 45342
rect 41468 44882 41524 45276
rect 41468 44830 41470 44882
rect 41522 44830 41524 44882
rect 41468 44818 41524 44830
rect 41132 44660 41188 44670
rect 41132 44566 41188 44604
rect 40908 43934 40910 43986
rect 40962 43934 40964 43986
rect 40908 43922 40964 43934
rect 41580 43986 41636 45500
rect 42252 44660 42308 44670
rect 41580 43934 41582 43986
rect 41634 43934 41636 43986
rect 41580 43922 41636 43934
rect 41804 44658 42308 44660
rect 41804 44606 42254 44658
rect 42306 44606 42308 44658
rect 41804 44604 42308 44606
rect 41244 43876 41300 43886
rect 41244 43782 41300 43820
rect 40124 43652 40404 43708
rect 40348 42866 40404 43652
rect 40348 42814 40350 42866
rect 40402 42814 40404 42866
rect 40348 42802 40404 42814
rect 41804 42866 41860 44604
rect 42252 44594 42308 44604
rect 41804 42814 41806 42866
rect 41858 42814 41860 42866
rect 41804 42802 41860 42814
rect 41916 43874 41972 43886
rect 41916 43822 41918 43874
rect 41970 43822 41972 43874
rect 40012 42702 40014 42754
rect 40066 42702 40068 42754
rect 40012 41860 40068 42702
rect 41132 42754 41188 42766
rect 41132 42702 41134 42754
rect 41186 42702 41188 42754
rect 40684 42644 40740 42654
rect 40684 42642 40852 42644
rect 40684 42590 40686 42642
rect 40738 42590 40852 42642
rect 40684 42588 40852 42590
rect 40684 42578 40740 42588
rect 40012 41794 40068 41804
rect 39900 41748 39956 41758
rect 37884 40850 37940 40908
rect 37884 40798 37886 40850
rect 37938 40798 37940 40850
rect 37884 40786 37940 40798
rect 38444 40908 38724 40964
rect 37660 40738 37716 40750
rect 37660 40686 37662 40738
rect 37714 40686 37716 40738
rect 37660 40516 37716 40686
rect 37716 40460 38164 40516
rect 37660 40450 37716 40460
rect 37548 40180 37604 40190
rect 37436 40178 37604 40180
rect 37436 40126 37550 40178
rect 37602 40126 37604 40178
rect 37436 40124 37604 40126
rect 37548 40114 37604 40124
rect 37884 39842 37940 39854
rect 37884 39790 37886 39842
rect 37938 39790 37940 39842
rect 37884 39732 37940 39790
rect 37324 39116 37716 39172
rect 37548 38948 37604 38958
rect 37212 38946 37380 38948
rect 37212 38894 37214 38946
rect 37266 38894 37380 38946
rect 37212 38892 37380 38894
rect 37212 38882 37268 38892
rect 36316 38162 36484 38164
rect 36316 38110 36318 38162
rect 36370 38110 36484 38162
rect 36316 38108 36484 38110
rect 36316 38098 36372 38108
rect 35308 37826 35364 37838
rect 35308 37774 35310 37826
rect 35362 37774 35364 37826
rect 35308 37716 35364 37774
rect 35308 37650 35364 37660
rect 36652 37826 36708 37838
rect 36652 37774 36654 37826
rect 36706 37774 36708 37826
rect 35196 37324 35460 37334
rect 35252 37268 35300 37324
rect 35356 37268 35404 37324
rect 35196 37258 35460 37268
rect 35980 36596 36036 36606
rect 36428 36596 36484 36606
rect 36652 36596 36708 37774
rect 37324 36932 37380 38892
rect 37324 36930 37492 36932
rect 37324 36878 37326 36930
rect 37378 36878 37492 36930
rect 37324 36876 37492 36878
rect 37324 36866 37380 36876
rect 35980 36594 36428 36596
rect 35980 36542 35982 36594
rect 36034 36542 36428 36594
rect 35980 36540 36428 36542
rect 36484 36540 36708 36596
rect 34972 35812 35028 35822
rect 34972 35718 35028 35756
rect 35980 35588 36036 36540
rect 36428 36502 36484 36540
rect 36428 36148 36484 36158
rect 36316 36036 36372 36046
rect 36428 36036 36484 36092
rect 36316 36034 36484 36036
rect 36316 35982 36318 36034
rect 36370 35982 36484 36034
rect 36316 35980 36484 35982
rect 36876 36148 36932 36158
rect 36316 35970 36372 35980
rect 35980 35522 36036 35532
rect 36204 35812 36260 35822
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34748 34862 34750 34914
rect 34802 34862 34804 34914
rect 34412 34580 34468 34590
rect 34412 32900 34468 34524
rect 34748 33460 34804 34862
rect 35644 34916 35700 34926
rect 35644 34822 35700 34860
rect 36092 34804 36148 34814
rect 36092 34710 36148 34748
rect 35196 34692 35252 34702
rect 35196 34598 35252 34636
rect 35196 34020 35252 34030
rect 34972 33908 35028 33918
rect 34860 33796 34916 33806
rect 34860 33702 34916 33740
rect 34748 33394 34804 33404
rect 34748 33122 34804 33134
rect 34748 33070 34750 33122
rect 34802 33070 34804 33122
rect 34748 32900 34804 33070
rect 34412 32898 34804 32900
rect 34412 32846 34750 32898
rect 34802 32846 34804 32898
rect 34412 32844 34804 32846
rect 34412 31778 34468 32844
rect 34748 32834 34804 32844
rect 34412 31726 34414 31778
rect 34466 31726 34468 31778
rect 34412 31714 34468 31726
rect 34748 31780 34804 31790
rect 34748 31686 34804 31724
rect 34412 30660 34468 30670
rect 34412 30566 34468 30604
rect 34748 30546 34804 30558
rect 34748 30494 34750 30546
rect 34802 30494 34804 30546
rect 34524 29876 34580 29886
rect 34748 29876 34804 30494
rect 34524 29874 34804 29876
rect 34524 29822 34526 29874
rect 34578 29822 34804 29874
rect 34524 29820 34804 29822
rect 34860 30212 34916 30222
rect 34524 29652 34580 29820
rect 34860 29764 34916 30156
rect 34524 29586 34580 29596
rect 34748 29762 34916 29764
rect 34748 29710 34862 29762
rect 34914 29710 34916 29762
rect 34748 29708 34916 29710
rect 34636 29316 34692 29326
rect 34748 29316 34804 29708
rect 34860 29698 34916 29708
rect 34692 29260 34804 29316
rect 34860 29540 34916 29550
rect 34636 29250 34692 29260
rect 34524 28980 34580 28990
rect 34412 28924 34524 28980
rect 34412 28754 34468 28924
rect 34524 28914 34580 28924
rect 34412 28702 34414 28754
rect 34466 28702 34468 28754
rect 34412 28690 34468 28702
rect 34636 28754 34692 28766
rect 34636 28702 34638 28754
rect 34690 28702 34692 28754
rect 34300 28476 34468 28532
rect 33964 28028 34244 28084
rect 33852 27860 33908 27870
rect 33852 27766 33908 27804
rect 33628 27122 33684 27132
rect 33964 26908 34020 28028
rect 34188 27858 34244 27870
rect 34188 27806 34190 27858
rect 34242 27806 34244 27858
rect 34188 27748 34244 27806
rect 34244 27692 34356 27748
rect 34188 27682 34244 27692
rect 33404 26852 33684 26908
rect 33292 26674 33348 26684
rect 33516 26626 33572 26638
rect 33516 26574 33518 26626
rect 33570 26574 33572 26626
rect 32956 26516 33012 26526
rect 33516 26516 33572 26574
rect 33012 26460 33572 26516
rect 33628 26516 33684 26852
rect 33740 26852 34020 26908
rect 33740 26850 33796 26852
rect 33740 26798 33742 26850
rect 33794 26798 33796 26850
rect 33740 26786 33796 26798
rect 34076 26850 34132 26862
rect 34076 26798 34078 26850
rect 34130 26798 34132 26850
rect 33964 26738 34020 26750
rect 33964 26686 33966 26738
rect 34018 26686 34020 26738
rect 33852 26516 33908 26526
rect 33628 26460 33852 26516
rect 32956 26450 33012 26460
rect 33516 26292 33572 26302
rect 32620 22542 32622 22594
rect 32674 22542 32676 22594
rect 32620 22530 32676 22542
rect 32732 24722 32788 24734
rect 32732 24670 32734 24722
rect 32786 24670 32788 24722
rect 32620 22372 32676 22382
rect 32732 22372 32788 24670
rect 32844 24610 32900 25564
rect 32844 24558 32846 24610
rect 32898 24558 32900 24610
rect 32844 23492 32900 24558
rect 33180 25954 33236 25966
rect 33180 25902 33182 25954
rect 33234 25902 33236 25954
rect 33180 24610 33236 25902
rect 33516 25844 33572 26236
rect 33516 25788 33684 25844
rect 33628 25730 33684 25788
rect 33628 25678 33630 25730
rect 33682 25678 33684 25730
rect 33180 24558 33182 24610
rect 33234 24558 33236 24610
rect 33180 23828 33236 24558
rect 33180 23762 33236 23772
rect 33404 25620 33460 25630
rect 33068 23716 33124 23726
rect 33068 23622 33124 23660
rect 33404 23714 33460 25564
rect 33628 25508 33684 25678
rect 33852 25732 33908 26460
rect 33852 25666 33908 25676
rect 33404 23662 33406 23714
rect 33458 23662 33460 23714
rect 33404 23650 33460 23662
rect 33516 25452 33684 25508
rect 33516 24610 33572 25452
rect 33964 25060 34020 26686
rect 33516 24558 33518 24610
rect 33570 24558 33572 24610
rect 32844 23426 32900 23436
rect 33516 23604 33572 24558
rect 33740 25004 34020 25060
rect 33628 24388 33684 24398
rect 33628 23716 33684 24332
rect 33740 23938 33796 25004
rect 33740 23886 33742 23938
rect 33794 23886 33796 23938
rect 33740 23874 33796 23886
rect 33628 23660 33796 23716
rect 33068 22484 33124 22494
rect 33516 22484 33572 23548
rect 33068 22482 33572 22484
rect 33068 22430 33070 22482
rect 33122 22430 33518 22482
rect 33570 22430 33572 22482
rect 33068 22428 33572 22430
rect 33068 22418 33124 22428
rect 32676 22316 32788 22372
rect 32620 22306 32676 22316
rect 32508 20862 32510 20914
rect 32562 20862 32564 20914
rect 32508 20850 32564 20862
rect 32284 20626 32340 20636
rect 32844 20690 32900 20702
rect 32844 20638 32846 20690
rect 32898 20638 32900 20690
rect 31836 20526 31838 20578
rect 31890 20526 31892 20578
rect 31836 20356 31892 20526
rect 31836 20290 31892 20300
rect 32060 20578 32116 20590
rect 32060 20526 32062 20578
rect 32114 20526 32116 20578
rect 32060 19796 32116 20526
rect 32844 20132 32900 20638
rect 33068 20692 33124 20702
rect 33068 20598 33124 20636
rect 33516 20468 33572 22428
rect 33516 20374 33572 20412
rect 33404 20132 33460 20142
rect 32844 20076 33236 20132
rect 33068 19908 33124 19918
rect 32956 19906 33124 19908
rect 32956 19854 33070 19906
rect 33122 19854 33124 19906
rect 32956 19852 33124 19854
rect 32060 19730 32116 19740
rect 32844 19796 32900 19806
rect 31724 19684 31780 19694
rect 31612 19628 31724 19684
rect 31388 18678 31390 18730
rect 31442 18678 31444 18730
rect 30492 17726 30494 17778
rect 30546 17726 30548 17778
rect 30492 17714 30548 17726
rect 30828 17892 30884 17902
rect 30828 17778 30884 17836
rect 30828 17726 30830 17778
rect 30882 17726 30884 17778
rect 30828 17714 30884 17726
rect 30380 17500 30660 17556
rect 30156 16606 30158 16658
rect 30210 16606 30212 16658
rect 30156 16594 30212 16606
rect 30492 16660 30548 16670
rect 30044 15764 30100 15774
rect 29932 15762 30100 15764
rect 29932 15710 30046 15762
rect 30098 15710 30100 15762
rect 29932 15708 30100 15710
rect 29484 15138 29540 15148
rect 29372 14702 29374 14754
rect 29426 14702 29428 14754
rect 29372 14690 29428 14702
rect 29708 14868 29764 14878
rect 29708 14754 29764 14812
rect 29708 14702 29710 14754
rect 29762 14702 29764 14754
rect 29260 13860 29316 14364
rect 29260 13766 29316 13804
rect 29708 13858 29764 14702
rect 29708 13806 29710 13858
rect 29762 13806 29764 13858
rect 29708 13794 29764 13806
rect 30044 14644 30100 15708
rect 30492 14978 30548 16604
rect 30604 16546 30660 17500
rect 31276 16660 31332 16670
rect 31388 16660 31444 18678
rect 31724 18676 31780 19628
rect 32284 19684 32340 19694
rect 32284 19590 32340 19628
rect 31724 18674 32004 18676
rect 31724 18622 31726 18674
rect 31778 18622 32004 18674
rect 31724 18620 32004 18622
rect 31724 18610 31780 18620
rect 30604 16494 30606 16546
rect 30658 16494 30660 16546
rect 30604 15092 30660 16494
rect 30604 15026 30660 15036
rect 31164 16658 31444 16660
rect 31164 16606 31278 16658
rect 31330 16606 31444 16658
rect 31164 16604 31444 16606
rect 30492 14926 30494 14978
rect 30546 14926 30548 14978
rect 30492 14914 30548 14926
rect 30604 14868 30660 14878
rect 30156 14644 30212 14654
rect 30044 14642 30212 14644
rect 30044 14590 30158 14642
rect 30210 14590 30212 14642
rect 30044 14588 30212 14590
rect 28588 13458 28644 13468
rect 28812 13636 28868 13646
rect 28812 13522 28868 13580
rect 30044 13636 30100 14588
rect 30156 14578 30212 14588
rect 30380 14642 30436 14654
rect 30380 14590 30382 14642
rect 30434 14590 30436 14642
rect 30380 13860 30436 14590
rect 30604 14642 30660 14812
rect 30604 14590 30606 14642
rect 30658 14590 30660 14642
rect 30604 14578 30660 14590
rect 30828 14644 30884 14654
rect 31164 14644 31220 16604
rect 31276 16594 31332 16604
rect 31948 16546 32004 18620
rect 32844 18674 32900 19740
rect 32844 18622 32846 18674
rect 32898 18622 32900 18674
rect 32844 18610 32900 18622
rect 31948 16494 31950 16546
rect 32002 16494 32004 16546
rect 31948 16482 32004 16494
rect 31948 15764 32004 15774
rect 31836 15762 32004 15764
rect 31836 15710 31950 15762
rect 32002 15710 32004 15762
rect 31836 15708 32004 15710
rect 31276 15650 31332 15662
rect 31276 15598 31278 15650
rect 31330 15598 31332 15650
rect 31276 15204 31332 15598
rect 31276 15138 31332 15148
rect 30828 14642 31220 14644
rect 30828 14590 30830 14642
rect 30882 14590 31220 14642
rect 30828 14588 31220 14590
rect 31836 15092 31892 15708
rect 31948 15698 32004 15708
rect 30380 13794 30436 13804
rect 30044 13570 30100 13580
rect 28812 13470 28814 13522
rect 28866 13470 28868 13522
rect 28364 12898 28420 12908
rect 28252 11454 28254 11506
rect 28306 11454 28308 11506
rect 27804 10946 27972 10948
rect 27804 10894 27806 10946
rect 27858 10894 27972 10946
rect 27804 10892 27972 10894
rect 28140 11394 28196 11406
rect 28140 11342 28142 11394
rect 28194 11342 28196 11394
rect 27804 10882 27860 10892
rect 28140 10724 28196 11342
rect 28140 10630 28196 10668
rect 28252 10500 28308 11454
rect 28700 11506 28756 11518
rect 28700 11454 28702 11506
rect 28754 11454 28756 11506
rect 28700 11282 28756 11454
rect 28812 11508 28868 13470
rect 30156 13524 30212 13534
rect 30156 13430 30212 13468
rect 30828 13524 30884 14588
rect 31836 14532 31892 15036
rect 31836 14466 31892 14476
rect 32284 15204 32340 15214
rect 32956 15148 33012 19852
rect 33068 19842 33124 19852
rect 33180 18898 33236 20076
rect 33404 19794 33460 20076
rect 33740 19906 33796 23660
rect 33964 22820 34020 22830
rect 33964 22726 34020 22764
rect 34076 22372 34132 26798
rect 34188 26628 34244 26638
rect 34188 26534 34244 26572
rect 34300 26626 34356 27692
rect 34300 26574 34302 26626
rect 34354 26574 34356 26626
rect 34300 26562 34356 26574
rect 34412 26180 34468 28476
rect 34636 28084 34692 28702
rect 34636 28018 34692 28028
rect 34524 27970 34580 27982
rect 34524 27918 34526 27970
rect 34578 27918 34580 27970
rect 34524 27860 34580 27918
rect 34524 27410 34580 27804
rect 34860 27748 34916 29484
rect 34972 28420 35028 33852
rect 35196 33794 35252 33964
rect 35868 34020 35924 34030
rect 35868 33906 35924 33964
rect 35868 33854 35870 33906
rect 35922 33854 35924 33906
rect 35868 33842 35924 33854
rect 36204 33906 36260 35756
rect 36764 35812 36820 35822
rect 36764 35718 36820 35756
rect 36876 35252 36932 36092
rect 37324 35812 37380 35822
rect 37324 35718 37380 35756
rect 36876 35196 37156 35252
rect 37100 34802 37156 35196
rect 37100 34750 37102 34802
rect 37154 34750 37156 34802
rect 37100 34738 37156 34750
rect 36204 33854 36206 33906
rect 36258 33854 36260 33906
rect 36204 33842 36260 33854
rect 36540 34018 36596 34030
rect 36540 33966 36542 34018
rect 36594 33966 36596 34018
rect 35196 33742 35198 33794
rect 35250 33742 35252 33794
rect 35196 33730 35252 33742
rect 35644 33796 35700 33806
rect 35532 33684 35588 33694
rect 35532 33590 35588 33628
rect 35196 33292 35460 33302
rect 35252 33236 35300 33292
rect 35356 33236 35404 33292
rect 35196 33226 35460 33236
rect 35196 33122 35252 33134
rect 35196 33070 35198 33122
rect 35250 33070 35252 33122
rect 35196 32898 35252 33070
rect 35196 32846 35198 32898
rect 35250 32846 35252 32898
rect 35196 32834 35252 32846
rect 35644 31892 35700 33740
rect 35756 33460 35812 33470
rect 35756 32898 35812 33404
rect 35756 32846 35758 32898
rect 35810 32846 35812 32898
rect 35756 32834 35812 32846
rect 35644 31826 35700 31836
rect 35756 31890 35812 31902
rect 35756 31838 35758 31890
rect 35810 31838 35812 31890
rect 35532 31780 35588 31790
rect 35196 31276 35460 31286
rect 35252 31220 35300 31276
rect 35356 31220 35404 31276
rect 35196 31210 35460 31220
rect 35532 30884 35588 31724
rect 35756 31780 35812 31838
rect 35756 31714 35812 31724
rect 36316 31778 36372 31790
rect 36316 31726 36318 31778
rect 36370 31726 36372 31778
rect 36316 30994 36372 31726
rect 36540 31444 36596 33966
rect 36988 34020 37044 34030
rect 37436 34020 37492 36876
rect 37548 34916 37604 38892
rect 37660 38946 37716 39116
rect 37660 38894 37662 38946
rect 37714 38894 37716 38946
rect 37660 38052 37716 38894
rect 37772 39058 37828 39070
rect 37772 39006 37774 39058
rect 37826 39006 37828 39058
rect 37772 38276 37828 39006
rect 37884 38724 37940 39676
rect 38108 38948 38164 40460
rect 38444 40180 38500 40908
rect 38668 40850 38724 40908
rect 38668 40798 38670 40850
rect 38722 40798 38724 40850
rect 38668 40786 38724 40798
rect 38780 41580 38892 41636
rect 38332 40124 38500 40180
rect 38556 40740 38612 40750
rect 38556 40180 38612 40684
rect 38556 40124 38668 40180
rect 38332 39954 38388 40124
rect 38612 39956 38668 40124
rect 38332 39902 38334 39954
rect 38386 39902 38388 39954
rect 38108 38854 38164 38892
rect 38220 39732 38276 39742
rect 37884 38658 37940 38668
rect 37772 38210 37828 38220
rect 37884 38052 37940 38062
rect 37660 37996 37884 38052
rect 37660 36706 37716 36718
rect 37660 36654 37662 36706
rect 37714 36654 37716 36706
rect 37660 36596 37716 36654
rect 37660 36530 37716 36540
rect 37548 34850 37604 34860
rect 37660 34804 37716 34814
rect 37660 34690 37716 34748
rect 37660 34638 37662 34690
rect 37714 34638 37716 34690
rect 37660 34626 37716 34638
rect 37884 34802 37940 37996
rect 37996 36932 38052 36942
rect 38220 36932 38276 39676
rect 38332 39170 38388 39902
rect 38332 39118 38334 39170
rect 38386 39118 38388 39170
rect 38332 39106 38388 39118
rect 38556 39900 38668 39956
rect 38556 38946 38612 39900
rect 38556 38894 38558 38946
rect 38610 38894 38612 38946
rect 38556 38882 38612 38894
rect 37996 36930 38276 36932
rect 37996 36878 37998 36930
rect 38050 36878 38276 36930
rect 37996 36876 38276 36878
rect 38556 38276 38612 38286
rect 37996 36866 38052 36876
rect 38332 36708 38388 36718
rect 37996 36706 38388 36708
rect 37996 36654 38334 36706
rect 38386 36654 38388 36706
rect 37996 36652 38388 36654
rect 37996 36146 38052 36652
rect 38332 36642 38388 36652
rect 37996 36094 37998 36146
rect 38050 36094 38052 36146
rect 37996 36082 38052 36094
rect 37884 34750 37886 34802
rect 37938 34750 37940 34802
rect 37884 34692 37940 34750
rect 37940 34636 38052 34692
rect 37884 34626 37940 34636
rect 37548 34020 37604 34030
rect 37044 34018 37940 34020
rect 37044 33966 37550 34018
rect 37602 33966 37940 34018
rect 37044 33964 37940 33966
rect 36988 33926 37044 33964
rect 37548 33954 37604 33964
rect 37324 33012 37380 33022
rect 37324 32898 37380 32956
rect 37324 32846 37326 32898
rect 37378 32846 37380 32898
rect 37324 32834 37380 32846
rect 37884 32786 37940 33964
rect 37996 33460 38052 34636
rect 37996 33394 38052 33404
rect 37884 32734 37886 32786
rect 37938 32734 37940 32786
rect 37884 32722 37940 32734
rect 38108 33012 38164 33022
rect 38108 32786 38164 32956
rect 38108 32734 38110 32786
rect 38162 32734 38164 32786
rect 38108 32722 38164 32734
rect 38444 32450 38500 32462
rect 38444 32398 38446 32450
rect 38498 32398 38500 32450
rect 37772 31892 37828 31902
rect 37548 31836 37772 31892
rect 36540 31378 36596 31388
rect 36652 31778 36708 31790
rect 36652 31726 36654 31778
rect 36706 31726 36708 31778
rect 36316 30942 36318 30994
rect 36370 30942 36372 30994
rect 36316 30930 36372 30942
rect 35084 30882 35588 30884
rect 35084 30830 35534 30882
rect 35586 30830 35588 30882
rect 35084 30828 35588 30830
rect 35084 28868 35140 30828
rect 35532 30548 35588 30828
rect 35532 30482 35588 30492
rect 35644 30770 35700 30782
rect 35644 30718 35646 30770
rect 35698 30718 35700 30770
rect 35532 30100 35588 30110
rect 35420 29764 35476 29774
rect 35420 29670 35476 29708
rect 35532 29762 35588 30044
rect 35532 29710 35534 29762
rect 35586 29710 35588 29762
rect 35196 29540 35252 29550
rect 35196 29446 35252 29484
rect 35196 29260 35460 29270
rect 35252 29204 35300 29260
rect 35356 29204 35404 29260
rect 35196 29194 35460 29204
rect 35196 28868 35252 28878
rect 35084 28866 35252 28868
rect 35084 28814 35198 28866
rect 35250 28814 35252 28866
rect 35084 28812 35252 28814
rect 35196 28802 35252 28812
rect 35532 28420 35588 29710
rect 35644 28978 35700 30718
rect 35756 30772 35812 30782
rect 35756 29874 35812 30716
rect 35756 29822 35758 29874
rect 35810 29822 35812 29874
rect 35756 29810 35812 29822
rect 35980 30324 36036 30334
rect 35644 28926 35646 28978
rect 35698 28926 35700 28978
rect 35644 28866 35700 28926
rect 35644 28814 35646 28866
rect 35698 28814 35700 28866
rect 35644 28802 35700 28814
rect 34972 28364 35140 28420
rect 35532 28364 35700 28420
rect 35084 27972 35140 28364
rect 34524 27358 34526 27410
rect 34578 27358 34580 27410
rect 34524 27346 34580 27358
rect 34636 27692 34916 27748
rect 34972 27916 35140 27972
rect 35196 28196 35252 28206
rect 35196 27970 35252 28140
rect 35532 28084 35588 28094
rect 35532 27990 35588 28028
rect 35196 27918 35198 27970
rect 35250 27918 35252 27970
rect 34300 26124 34468 26180
rect 34188 23828 34244 23838
rect 34188 23734 34244 23772
rect 33964 22316 34132 22372
rect 33964 20802 34020 22316
rect 34300 21812 34356 26124
rect 34412 25956 34468 25966
rect 34412 25862 34468 25900
rect 34636 23828 34692 27692
rect 34748 27410 34804 27422
rect 34748 27358 34750 27410
rect 34802 27358 34804 27410
rect 34748 26626 34804 27358
rect 34972 26908 35028 27916
rect 35196 27906 35252 27918
rect 35084 27748 35140 27758
rect 35084 27654 35140 27692
rect 35308 27748 35364 27758
rect 35644 27748 35700 28364
rect 35308 27746 35588 27748
rect 35308 27694 35310 27746
rect 35362 27694 35588 27746
rect 35308 27692 35588 27694
rect 35308 27682 35364 27692
rect 34860 26852 35028 26908
rect 35084 27524 35140 27534
rect 34860 26850 34916 26852
rect 34860 26798 34862 26850
rect 34914 26798 34916 26850
rect 34860 26786 34916 26798
rect 34748 26574 34750 26626
rect 34802 26574 34804 26626
rect 34748 24612 34804 26574
rect 34972 26738 35028 26750
rect 34972 26686 34974 26738
rect 35026 26686 35028 26738
rect 34972 26626 35028 26686
rect 34972 26574 34974 26626
rect 35026 26574 35028 26626
rect 34972 26562 35028 26574
rect 35084 26402 35140 27468
rect 35196 27244 35460 27254
rect 35252 27188 35300 27244
rect 35356 27188 35404 27244
rect 35196 27178 35460 27188
rect 35532 26852 35588 27692
rect 35644 27654 35700 27692
rect 35868 27746 35924 27758
rect 35868 27694 35870 27746
rect 35922 27694 35924 27746
rect 35532 26786 35588 26796
rect 35868 26740 35924 27694
rect 35868 26674 35924 26684
rect 35532 26626 35588 26638
rect 35532 26574 35534 26626
rect 35586 26574 35588 26626
rect 35196 26516 35252 26526
rect 35196 26422 35252 26460
rect 35084 26350 35086 26402
rect 35138 26350 35140 26402
rect 35084 26338 35140 26350
rect 35532 25956 35588 26574
rect 35868 26516 35924 26526
rect 35868 26422 35924 26460
rect 35980 26516 36036 30268
rect 36652 30324 36708 31726
rect 36988 31780 37044 31790
rect 36988 31686 37044 31724
rect 37324 31778 37380 31790
rect 37324 31726 37326 31778
rect 37378 31726 37380 31778
rect 37324 30772 37380 31726
rect 37324 30706 37380 30716
rect 36988 30660 37044 30670
rect 36988 30658 37268 30660
rect 36988 30606 36990 30658
rect 37042 30606 37268 30658
rect 36988 30604 37268 30606
rect 36988 30594 37044 30604
rect 36652 30258 36708 30268
rect 36540 30212 36596 30222
rect 36540 29988 36596 30156
rect 36652 29988 36708 29998
rect 36540 29986 36708 29988
rect 36540 29934 36654 29986
rect 36706 29934 36708 29986
rect 36540 29932 36708 29934
rect 36652 29922 36708 29932
rect 36204 29876 36260 29886
rect 36204 29782 36260 29820
rect 36988 29876 37044 29886
rect 36092 28980 36148 28990
rect 36092 28866 36148 28924
rect 36092 28814 36094 28866
rect 36146 28814 36148 28866
rect 36092 28802 36148 28814
rect 36428 28978 36484 28990
rect 36428 28926 36430 28978
rect 36482 28926 36484 28978
rect 35980 26514 36148 26516
rect 35980 26462 35982 26514
rect 36034 26462 36148 26514
rect 35980 26460 36148 26462
rect 35980 26450 36036 26460
rect 35532 25890 35588 25900
rect 35420 25842 35476 25854
rect 35420 25790 35422 25842
rect 35474 25790 35476 25842
rect 34972 25620 35028 25658
rect 34972 25554 35028 25564
rect 34972 25396 35028 25406
rect 35420 25396 35476 25790
rect 35868 25730 35924 25742
rect 35868 25678 35870 25730
rect 35922 25678 35924 25730
rect 35644 25620 35700 25630
rect 35420 25340 35588 25396
rect 34972 24946 35028 25340
rect 35196 25228 35460 25238
rect 35252 25172 35300 25228
rect 35356 25172 35404 25228
rect 35196 25162 35460 25172
rect 34972 24894 34974 24946
rect 35026 24894 35028 24946
rect 34972 24882 35028 24894
rect 34748 24546 34804 24556
rect 35532 24500 35588 25340
rect 35532 24406 35588 24444
rect 34636 23772 34804 23828
rect 34636 23604 34692 23614
rect 34636 23510 34692 23548
rect 34412 21812 34468 21822
rect 34300 21756 34412 21812
rect 34412 21718 34468 21756
rect 34076 21588 34132 21598
rect 34076 21494 34132 21532
rect 34748 20916 34804 23772
rect 35532 23604 35588 23614
rect 35644 23604 35700 25564
rect 35868 25508 35924 25678
rect 35868 25442 35924 25452
rect 36092 25508 36148 26460
rect 36428 26514 36484 28926
rect 36988 28868 37044 29820
rect 37100 29652 37156 29662
rect 37100 29558 37156 29596
rect 37212 29540 37268 30604
rect 37324 30548 37380 30558
rect 37548 30548 37604 31836
rect 37772 31798 37828 31836
rect 38444 31890 38500 32398
rect 38444 31838 38446 31890
rect 38498 31838 38500 31890
rect 38444 31826 38500 31838
rect 37660 31444 37716 31454
rect 37660 30772 37716 31388
rect 37660 30770 37940 30772
rect 37660 30718 37662 30770
rect 37714 30718 37940 30770
rect 37660 30716 37940 30718
rect 37660 30706 37716 30716
rect 37324 30546 37604 30548
rect 37324 30494 37326 30546
rect 37378 30494 37604 30546
rect 37324 30492 37604 30494
rect 37324 30482 37380 30492
rect 37884 29988 37940 30716
rect 38444 30548 38500 30558
rect 37996 30434 38052 30446
rect 37996 30382 37998 30434
rect 38050 30382 38052 30434
rect 37996 30324 38052 30382
rect 37996 30258 38052 30268
rect 37996 29988 38052 29998
rect 37884 29986 38052 29988
rect 37884 29934 37998 29986
rect 38050 29934 38052 29986
rect 37884 29932 38052 29934
rect 37996 29922 38052 29932
rect 38444 29986 38500 30492
rect 38444 29934 38446 29986
rect 38498 29934 38500 29986
rect 37212 29474 37268 29484
rect 37548 29650 37604 29662
rect 37548 29598 37550 29650
rect 37602 29598 37604 29650
rect 37548 29540 37604 29598
rect 37548 29474 37604 29484
rect 37100 28868 37156 28878
rect 36988 28866 37156 28868
rect 36988 28814 37102 28866
rect 37154 28814 37156 28866
rect 36988 28812 37156 28814
rect 37100 28802 37156 28812
rect 38332 28644 38388 28654
rect 37100 26852 37156 26862
rect 37100 26850 37940 26852
rect 37100 26798 37102 26850
rect 37154 26798 37940 26850
rect 37100 26796 37940 26798
rect 37100 26786 37156 26796
rect 36428 26462 36430 26514
rect 36482 26462 36484 26514
rect 36092 25442 36148 25452
rect 36204 25730 36260 25742
rect 36204 25678 36206 25730
rect 36258 25678 36260 25730
rect 36204 25396 36260 25678
rect 36428 25732 36484 26462
rect 36540 26628 36596 26638
rect 36540 25954 36596 26572
rect 37660 26628 37716 26638
rect 37548 26516 37604 26526
rect 37436 26514 37604 26516
rect 37436 26462 37550 26514
rect 37602 26462 37604 26514
rect 37436 26460 37604 26462
rect 36540 25902 36542 25954
rect 36594 25902 36596 25954
rect 36540 25890 36596 25902
rect 36988 26402 37044 26414
rect 36988 26350 36990 26402
rect 37042 26350 37044 26402
rect 36988 25954 37044 26350
rect 36988 25902 36990 25954
rect 37042 25902 37044 25954
rect 36988 25890 37044 25902
rect 36428 25666 36484 25676
rect 36876 25732 36932 25742
rect 36204 25330 36260 25340
rect 36428 24836 36484 24846
rect 36652 24836 36708 24846
rect 36204 24834 36652 24836
rect 36204 24782 36430 24834
rect 36482 24782 36652 24834
rect 36204 24780 36652 24782
rect 35980 24500 36036 24510
rect 35980 24406 36036 24444
rect 35588 23548 35700 23604
rect 35532 23538 35588 23548
rect 35196 23212 35460 23222
rect 35252 23156 35300 23212
rect 35356 23156 35404 23212
rect 35196 23146 35460 23156
rect 35532 22820 35588 22830
rect 34972 21812 35028 21822
rect 34972 21718 35028 21756
rect 33964 20750 33966 20802
rect 34018 20750 34020 20802
rect 33740 19854 33742 19906
rect 33794 19854 33796 19906
rect 33740 19842 33796 19854
rect 33852 20356 33908 20366
rect 33404 19742 33406 19794
rect 33458 19742 33460 19794
rect 33404 19730 33460 19742
rect 33180 18846 33182 18898
rect 33234 18846 33236 18898
rect 33180 18834 33236 18846
rect 33852 18562 33908 20300
rect 33964 20132 34020 20750
rect 34636 20860 34804 20916
rect 35084 21476 35140 21486
rect 33964 20066 34020 20076
rect 34300 20692 34356 20702
rect 34300 19908 34356 20636
rect 34412 19908 34468 19918
rect 34300 19906 34468 19908
rect 34300 19854 34414 19906
rect 34466 19854 34468 19906
rect 34300 19852 34468 19854
rect 34412 19842 34468 19852
rect 33852 18510 33854 18562
rect 33906 18510 33908 18562
rect 33852 18498 33908 18510
rect 34076 19794 34132 19806
rect 34076 19742 34078 19794
rect 34130 19742 34132 19794
rect 34076 18228 34132 19742
rect 34636 18564 34692 20860
rect 34972 20804 35028 20814
rect 35084 20804 35140 21420
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 21028 35252 21038
rect 35196 20934 35252 20972
rect 34748 20802 35140 20804
rect 34748 20750 34974 20802
rect 35026 20750 35140 20802
rect 34748 20748 35140 20750
rect 34748 19794 34804 20748
rect 34972 20738 35028 20748
rect 35196 20356 35252 20366
rect 35196 19906 35252 20300
rect 35196 19854 35198 19906
rect 35250 19854 35252 19906
rect 35196 19842 35252 19854
rect 34748 19742 34750 19794
rect 34802 19742 34804 19794
rect 34748 19730 34804 19742
rect 35196 19180 35460 19190
rect 35252 19124 35300 19180
rect 35356 19124 35404 19180
rect 35196 19114 35460 19124
rect 35532 18786 35588 22764
rect 36204 22820 36260 24780
rect 36428 24770 36484 24780
rect 36652 24770 36708 24780
rect 36876 24500 36932 25676
rect 37436 25620 37492 26460
rect 37548 26450 37604 26460
rect 37548 25732 37604 25770
rect 37548 25666 37604 25676
rect 37436 25554 37492 25564
rect 37548 25508 37604 25518
rect 37660 25508 37716 26572
rect 37772 25730 37828 25742
rect 37772 25678 37774 25730
rect 37826 25678 37828 25730
rect 37772 25620 37828 25678
rect 37772 25554 37828 25564
rect 37884 25730 37940 26796
rect 38220 26740 38276 26750
rect 37884 25678 37886 25730
rect 37938 25678 37940 25730
rect 37604 25452 37716 25508
rect 37324 24500 37380 24510
rect 36204 22726 36260 22764
rect 36428 23604 36484 23614
rect 35756 22484 35812 22494
rect 36428 22484 36484 23548
rect 35756 22482 36484 22484
rect 35756 22430 35758 22482
rect 35810 22430 36484 22482
rect 35756 22428 36484 22430
rect 36876 23602 36932 24444
rect 37212 24498 37380 24500
rect 37212 24446 37326 24498
rect 37378 24446 37380 24498
rect 37212 24444 37380 24446
rect 37212 23826 37268 24444
rect 37324 24434 37380 24444
rect 37212 23774 37214 23826
rect 37266 23774 37268 23826
rect 37212 23762 37268 23774
rect 37548 23826 37604 25452
rect 37884 24836 37940 25678
rect 37996 26514 38052 26526
rect 37996 26462 37998 26514
rect 38050 26462 38052 26514
rect 37996 26292 38052 26462
rect 37996 25732 38052 26236
rect 37996 25666 38052 25676
rect 38108 26402 38164 26414
rect 38108 26350 38110 26402
rect 38162 26350 38164 26402
rect 38108 25730 38164 26350
rect 38108 25678 38110 25730
rect 38162 25678 38164 25730
rect 37884 24724 37940 24780
rect 37996 24724 38052 24734
rect 37884 24722 38052 24724
rect 37884 24670 37998 24722
rect 38050 24670 38052 24722
rect 37884 24668 38052 24670
rect 37548 23774 37550 23826
rect 37602 23774 37604 23826
rect 37548 23762 37604 23774
rect 37884 23716 37940 23726
rect 36876 23550 36878 23602
rect 36930 23550 36932 23602
rect 35756 22418 35812 22428
rect 35980 21924 36036 22428
rect 35980 21858 36036 21868
rect 35644 21812 35700 21822
rect 35868 21812 35924 21822
rect 35700 21810 35924 21812
rect 35700 21758 35870 21810
rect 35922 21758 35924 21810
rect 35700 21756 35924 21758
rect 35644 21718 35700 21756
rect 35868 21746 35924 21756
rect 36652 21586 36708 21598
rect 36652 21534 36654 21586
rect 36706 21534 36708 21586
rect 36204 21476 36260 21486
rect 36204 21382 36260 21420
rect 36652 21474 36708 21534
rect 36652 21422 36654 21474
rect 36706 21422 36708 21474
rect 36652 21410 36708 21422
rect 36876 21474 36932 23550
rect 37660 23714 37940 23716
rect 37660 23662 37886 23714
rect 37938 23662 37940 23714
rect 37660 23660 37940 23662
rect 37660 23156 37716 23660
rect 37884 23650 37940 23660
rect 37324 23100 37716 23156
rect 37324 23042 37380 23100
rect 37324 22990 37326 23042
rect 37378 22990 37380 23042
rect 37324 22978 37380 22990
rect 37884 22708 37940 22718
rect 37996 22708 38052 24668
rect 37884 22706 38052 22708
rect 37884 22654 37886 22706
rect 37938 22654 38052 22706
rect 37884 22652 38052 22654
rect 37884 22642 37940 22652
rect 37996 22596 38052 22652
rect 37996 22530 38052 22540
rect 36876 21422 36878 21474
rect 36930 21422 36932 21474
rect 36876 21410 36932 21422
rect 37100 21812 37156 21822
rect 38108 21812 38164 25678
rect 38220 23938 38276 26684
rect 38220 23886 38222 23938
rect 38274 23886 38276 23938
rect 38220 23874 38276 23886
rect 38220 21812 38276 21822
rect 38108 21810 38276 21812
rect 38108 21758 38222 21810
rect 38274 21758 38276 21810
rect 38108 21756 38276 21758
rect 37100 21586 37156 21756
rect 37100 21534 37102 21586
rect 37154 21534 37156 21586
rect 36316 20804 36372 20814
rect 36316 20710 36372 20748
rect 35644 20578 35700 20590
rect 35644 20526 35646 20578
rect 35698 20526 35700 20578
rect 35644 19348 35700 20526
rect 36204 20578 36260 20590
rect 36204 20526 36206 20578
rect 36258 20526 36260 20578
rect 35644 19282 35700 19292
rect 35980 19682 36036 19694
rect 35980 19630 35982 19682
rect 36034 19630 36036 19682
rect 35980 18898 36036 19630
rect 35980 18846 35982 18898
rect 36034 18846 36036 18898
rect 35980 18834 36036 18846
rect 35532 18734 35534 18786
rect 35586 18734 35588 18786
rect 35532 18722 35588 18734
rect 35980 18676 36036 18686
rect 35980 18582 36036 18620
rect 34748 18564 34804 18574
rect 34636 18562 34804 18564
rect 34636 18510 34750 18562
rect 34802 18510 34804 18562
rect 34636 18508 34804 18510
rect 34748 18452 34804 18508
rect 36204 18564 36260 20526
rect 37100 20468 37156 21534
rect 37548 21586 37604 21598
rect 37548 21534 37550 21586
rect 37602 21534 37604 21586
rect 37548 21474 37604 21534
rect 37548 21422 37550 21474
rect 37602 21422 37604 21474
rect 37212 20804 37268 20814
rect 37212 20710 37268 20748
rect 37548 20690 37604 21422
rect 38220 21474 38276 21756
rect 38220 21422 38222 21474
rect 38274 21422 38276 21474
rect 38220 21410 38276 21422
rect 38332 20804 38388 28588
rect 38444 28082 38500 29934
rect 38556 28644 38612 38220
rect 38780 38050 38836 41580
rect 38892 41570 38948 41580
rect 39788 41692 39900 41748
rect 39228 39060 39284 39070
rect 39228 38966 39284 39004
rect 38892 38724 38948 38734
rect 39788 38668 39844 41692
rect 39900 41654 39956 41692
rect 40460 41746 40516 41758
rect 40460 41694 40462 41746
rect 40514 41694 40516 41746
rect 40348 40964 40404 40974
rect 39900 40068 39956 40078
rect 39900 39974 39956 40012
rect 40348 38724 40404 40908
rect 40460 39060 40516 41694
rect 40460 38994 40516 39004
rect 40460 38724 40516 38734
rect 40348 38722 40516 38724
rect 40348 38670 40462 38722
rect 40514 38670 40516 38722
rect 40348 38668 40516 38670
rect 38892 38630 38948 38668
rect 39676 38612 39844 38668
rect 38780 37998 38782 38050
rect 38834 37998 38836 38050
rect 38780 37986 38836 37998
rect 39228 38162 39284 38174
rect 39228 38110 39230 38162
rect 39282 38110 39284 38162
rect 39228 37714 39284 38110
rect 39228 37662 39230 37714
rect 39282 37662 39284 37714
rect 38668 36706 38724 36718
rect 39004 36708 39060 36718
rect 38668 36654 38670 36706
rect 38722 36654 38724 36706
rect 38668 33684 38724 36654
rect 38780 36706 39060 36708
rect 38780 36654 39006 36706
rect 39058 36654 39060 36706
rect 38780 36652 39060 36654
rect 38780 34914 38836 36652
rect 39004 36642 39060 36652
rect 38892 36036 38948 36046
rect 38892 35810 38948 35980
rect 38892 35758 38894 35810
rect 38946 35758 38948 35810
rect 38892 35746 38948 35758
rect 39228 35812 39284 37662
rect 39676 37714 39732 38612
rect 39788 38610 39844 38612
rect 39788 38558 39790 38610
rect 39842 38558 39844 38610
rect 39788 38546 39844 38558
rect 40236 38612 40404 38668
rect 40460 38658 40516 38668
rect 39788 38164 39844 38174
rect 40236 38164 40292 38612
rect 39788 38162 40292 38164
rect 39788 38110 39790 38162
rect 39842 38110 40292 38162
rect 39788 38108 40292 38110
rect 39788 38098 39844 38108
rect 40348 38052 40404 38062
rect 39676 37662 39678 37714
rect 39730 37662 39732 37714
rect 38780 34862 38782 34914
rect 38834 34862 38836 34914
rect 38780 34850 38836 34862
rect 38780 34132 38836 34142
rect 38780 34018 38836 34076
rect 38780 33966 38782 34018
rect 38834 33966 38836 34018
rect 38780 33954 38836 33966
rect 39228 34020 39284 35756
rect 38668 33618 38724 33628
rect 39116 33460 39172 33470
rect 39116 32900 39172 33404
rect 39228 33012 39284 33964
rect 39340 36594 39396 36606
rect 39340 36542 39342 36594
rect 39394 36542 39396 36594
rect 39340 33572 39396 36542
rect 39676 36036 39732 37662
rect 39788 37828 39844 37838
rect 39788 36146 39844 37772
rect 40348 37714 40404 37996
rect 40348 37662 40350 37714
rect 40402 37662 40404 37714
rect 40348 37604 40404 37662
rect 40348 37538 40404 37548
rect 40796 36820 40852 42588
rect 41132 41972 41188 42702
rect 41132 41906 41188 41916
rect 40908 41860 40964 41870
rect 40908 41766 40964 41804
rect 41580 41636 41636 41646
rect 41356 41524 41412 41534
rect 41356 41522 41524 41524
rect 41356 41470 41358 41522
rect 41410 41470 41524 41522
rect 41356 41468 41524 41470
rect 41356 41458 41412 41468
rect 41244 40740 41300 40750
rect 41244 40646 41300 40684
rect 40908 40068 40964 40078
rect 40908 39954 40964 40012
rect 40908 39902 40910 39954
rect 40962 39902 40964 39954
rect 40908 39890 40964 39902
rect 41468 39956 41524 41468
rect 41580 40850 41636 41580
rect 41580 40798 41582 40850
rect 41634 40798 41636 40850
rect 41580 40786 41636 40798
rect 41916 40068 41972 43822
rect 42364 42756 42420 45612
rect 42924 45332 42980 46622
rect 42924 45266 42980 45276
rect 43036 46564 43092 46574
rect 43036 43986 43092 46508
rect 43036 43934 43038 43986
rect 43090 43934 43092 43986
rect 43036 43922 43092 43934
rect 43148 45666 43204 45678
rect 43148 45614 43150 45666
rect 43202 45614 43204 45666
rect 42476 43874 42532 43886
rect 42476 43822 42478 43874
rect 42530 43822 42532 43874
rect 42476 43708 42532 43822
rect 43148 43764 43204 45614
rect 43708 44100 43764 44110
rect 43820 44100 43876 48636
rect 44156 48626 44212 48636
rect 50556 48412 50820 48422
rect 50612 48356 50660 48412
rect 50716 48356 50764 48412
rect 50556 48346 50820 48356
rect 44044 46564 44100 46574
rect 44044 46470 44100 46508
rect 50556 46396 50820 46406
rect 50612 46340 50660 46396
rect 50716 46340 50764 46396
rect 50556 46330 50820 46340
rect 46060 45890 46116 45902
rect 46060 45838 46062 45890
rect 46114 45838 46116 45890
rect 45612 44884 45668 44894
rect 45388 44882 45668 44884
rect 45388 44830 45614 44882
rect 45666 44830 45668 44882
rect 45388 44828 45668 44830
rect 45164 44660 45220 44670
rect 45164 44566 45220 44604
rect 43708 44098 43876 44100
rect 43708 44046 43710 44098
rect 43762 44046 43876 44098
rect 43708 44044 43876 44046
rect 45388 44098 45444 44828
rect 45612 44818 45668 44828
rect 45388 44046 45390 44098
rect 45442 44046 45444 44098
rect 43708 44034 43764 44044
rect 42476 43652 42644 43708
rect 42476 42756 42532 42766
rect 42364 42754 42532 42756
rect 42364 42702 42478 42754
rect 42530 42702 42532 42754
rect 42364 42700 42532 42702
rect 42476 42690 42532 42700
rect 42588 41972 42644 43652
rect 42588 41074 42644 41916
rect 42588 41022 42590 41074
rect 42642 41022 42644 41074
rect 41692 40012 41972 40068
rect 42364 40626 42420 40638
rect 42364 40574 42366 40626
rect 42418 40574 42420 40626
rect 42364 40068 42420 40574
rect 41580 39956 41636 39966
rect 41468 39954 41636 39956
rect 41468 39902 41582 39954
rect 41634 39902 41636 39954
rect 41468 39900 41636 39902
rect 41580 39890 41636 39900
rect 41244 39844 41300 39854
rect 41244 39842 41412 39844
rect 41244 39790 41246 39842
rect 41298 39790 41412 39842
rect 41244 39788 41412 39790
rect 41244 39778 41300 39788
rect 41356 39060 41412 39788
rect 41132 38948 41188 38958
rect 41132 38722 41188 38892
rect 41132 38670 41134 38722
rect 41186 38670 41188 38722
rect 41132 38658 41188 38670
rect 41244 38724 41300 38734
rect 41244 37938 41300 38668
rect 41244 37886 41246 37938
rect 41298 37886 41300 37938
rect 41244 37874 41300 37886
rect 40908 37828 40964 37838
rect 40908 37734 40964 37772
rect 40796 36764 40964 36820
rect 39788 36094 39790 36146
rect 39842 36094 39844 36146
rect 39788 36082 39844 36094
rect 39900 36706 39956 36718
rect 39900 36654 39902 36706
rect 39954 36654 39956 36706
rect 39340 33506 39396 33516
rect 39452 34916 39508 34926
rect 39452 34690 39508 34860
rect 39452 34638 39454 34690
rect 39506 34638 39508 34690
rect 39228 32946 39284 32956
rect 39116 32806 39172 32844
rect 39228 32676 39284 32686
rect 39116 31890 39172 31902
rect 39116 31838 39118 31890
rect 39170 31838 39172 31890
rect 39116 30546 39172 31838
rect 39116 30494 39118 30546
rect 39170 30494 39172 30546
rect 39116 30482 39172 30494
rect 39228 30772 39284 32620
rect 39228 30658 39284 30716
rect 39228 30606 39230 30658
rect 39282 30606 39284 30658
rect 39228 30324 39284 30606
rect 38892 30268 39284 30324
rect 38892 29986 38948 30268
rect 39452 30100 39508 34638
rect 39676 34018 39732 35980
rect 39676 33966 39678 34018
rect 39730 33966 39732 34018
rect 39676 32676 39732 33966
rect 39676 32610 39732 32620
rect 39900 31892 39956 36654
rect 40460 36708 40516 36718
rect 40460 36706 40852 36708
rect 40460 36654 40462 36706
rect 40514 36654 40852 36706
rect 40460 36652 40852 36654
rect 40460 36642 40516 36652
rect 40348 36148 40404 36158
rect 40348 35700 40404 36092
rect 40796 36034 40852 36652
rect 40796 35982 40798 36034
rect 40850 35982 40852 36034
rect 40796 35970 40852 35982
rect 40124 34802 40180 34814
rect 40124 34750 40126 34802
rect 40178 34750 40180 34802
rect 40124 34020 40180 34750
rect 40348 34244 40404 35644
rect 40796 34692 40852 34702
rect 40796 34578 40852 34636
rect 40796 34526 40798 34578
rect 40850 34526 40852 34578
rect 40796 34514 40852 34526
rect 40572 34244 40628 34254
rect 40348 34178 40404 34188
rect 40460 34188 40572 34244
rect 40348 34020 40404 34030
rect 40124 33964 40348 34020
rect 40236 32786 40292 33964
rect 40348 33926 40404 33964
rect 40236 32734 40238 32786
rect 40290 32734 40292 32786
rect 40124 32676 40180 32686
rect 40124 32582 40180 32620
rect 40236 31948 40292 32734
rect 39900 31826 39956 31836
rect 40012 31892 40292 31948
rect 39900 31668 39956 31678
rect 40012 31668 40068 31892
rect 40236 31816 40292 31836
rect 39676 31666 40068 31668
rect 39676 31614 39902 31666
rect 39954 31614 40068 31666
rect 39676 31612 40068 31614
rect 40348 31668 40404 31678
rect 39676 30770 39732 31612
rect 39900 31602 39956 31612
rect 40348 31332 40404 31612
rect 40348 31266 40404 31276
rect 39676 30718 39678 30770
rect 39730 30718 39732 30770
rect 39676 30548 39732 30718
rect 39676 30482 39732 30492
rect 39900 30772 39956 30782
rect 39452 30034 39508 30044
rect 38892 29934 38894 29986
rect 38946 29934 38948 29986
rect 38892 29922 38948 29934
rect 39900 29986 39956 30716
rect 40348 30548 40404 30558
rect 39900 29934 39902 29986
rect 39954 29934 39956 29986
rect 39900 29922 39956 29934
rect 40124 30324 40180 30334
rect 39452 29650 39508 29662
rect 39452 29598 39454 29650
rect 39506 29598 39508 29650
rect 39116 28868 39172 28878
rect 39452 28868 39508 29598
rect 40124 29090 40180 30268
rect 40348 29986 40404 30492
rect 40348 29934 40350 29986
rect 40402 29934 40404 29986
rect 40348 29922 40404 29934
rect 40124 29038 40126 29090
rect 40178 29038 40180 29090
rect 40124 29026 40180 29038
rect 39900 28868 39956 28878
rect 39116 28866 39900 28868
rect 39116 28814 39118 28866
rect 39170 28814 39900 28866
rect 39116 28812 39900 28814
rect 38556 28578 38612 28588
rect 38780 28642 38836 28654
rect 38780 28590 38782 28642
rect 38834 28590 38836 28642
rect 38780 28532 38836 28590
rect 39116 28644 39172 28812
rect 39900 28774 39956 28812
rect 40460 28756 40516 34188
rect 40572 34178 40628 34188
rect 40908 33348 40964 36764
rect 41132 36594 41188 36606
rect 41132 36542 41134 36594
rect 41186 36542 41188 36594
rect 41020 34804 41076 34814
rect 41020 34020 41076 34748
rect 41020 33926 41076 33964
rect 40684 33292 40964 33348
rect 40684 31332 40740 33292
rect 40796 33124 40852 33134
rect 41132 33124 41188 36542
rect 41244 36036 41300 36046
rect 41244 35810 41300 35980
rect 41244 35758 41246 35810
rect 41298 35758 41300 35810
rect 41244 35746 41300 35758
rect 40796 33122 41188 33124
rect 40796 33070 40798 33122
rect 40850 33070 41188 33122
rect 40796 33068 41188 33070
rect 41244 33684 41300 33694
rect 40796 33058 40852 33068
rect 41244 32114 41300 33628
rect 41356 33460 41412 39004
rect 41692 38836 41748 40012
rect 42364 40002 42420 40012
rect 42476 39956 42532 39966
rect 42588 39956 42644 41022
rect 43036 41746 43092 41758
rect 43036 41694 43038 41746
rect 43090 41694 43092 41746
rect 43036 40964 43092 41694
rect 43036 40898 43092 40908
rect 42924 40850 42980 40862
rect 42924 40798 42926 40850
rect 42978 40798 42980 40850
rect 42476 39954 42644 39956
rect 42476 39902 42478 39954
rect 42530 39902 42644 39954
rect 42476 39900 42644 39902
rect 42700 40740 42756 40750
rect 42924 40740 42980 40798
rect 43036 40740 43092 40750
rect 42924 40738 43092 40740
rect 42924 40686 43038 40738
rect 43090 40686 43092 40738
rect 42924 40684 43092 40686
rect 42476 39890 42532 39900
rect 41916 39844 41972 39854
rect 41916 39750 41972 39788
rect 41468 38780 41748 38836
rect 42252 38834 42308 38846
rect 42252 38782 42254 38834
rect 42306 38782 42308 38834
rect 41468 34244 41524 38780
rect 42028 38724 42084 38734
rect 41916 38612 41972 38622
rect 41580 38610 41972 38612
rect 41580 38558 41918 38610
rect 41970 38558 41972 38610
rect 41580 38556 41972 38558
rect 41580 37938 41636 38556
rect 41916 38546 41972 38556
rect 42028 38388 42084 38668
rect 41916 38332 42084 38388
rect 41916 38050 41972 38332
rect 41916 37998 41918 38050
rect 41970 37998 41972 38050
rect 41916 37986 41972 37998
rect 41580 37886 41582 37938
rect 41634 37886 41636 37938
rect 41580 37874 41636 37886
rect 42252 37604 42308 38782
rect 42700 38722 42756 40684
rect 43036 40674 43092 40684
rect 43036 39956 43092 39966
rect 43148 39956 43204 43708
rect 43932 42644 43988 42654
rect 43932 42642 44100 42644
rect 43932 42590 43934 42642
rect 43986 42590 44100 42642
rect 43932 42588 44100 42590
rect 43932 42578 43988 42588
rect 43932 41972 43988 41982
rect 43484 41746 43540 41758
rect 43484 41694 43486 41746
rect 43538 41694 43540 41746
rect 43484 41636 43540 41694
rect 43484 40852 43540 41580
rect 43932 40964 43988 41916
rect 44044 41860 44100 42588
rect 44940 42642 44996 42654
rect 44940 42590 44942 42642
rect 44994 42590 44996 42642
rect 44940 42530 44996 42590
rect 44940 42478 44942 42530
rect 44994 42478 44996 42530
rect 44380 41972 44436 41982
rect 44716 41972 44772 41982
rect 44436 41916 44548 41972
rect 44380 41906 44436 41916
rect 44268 41860 44324 41870
rect 44044 41804 44268 41860
rect 44268 41766 44324 41804
rect 44492 41858 44548 41916
rect 44492 41806 44494 41858
rect 44546 41806 44548 41858
rect 44492 41748 44548 41806
rect 44716 41858 44772 41916
rect 44716 41806 44718 41858
rect 44770 41806 44772 41858
rect 44716 41794 44772 41806
rect 44940 41860 44996 42478
rect 44940 41794 44996 41804
rect 45388 42642 45444 44046
rect 45500 44660 45556 44670
rect 45500 43652 45556 44604
rect 45724 43764 45780 43802
rect 46060 43708 46116 45838
rect 48188 45890 48244 45902
rect 48188 45838 48190 45890
rect 48242 45838 48244 45890
rect 45724 43698 45780 43708
rect 45500 43586 45556 43596
rect 45836 43652 46116 43708
rect 46508 44770 46564 44782
rect 46508 44718 46510 44770
rect 46562 44718 46564 44770
rect 46508 43764 46564 44718
rect 47292 44770 47348 44782
rect 47292 44718 47294 44770
rect 47346 44718 47348 44770
rect 46508 43698 46564 43708
rect 46956 43762 47012 43774
rect 46956 43710 46958 43762
rect 47010 43710 47012 43762
rect 45388 42590 45390 42642
rect 45442 42590 45444 42642
rect 45388 42196 45444 42590
rect 45388 41972 45444 42140
rect 44492 41682 44548 41692
rect 43932 40898 43988 40908
rect 45052 41522 45108 41534
rect 45052 41470 45054 41522
rect 45106 41470 45108 41522
rect 43036 39954 43204 39956
rect 43036 39902 43038 39954
rect 43090 39902 43204 39954
rect 43036 39900 43204 39902
rect 43260 40796 43484 40852
rect 43036 39890 43092 39900
rect 43260 39060 43316 40796
rect 43484 40786 43540 40796
rect 44044 40852 44100 40862
rect 44044 40758 44100 40796
rect 43036 39004 43316 39060
rect 43484 40626 43540 40638
rect 43484 40574 43486 40626
rect 43538 40574 43540 40626
rect 43484 40514 43540 40574
rect 43484 40462 43486 40514
rect 43538 40462 43540 40514
rect 43036 38948 43092 39004
rect 42700 38670 42702 38722
rect 42754 38670 42756 38722
rect 42700 38668 42756 38670
rect 42588 38612 42756 38668
rect 42924 38946 43092 38948
rect 42924 38894 43038 38946
rect 43090 38894 43092 38946
rect 42924 38892 43092 38894
rect 42476 37828 42532 37838
rect 42476 37734 42532 37772
rect 42252 37538 42308 37548
rect 42588 37716 42644 38612
rect 41916 36594 41972 36606
rect 41916 36542 41918 36594
rect 41970 36542 41972 36594
rect 41916 36036 41972 36542
rect 41916 35970 41972 35980
rect 42252 36036 42308 36046
rect 41580 34804 41636 34814
rect 41580 34710 41636 34748
rect 41468 34178 41524 34188
rect 41692 34692 41748 34702
rect 41692 34132 41748 34636
rect 42252 34692 42308 35980
rect 42588 34916 42644 37660
rect 42924 36818 42980 38892
rect 43036 38882 43092 38892
rect 43036 37828 43092 37838
rect 43484 37828 43540 40462
rect 44940 40626 44996 40638
rect 44940 40574 44942 40626
rect 44994 40574 44996 40626
rect 43708 40068 43764 40078
rect 43708 39974 43764 40012
rect 44940 39956 44996 40574
rect 44940 39890 44996 39900
rect 45052 39954 45108 41470
rect 45388 40852 45444 41916
rect 45836 42642 45892 43652
rect 46060 43540 46116 43652
rect 46060 43474 46116 43484
rect 46732 43652 46788 43662
rect 46732 42978 46788 43596
rect 46732 42926 46734 42978
rect 46786 42926 46788 42978
rect 46732 42914 46788 42926
rect 45836 42590 45838 42642
rect 45890 42590 45892 42642
rect 45612 41860 45668 41870
rect 45836 41860 45892 42590
rect 46284 42642 46340 42654
rect 46284 42590 46286 42642
rect 46338 42590 46340 42642
rect 46284 42530 46340 42590
rect 46284 42478 46286 42530
rect 46338 42478 46340 42530
rect 46284 42466 46340 42478
rect 46732 42196 46788 42206
rect 46956 42196 47012 43710
rect 47292 43652 47348 44718
rect 48188 44098 48244 45838
rect 50556 44380 50820 44390
rect 50612 44324 50660 44380
rect 50716 44324 50764 44380
rect 50556 44314 50820 44324
rect 48188 44046 48190 44098
rect 48242 44046 48244 44098
rect 47292 42756 47348 43596
rect 47404 43762 47460 43774
rect 47404 43710 47406 43762
rect 47458 43710 47460 43762
rect 47404 43540 47460 43710
rect 47404 43474 47460 43484
rect 47964 43540 48020 43550
rect 47964 42868 48020 43484
rect 47964 42774 48020 42812
rect 48076 42978 48132 42990
rect 48076 42926 48078 42978
rect 48130 42926 48132 42978
rect 47516 42756 47572 42766
rect 47292 42700 47516 42756
rect 47516 42662 47572 42700
rect 47740 42754 47796 42766
rect 47740 42702 47742 42754
rect 47794 42702 47796 42754
rect 47180 42644 47236 42654
rect 47180 42642 47348 42644
rect 47180 42590 47182 42642
rect 47234 42590 47348 42642
rect 47180 42588 47348 42590
rect 47180 42578 47236 42588
rect 46788 42140 47012 42196
rect 47292 42530 47348 42588
rect 47292 42478 47294 42530
rect 47346 42478 47348 42530
rect 46732 41970 46788 42140
rect 46732 41918 46734 41970
rect 46786 41918 46788 41970
rect 46732 41906 46788 41918
rect 47180 42082 47236 42094
rect 47180 42030 47182 42082
rect 47234 42030 47236 42082
rect 45612 41858 46228 41860
rect 45612 41806 45614 41858
rect 45666 41806 46228 41858
rect 45612 41804 46228 41806
rect 45612 41748 45668 41804
rect 45612 41682 45668 41692
rect 45388 40758 45444 40796
rect 46172 40850 46228 41804
rect 46172 40798 46174 40850
rect 46226 40798 46228 40850
rect 46172 40786 46228 40798
rect 46732 40852 46788 40862
rect 46732 40758 46788 40796
rect 46732 40180 46788 40190
rect 45052 39902 45054 39954
rect 45106 39902 45108 39954
rect 45052 39890 45108 39902
rect 45724 39956 45780 39966
rect 45724 39862 45780 39900
rect 46508 39954 46564 39966
rect 46508 39902 46510 39954
rect 46562 39902 46564 39954
rect 44492 39844 44548 39854
rect 44492 39750 44548 39788
rect 45388 39844 45444 39854
rect 46060 39844 46116 39854
rect 45388 39750 45444 39788
rect 45948 39842 46116 39844
rect 45948 39790 46062 39842
rect 46114 39790 46116 39842
rect 45948 39788 46116 39790
rect 44940 38836 44996 38846
rect 44940 38610 44996 38780
rect 44940 38558 44942 38610
rect 44994 38558 44996 38610
rect 43708 37940 43764 37950
rect 44940 37940 44996 38558
rect 43708 37938 43876 37940
rect 43708 37886 43710 37938
rect 43762 37886 43876 37938
rect 43708 37884 43876 37886
rect 43708 37874 43764 37884
rect 43036 37826 43204 37828
rect 43036 37774 43038 37826
rect 43090 37774 43204 37826
rect 43036 37772 43204 37774
rect 43036 37762 43092 37772
rect 42924 36766 42926 36818
rect 42978 36766 42980 36818
rect 42924 35924 42980 36766
rect 43036 37604 43092 37614
rect 43036 36818 43092 37548
rect 43036 36766 43038 36818
rect 43090 36766 43092 36818
rect 43036 36754 43092 36766
rect 43148 36596 43204 37772
rect 43484 37762 43540 37772
rect 43820 37154 43876 37884
rect 44828 37884 44996 37940
rect 45948 37940 46004 39788
rect 46060 39778 46116 39788
rect 46508 38836 46564 39902
rect 46508 38770 46564 38780
rect 46732 38834 46788 40124
rect 47180 39954 47236 42030
rect 47292 41972 47348 42478
rect 47740 42196 47796 42702
rect 47740 42130 47796 42140
rect 47516 41972 47572 41982
rect 47292 41970 47572 41972
rect 47292 41918 47518 41970
rect 47570 41918 47572 41970
rect 47292 41916 47572 41918
rect 47516 41860 47572 41916
rect 47516 40852 47572 41804
rect 47516 40758 47572 40796
rect 47852 40068 47908 40078
rect 48076 40068 48132 42926
rect 48188 42866 48244 44046
rect 54124 43874 54180 43886
rect 54124 43822 54126 43874
rect 54178 43822 54180 43874
rect 51772 43762 51828 43774
rect 51772 43710 51774 43762
rect 51826 43710 51828 43762
rect 48188 42814 48190 42866
rect 48242 42814 48244 42866
rect 48188 42644 48244 42814
rect 49420 42868 49476 42878
rect 48860 42756 48916 42766
rect 48636 42644 48692 42654
rect 48188 42642 48692 42644
rect 48188 42590 48638 42642
rect 48690 42590 48692 42642
rect 48188 42588 48692 42590
rect 48636 41860 48692 42588
rect 48860 42084 48916 42700
rect 49084 42642 49140 42654
rect 49084 42590 49086 42642
rect 49138 42590 49140 42642
rect 49084 42196 49140 42590
rect 49084 42130 49140 42140
rect 49420 42644 49476 42812
rect 49532 42644 49588 42654
rect 49420 42642 49588 42644
rect 49420 42590 49534 42642
rect 49586 42590 49588 42642
rect 49420 42588 49588 42590
rect 48860 41970 48916 42028
rect 48860 41918 48862 41970
rect 48914 41918 48916 41970
rect 48860 41906 48916 41918
rect 49308 42084 49364 42094
rect 48636 41794 48692 41804
rect 49196 41860 49252 41870
rect 49196 41766 49252 41804
rect 47852 40066 48132 40068
rect 47852 40014 47854 40066
rect 47906 40014 48132 40066
rect 47852 40012 48132 40014
rect 47852 40002 47908 40012
rect 47180 39902 47182 39954
rect 47234 39902 47236 39954
rect 47180 39890 47236 39902
rect 48748 39956 48804 39966
rect 46732 38782 46734 38834
rect 46786 38782 46788 38834
rect 46732 38770 46788 38782
rect 46844 39844 46900 39854
rect 46284 38500 46340 38510
rect 43820 37102 43822 37154
rect 43874 37102 43876 37154
rect 43820 37090 43876 37102
rect 44492 37828 44548 37838
rect 43932 36820 43988 36830
rect 43820 36818 43988 36820
rect 43820 36766 43934 36818
rect 43986 36766 43988 36818
rect 43820 36764 43988 36766
rect 43148 36530 43204 36540
rect 43484 36708 43540 36718
rect 43148 35924 43204 35934
rect 42924 35922 43204 35924
rect 42924 35870 43150 35922
rect 43202 35870 43204 35922
rect 42924 35868 43204 35870
rect 43148 35700 43204 35868
rect 43484 35810 43540 36652
rect 43820 36036 43876 36764
rect 43932 36754 43988 36764
rect 44044 36818 44100 36830
rect 44044 36766 44046 36818
rect 44098 36766 44100 36818
rect 44044 36708 44100 36766
rect 44100 36652 44324 36708
rect 44044 36642 44100 36652
rect 43820 35970 43876 35980
rect 43932 36596 43988 36606
rect 43484 35758 43486 35810
rect 43538 35758 43540 35810
rect 43484 35746 43540 35758
rect 43148 35634 43204 35644
rect 43932 35698 43988 36540
rect 43932 35646 43934 35698
rect 43986 35646 43988 35698
rect 43932 35634 43988 35646
rect 42588 34850 42644 34860
rect 43596 34916 43652 34926
rect 42252 34598 42308 34636
rect 42364 34804 42420 34814
rect 41580 34076 41748 34132
rect 41804 34132 41860 34142
rect 41468 34020 41524 34030
rect 41580 34020 41636 34076
rect 41468 34018 41636 34020
rect 41468 33966 41470 34018
rect 41522 33966 41636 34018
rect 41468 33964 41636 33966
rect 41468 33954 41524 33964
rect 41804 33684 41860 34076
rect 42364 34018 42420 34748
rect 42364 33966 42366 34018
rect 42418 33966 42420 34018
rect 42364 33954 42420 33966
rect 42812 34692 42868 34702
rect 42812 33906 42868 34636
rect 42812 33854 42814 33906
rect 42866 33854 42868 33906
rect 42812 33842 42868 33854
rect 43260 34580 43316 34590
rect 43148 33794 43204 33806
rect 43148 33742 43150 33794
rect 43202 33742 43204 33794
rect 41916 33684 41972 33694
rect 41804 33682 41972 33684
rect 41804 33630 41918 33682
rect 41970 33630 41972 33682
rect 41804 33628 41972 33630
rect 41356 33404 41636 33460
rect 41244 32062 41246 32114
rect 41298 32062 41300 32114
rect 41244 32050 41300 32062
rect 40908 31778 40964 31790
rect 40908 31726 40910 31778
rect 40962 31726 40964 31778
rect 40908 31668 40964 31726
rect 40908 31602 40964 31612
rect 40684 31276 41300 31332
rect 40572 31108 40628 31118
rect 40572 30882 40628 31052
rect 40572 30830 40574 30882
rect 40626 30830 40628 30882
rect 40572 30818 40628 30830
rect 41132 31108 41188 31118
rect 41132 30770 41188 31052
rect 41132 30718 41134 30770
rect 41186 30718 41188 30770
rect 41132 30706 41188 30718
rect 41244 29874 41300 31276
rect 41356 30772 41412 30782
rect 41356 30678 41412 30716
rect 41244 29822 41246 29874
rect 41298 29822 41300 29874
rect 41244 29810 41300 29822
rect 41468 29764 41524 29774
rect 41356 29762 41524 29764
rect 41356 29710 41470 29762
rect 41522 29710 41524 29762
rect 41356 29708 41524 29710
rect 40796 29428 40852 29438
rect 40796 29334 40852 29372
rect 41244 28868 41300 28878
rect 41356 28868 41412 29708
rect 41468 29698 41524 29708
rect 41300 28812 41412 28868
rect 41244 28774 41300 28812
rect 40572 28756 40628 28766
rect 40460 28754 40628 28756
rect 40460 28702 40574 28754
rect 40626 28702 40628 28754
rect 40460 28700 40628 28702
rect 40572 28690 40628 28700
rect 41020 28644 41076 28654
rect 39116 28578 39172 28588
rect 40908 28642 41076 28644
rect 40908 28590 41022 28642
rect 41074 28590 41076 28642
rect 40908 28588 41076 28590
rect 38780 28466 38836 28476
rect 38444 28030 38446 28082
rect 38498 28030 38500 28082
rect 38444 27972 38500 28030
rect 39452 28082 39508 28094
rect 39452 28030 39454 28082
rect 39506 28030 39508 28082
rect 38556 27972 38612 27982
rect 39452 27972 39508 28030
rect 38444 27970 38612 27972
rect 38444 27918 38558 27970
rect 38610 27918 38612 27970
rect 38444 27916 38612 27918
rect 38556 27906 38612 27916
rect 39340 27970 39508 27972
rect 39340 27918 39454 27970
rect 39506 27918 39508 27970
rect 39340 27916 39508 27918
rect 39004 27634 39060 27646
rect 39004 27582 39006 27634
rect 39058 27582 39060 27634
rect 38444 26626 38500 26638
rect 38444 26574 38446 26626
rect 38498 26574 38500 26626
rect 38444 25620 38500 26574
rect 38780 26628 38836 26638
rect 38780 26534 38836 26572
rect 38668 26292 38724 26302
rect 39004 26292 39060 27582
rect 39340 27076 39396 27916
rect 39452 27906 39508 27916
rect 38724 26236 39060 26292
rect 39116 26626 39172 26638
rect 39116 26574 39118 26626
rect 39170 26574 39172 26626
rect 38668 25732 38724 26236
rect 38556 25620 38612 25630
rect 38444 25618 38612 25620
rect 38444 25566 38558 25618
rect 38610 25566 38612 25618
rect 38444 25564 38612 25566
rect 38556 25554 38612 25564
rect 38668 24722 38724 25676
rect 39116 25730 39172 26574
rect 39116 25678 39118 25730
rect 39170 25678 39172 25730
rect 39116 25666 39172 25678
rect 39340 25732 39396 27020
rect 40348 27634 40404 27646
rect 40348 27582 40350 27634
rect 40402 27582 40404 27634
rect 40348 26964 40404 27582
rect 39452 26852 39508 26862
rect 39452 26738 39508 26796
rect 39452 26686 39454 26738
rect 39506 26686 39508 26738
rect 39452 26674 39508 26686
rect 39900 26626 39956 26638
rect 39900 26574 39902 26626
rect 39954 26574 39956 26626
rect 39676 25732 39732 25742
rect 39340 25730 39620 25732
rect 39340 25678 39342 25730
rect 39394 25678 39620 25730
rect 39340 25676 39620 25678
rect 39340 25666 39396 25676
rect 39564 25508 39620 25676
rect 39676 25638 39732 25676
rect 39564 25452 39844 25508
rect 38668 24670 38670 24722
rect 38722 24670 38724 24722
rect 38668 22596 38724 24670
rect 38892 24724 38948 24734
rect 38892 24612 38948 24668
rect 39788 24724 39844 25452
rect 39788 24630 39844 24668
rect 38892 24610 39060 24612
rect 38892 24558 38894 24610
rect 38946 24558 39060 24610
rect 38892 24556 39060 24558
rect 38892 24546 38948 24556
rect 38780 23828 38836 23838
rect 38780 23734 38836 23772
rect 38892 22820 38948 22830
rect 39004 22820 39060 24556
rect 39900 23828 39956 26574
rect 40348 25732 40404 26908
rect 40348 24724 40404 25676
rect 40236 24722 40404 24724
rect 40236 24670 40350 24722
rect 40402 24670 40404 24722
rect 40236 24668 40404 24670
rect 39900 23762 39956 23772
rect 40012 23826 40068 23838
rect 40012 23774 40014 23826
rect 40066 23774 40068 23826
rect 39340 23714 39396 23726
rect 39340 23662 39342 23714
rect 39394 23662 39396 23714
rect 39340 23044 39396 23662
rect 40012 23492 40068 23774
rect 40012 23426 40068 23436
rect 39340 22978 39396 22988
rect 40124 23044 40180 23054
rect 40124 22950 40180 22988
rect 38892 22818 39060 22820
rect 38892 22766 38894 22818
rect 38946 22766 39060 22818
rect 38892 22764 39060 22766
rect 38892 22754 38948 22764
rect 39116 22596 39172 22606
rect 38668 22594 39620 22596
rect 38668 22542 39118 22594
rect 39170 22542 39620 22594
rect 38668 22540 39620 22542
rect 39116 22530 39172 22540
rect 39564 21922 39620 22540
rect 40236 22594 40292 24668
rect 40348 24658 40404 24668
rect 40572 26626 40628 26638
rect 40572 26574 40574 26626
rect 40626 26574 40628 26626
rect 40572 24388 40628 26574
rect 40572 24322 40628 24332
rect 40572 23940 40628 23950
rect 40460 23884 40572 23940
rect 40460 22706 40516 23884
rect 40572 23874 40628 23884
rect 40796 23492 40852 23502
rect 40908 23492 40964 28588
rect 41020 28578 41076 28588
rect 41020 27634 41076 27646
rect 41020 27582 41022 27634
rect 41074 27582 41076 27634
rect 41020 27076 41076 27582
rect 41020 25730 41076 27020
rect 41244 26516 41300 26526
rect 41132 26514 41300 26516
rect 41132 26462 41246 26514
rect 41298 26462 41300 26514
rect 41132 26460 41300 26462
rect 41132 26066 41188 26460
rect 41244 26450 41300 26460
rect 41132 26014 41134 26066
rect 41186 26014 41188 26066
rect 41132 26002 41188 26014
rect 41020 25678 41022 25730
rect 41074 25678 41076 25730
rect 41020 23940 41076 25678
rect 41244 25842 41300 25854
rect 41244 25790 41246 25842
rect 41298 25790 41300 25842
rect 41244 25732 41300 25790
rect 41300 25676 41412 25732
rect 41244 25666 41300 25676
rect 41356 24164 41412 25676
rect 41468 24388 41524 24398
rect 41468 24294 41524 24332
rect 41356 24108 41524 24164
rect 41020 23874 41076 23884
rect 41356 23940 41412 23950
rect 41132 23716 41188 23726
rect 41132 23714 41300 23716
rect 41132 23662 41134 23714
rect 41186 23662 41300 23714
rect 41132 23660 41300 23662
rect 41132 23650 41188 23660
rect 41244 23604 41300 23660
rect 40908 23436 41188 23492
rect 40796 23398 40852 23436
rect 40908 22818 40964 22830
rect 40908 22766 40910 22818
rect 40962 22766 40964 22818
rect 40460 22654 40462 22706
rect 40514 22654 40516 22706
rect 40460 22642 40516 22654
rect 40684 22706 40740 22718
rect 40684 22654 40686 22706
rect 40738 22654 40740 22706
rect 40236 22542 40238 22594
rect 40290 22542 40292 22594
rect 40236 22530 40292 22542
rect 40572 22596 40628 22606
rect 40684 22596 40740 22654
rect 40628 22540 40740 22596
rect 40908 22706 40964 22766
rect 40908 22654 40910 22706
rect 40962 22654 40964 22706
rect 40572 22530 40628 22540
rect 39564 21870 39566 21922
rect 39618 21870 39620 21922
rect 39564 21858 39620 21870
rect 38332 20738 38388 20748
rect 38668 21586 38724 21598
rect 38668 21534 38670 21586
rect 38722 21534 38724 21586
rect 38668 21474 38724 21534
rect 38668 21422 38670 21474
rect 38722 21422 38724 21474
rect 37548 20638 37550 20690
rect 37602 20638 37604 20690
rect 37548 20626 37604 20638
rect 37100 20402 37156 20412
rect 38332 20468 38388 20478
rect 36316 19682 36372 19694
rect 36316 19630 36318 19682
rect 36370 19630 36372 19682
rect 36316 18676 36372 19630
rect 36316 18610 36372 18620
rect 36428 18898 36484 18910
rect 36428 18846 36430 18898
rect 36482 18846 36484 18898
rect 36428 18786 36484 18846
rect 36428 18734 36430 18786
rect 36482 18734 36484 18786
rect 36204 18498 36260 18508
rect 34748 18386 34804 18396
rect 35084 18450 35140 18462
rect 35084 18398 35086 18450
rect 35138 18398 35140 18450
rect 35084 18228 35140 18398
rect 34076 18172 35140 18228
rect 34972 16772 35028 16782
rect 34972 16678 35028 16716
rect 33852 16546 33908 16558
rect 33852 16494 33854 16546
rect 33906 16494 33908 16546
rect 33516 16436 33572 16446
rect 33852 16436 33908 16494
rect 33516 16434 33908 16436
rect 33516 16382 33518 16434
rect 33570 16382 33908 16434
rect 33516 16380 33908 16382
rect 32284 14418 32340 15148
rect 32844 15092 33012 15148
rect 33068 15764 33124 15774
rect 33516 15764 33572 16380
rect 33068 15762 33572 15764
rect 33068 15710 33070 15762
rect 33122 15710 33572 15762
rect 33068 15708 33572 15710
rect 32732 14868 32788 14878
rect 32732 14754 32788 14812
rect 32732 14702 32734 14754
rect 32786 14702 32788 14754
rect 32732 14690 32788 14702
rect 32284 14366 32286 14418
rect 32338 14366 32340 14418
rect 32060 13860 32116 13870
rect 32060 13766 32116 13804
rect 32284 13636 32340 14366
rect 32508 13636 32564 13646
rect 32284 13580 32508 13636
rect 32508 13542 32564 13580
rect 30828 13458 30884 13468
rect 32844 13412 32900 15092
rect 33068 14868 33124 15708
rect 35084 15652 35140 18172
rect 35308 18452 35364 18462
rect 35308 17890 35364 18396
rect 36428 18340 36484 18734
rect 37660 18676 37716 18686
rect 36428 18274 36484 18284
rect 37548 18564 37604 18574
rect 35308 17838 35310 17890
rect 35362 17838 35364 17890
rect 35308 17826 35364 17838
rect 35196 17164 35460 17174
rect 35252 17108 35300 17164
rect 35356 17108 35404 17164
rect 35196 17098 35460 17108
rect 36764 16772 36820 16782
rect 37436 16772 37492 16782
rect 36204 15764 36260 15774
rect 36204 15670 36260 15708
rect 36764 15762 36820 16716
rect 36764 15710 36766 15762
rect 36818 15710 36820 15762
rect 36764 15698 36820 15710
rect 37324 16716 37436 16772
rect 37324 16658 37380 16716
rect 37436 16706 37492 16716
rect 37324 16606 37326 16658
rect 37378 16606 37380 16658
rect 35084 15148 35140 15596
rect 37100 15650 37156 15662
rect 37100 15598 37102 15650
rect 37154 15598 37156 15650
rect 33068 14802 33124 14812
rect 34636 15092 35140 15148
rect 35196 15148 35460 15158
rect 35252 15092 35300 15148
rect 35356 15092 35404 15148
rect 37100 15148 37156 15598
rect 37100 15092 37268 15148
rect 33180 14644 33236 14654
rect 33180 14550 33236 14588
rect 34076 14532 34132 14542
rect 34076 14438 34132 14476
rect 33516 14308 33572 14318
rect 33404 14252 33516 14308
rect 31948 12964 32004 12974
rect 31948 12870 32004 12908
rect 32844 12740 32900 13356
rect 32732 12684 32844 12740
rect 32732 12626 32788 12684
rect 32844 12674 32900 12684
rect 33180 13748 33236 13758
rect 33180 13522 33236 13692
rect 33180 13470 33182 13522
rect 33234 13470 33236 13522
rect 32732 12574 32734 12626
rect 32786 12574 32788 12626
rect 32732 12562 32788 12574
rect 32396 12516 32452 12526
rect 32172 12514 32452 12516
rect 32172 12462 32398 12514
rect 32450 12462 32452 12514
rect 32172 12460 32452 12462
rect 30940 11618 30996 11630
rect 30940 11566 30942 11618
rect 30994 11566 30996 11618
rect 29148 11508 29204 11518
rect 28812 11506 29204 11508
rect 28812 11454 29150 11506
rect 29202 11454 29204 11506
rect 28812 11452 29204 11454
rect 28700 11230 28702 11282
rect 28754 11230 28756 11282
rect 28700 11218 28756 11230
rect 28252 10434 28308 10444
rect 27468 9714 27524 10108
rect 27468 9662 27470 9714
rect 27522 9662 27524 9714
rect 27468 9650 27524 9662
rect 28588 10386 28644 10398
rect 28588 10334 28590 10386
rect 28642 10334 28644 10386
rect 28588 9716 28644 10334
rect 28588 9650 28644 9660
rect 28700 9714 28756 9726
rect 28700 9662 28702 9714
rect 28754 9662 28756 9714
rect 28028 9604 28084 9614
rect 28028 9602 28308 9604
rect 28028 9550 28030 9602
rect 28082 9550 28308 9602
rect 28028 9548 28308 9550
rect 28028 9538 28084 9548
rect 28252 8818 28308 9548
rect 28252 8766 28254 8818
rect 28306 8766 28308 8818
rect 28252 8754 28308 8766
rect 27356 7746 27412 7756
rect 28700 7700 28756 9662
rect 29148 8596 29204 11452
rect 30604 11508 30660 11518
rect 30940 11508 30996 11566
rect 30604 11506 30996 11508
rect 30604 11454 30606 11506
rect 30658 11454 30996 11506
rect 30604 11452 30996 11454
rect 29260 11284 29316 11294
rect 29260 11282 29428 11284
rect 29260 11230 29262 11282
rect 29314 11230 29428 11282
rect 29260 11228 29428 11230
rect 29260 11218 29316 11228
rect 29372 10498 29428 11228
rect 30044 10724 30100 10734
rect 29372 10446 29374 10498
rect 29426 10446 29428 10498
rect 29148 8530 29204 8540
rect 29260 9716 29316 9726
rect 29260 8594 29316 9660
rect 29372 8708 29428 10446
rect 29708 10500 29764 10510
rect 29708 10406 29764 10444
rect 30044 10498 30100 10668
rect 30044 10446 30046 10498
rect 30098 10446 30100 10498
rect 30044 10434 30100 10446
rect 30604 10610 30660 11452
rect 30604 10558 30606 10610
rect 30658 10558 30660 10610
rect 29596 9716 29652 9726
rect 29596 9622 29652 9660
rect 30604 9716 30660 10558
rect 29372 8642 29428 8652
rect 30268 8708 30324 8718
rect 30324 8652 30436 8708
rect 30268 8614 30324 8652
rect 29260 8542 29262 8594
rect 29314 8542 29316 8594
rect 29260 8428 29316 8542
rect 29820 8596 29876 8606
rect 29820 8502 29876 8540
rect 29260 8372 29428 8428
rect 29260 7700 29316 7710
rect 28700 7698 29316 7700
rect 28700 7646 29262 7698
rect 29314 7646 29316 7698
rect 28700 7644 29316 7646
rect 29260 7634 29316 7644
rect 27468 6692 27524 6702
rect 27020 6580 27076 6590
rect 27020 5906 27076 6524
rect 27020 5854 27022 5906
rect 27074 5854 27076 5906
rect 27020 5794 27076 5854
rect 27020 5742 27022 5794
rect 27074 5742 27076 5794
rect 27020 5730 27076 5742
rect 27468 5794 27524 6636
rect 28924 6692 28980 6702
rect 28812 6580 28868 6590
rect 28476 6466 28532 6478
rect 28476 6414 28478 6466
rect 28530 6414 28532 6466
rect 27468 5742 27470 5794
rect 27522 5742 27524 5794
rect 27468 5730 27524 5742
rect 27916 5906 27972 5918
rect 27916 5854 27918 5906
rect 27970 5854 27972 5906
rect 27916 5796 27972 5854
rect 27916 5702 27972 5740
rect 28364 5796 28420 5806
rect 28476 5796 28532 6414
rect 28364 5794 28532 5796
rect 28364 5742 28366 5794
rect 28418 5742 28532 5794
rect 28364 5740 28532 5742
rect 28364 5730 28420 5740
rect 28476 5572 28532 5740
rect 28812 5572 28868 6524
rect 28476 5570 28868 5572
rect 28476 5518 28814 5570
rect 28866 5518 28868 5570
rect 28476 5516 28868 5518
rect 28476 5460 28532 5516
rect 28812 5506 28868 5516
rect 26684 4610 26740 4620
rect 27692 4676 27748 4686
rect 27692 4582 27748 4620
rect 28476 4674 28532 5404
rect 28476 4622 28478 4674
rect 28530 4622 28532 4674
rect 28476 4610 28532 4622
rect 28924 4674 28980 6636
rect 29260 6580 29316 6590
rect 29372 6580 29428 8372
rect 30268 7924 30324 7934
rect 30268 7810 30324 7868
rect 30268 7758 30270 7810
rect 30322 7758 30324 7810
rect 30268 7746 30324 7758
rect 30380 6692 30436 8652
rect 30604 7812 30660 9660
rect 30716 10724 30772 10734
rect 30716 8708 30772 10668
rect 30716 8614 30772 8652
rect 31276 10500 31332 10510
rect 31276 8820 31332 10444
rect 32172 9828 32228 12460
rect 32396 12450 32452 12460
rect 32844 12514 32900 12526
rect 32844 12462 32846 12514
rect 32898 12462 32900 12514
rect 32844 11844 32900 12462
rect 32844 11778 32900 11788
rect 32284 11620 32340 11630
rect 33068 11620 33124 11630
rect 32284 11618 33124 11620
rect 32284 11566 32286 11618
rect 32338 11566 33070 11618
rect 33122 11566 33124 11618
rect 32284 11564 33124 11566
rect 32284 11554 32340 11564
rect 33068 11554 33124 11564
rect 32172 9762 32228 9772
rect 32396 10500 32452 10510
rect 31276 8764 31668 8820
rect 31164 8484 31220 8494
rect 30716 7812 30772 7822
rect 31164 7812 31220 8428
rect 31276 7922 31332 8764
rect 31276 7870 31278 7922
rect 31330 7870 31332 7922
rect 31276 7858 31332 7870
rect 31388 8596 31444 8606
rect 30604 7810 31220 7812
rect 30604 7758 30718 7810
rect 30770 7758 31166 7810
rect 31218 7758 31220 7810
rect 30604 7756 31220 7758
rect 30716 7746 30772 7756
rect 31164 7746 31220 7756
rect 30380 6626 30436 6636
rect 29316 6524 29428 6580
rect 29260 6486 29316 6524
rect 29932 6468 29988 6478
rect 29820 6466 29988 6468
rect 29820 6414 29934 6466
rect 29986 6414 29988 6466
rect 29820 6412 29988 6414
rect 31388 6468 31444 8540
rect 31612 8594 31668 8764
rect 31612 8542 31614 8594
rect 31666 8542 31668 8594
rect 31612 8530 31668 8542
rect 32060 8708 32116 8718
rect 32060 8594 32116 8652
rect 32060 8542 32062 8594
rect 32114 8542 32116 8594
rect 32060 8530 32116 8542
rect 31948 7476 32004 7486
rect 31836 7474 32004 7476
rect 31836 7422 31950 7474
rect 32002 7422 32004 7474
rect 31836 7420 32004 7422
rect 31836 6580 31892 7420
rect 31948 7410 32004 7420
rect 32396 7474 32452 10444
rect 33068 10500 33124 10510
rect 33180 10500 33236 13470
rect 33124 10444 33236 10500
rect 33404 11730 33460 14252
rect 33516 14214 33572 14252
rect 33740 13748 33796 13758
rect 33740 13634 33796 13692
rect 33740 13582 33742 13634
rect 33794 13582 33796 13634
rect 33740 13570 33796 13582
rect 33964 13636 34020 13646
rect 33964 13542 34020 13580
rect 33628 13524 33684 13534
rect 33628 12962 33684 13468
rect 33628 12910 33630 12962
rect 33682 12910 33684 12962
rect 33628 12738 33684 12910
rect 33628 12686 33630 12738
rect 33682 12686 33684 12738
rect 33628 12674 33684 12686
rect 34076 13524 34132 13534
rect 34076 12738 34132 13468
rect 34300 13522 34356 13534
rect 34300 13470 34302 13522
rect 34354 13470 34356 13522
rect 34300 12962 34356 13470
rect 34300 12910 34302 12962
rect 34354 12910 34356 12962
rect 34300 12898 34356 12910
rect 34076 12686 34078 12738
rect 34130 12686 34132 12738
rect 34076 12674 34132 12686
rect 34524 12740 34580 12750
rect 34524 12646 34580 12684
rect 33404 11678 33406 11730
rect 33458 11678 33460 11730
rect 33068 10406 33124 10444
rect 32508 10388 32564 10398
rect 32508 9490 32564 10332
rect 32508 9438 32510 9490
rect 32562 9438 32564 9490
rect 32508 9426 32564 9438
rect 32732 9604 32788 9614
rect 32732 8594 32788 9548
rect 32732 8542 32734 8594
rect 32786 8542 32788 8594
rect 32732 8484 32788 8542
rect 32396 7422 32398 7474
rect 32450 7422 32452 7474
rect 31612 6468 31668 6478
rect 31388 6412 31612 6468
rect 29148 5796 29204 5806
rect 29820 5796 29876 6412
rect 29932 6402 29988 6412
rect 29204 5740 29316 5796
rect 29148 5730 29204 5740
rect 29260 5570 29316 5740
rect 29820 5730 29876 5740
rect 29260 5518 29262 5570
rect 29314 5518 29316 5570
rect 29260 5506 29316 5518
rect 31500 5458 31556 6412
rect 31612 6402 31668 6412
rect 31836 5570 31892 6524
rect 32396 6468 32452 7422
rect 32396 6402 32452 6412
rect 32508 7588 32564 7598
rect 32396 5796 32452 5806
rect 32508 5796 32564 7532
rect 32732 6692 32788 8428
rect 33292 8708 33348 8718
rect 33068 7588 33124 7598
rect 32844 7586 33124 7588
rect 32844 7534 33070 7586
rect 33122 7534 33124 7586
rect 32844 7532 33124 7534
rect 32844 6802 32900 7532
rect 33068 7522 33124 7532
rect 32844 6750 32846 6802
rect 32898 6750 32900 6802
rect 32844 6738 32900 6750
rect 32732 6626 32788 6636
rect 33068 6692 33124 6702
rect 32396 5794 32564 5796
rect 32396 5742 32398 5794
rect 32450 5742 32564 5794
rect 32396 5740 32564 5742
rect 32396 5730 32452 5740
rect 31836 5518 31838 5570
rect 31890 5518 31892 5570
rect 31836 5506 31892 5518
rect 33068 5572 33124 6636
rect 33292 6356 33348 8652
rect 33404 7698 33460 11678
rect 34076 11732 34132 11742
rect 34636 11732 34692 15092
rect 35196 15082 35460 15092
rect 34860 14868 34916 14878
rect 34748 14642 34804 14654
rect 34748 14590 34750 14642
rect 34802 14590 34804 14642
rect 34748 13636 34804 14590
rect 34748 13570 34804 13580
rect 34860 13634 34916 14812
rect 36428 14756 36484 14766
rect 36428 14662 36484 14700
rect 37100 14644 37156 14654
rect 37100 14550 37156 14588
rect 35644 14532 35700 14542
rect 35644 14438 35700 14476
rect 34860 13582 34862 13634
rect 34914 13582 34916 13634
rect 34860 13524 34916 13582
rect 34860 13458 34916 13468
rect 37212 14308 37268 15092
rect 35196 13132 35460 13142
rect 35252 13076 35300 13132
rect 35356 13076 35404 13132
rect 35196 13066 35460 13076
rect 36428 12852 36484 12862
rect 36428 12738 36484 12796
rect 36428 12686 36430 12738
rect 36482 12686 36484 12738
rect 36428 12674 36484 12686
rect 37100 12628 37156 12638
rect 37100 12534 37156 12572
rect 35868 11732 35924 11742
rect 33740 11618 33796 11630
rect 33740 11566 33742 11618
rect 33794 11566 33796 11618
rect 33740 10388 33796 11566
rect 34076 11618 34132 11676
rect 34076 11566 34078 11618
rect 34130 11566 34132 11618
rect 34076 11554 34132 11566
rect 34412 11730 34692 11732
rect 34412 11678 34638 11730
rect 34690 11678 34692 11730
rect 34412 11676 34692 11678
rect 33740 10322 33796 10332
rect 33404 7646 33406 7698
rect 33458 7646 33460 7698
rect 33404 7634 33460 7646
rect 33516 8148 33572 8158
rect 33516 6692 33572 8092
rect 34076 7812 34132 7822
rect 34076 7718 34132 7756
rect 34412 7700 34468 11676
rect 34636 11666 34692 11676
rect 35532 11730 35924 11732
rect 35532 11678 35870 11730
rect 35922 11678 35924 11730
rect 35532 11676 35924 11678
rect 35196 11620 35252 11630
rect 34748 11618 35252 11620
rect 34748 11566 35198 11618
rect 35250 11566 35252 11618
rect 34748 11564 35252 11566
rect 34748 10948 34804 11564
rect 35196 11554 35252 11564
rect 35196 11116 35460 11126
rect 35252 11060 35300 11116
rect 35356 11060 35404 11116
rect 35196 11050 35460 11060
rect 34524 10892 34804 10948
rect 34524 10386 34580 10892
rect 34524 10334 34526 10386
rect 34578 10334 34580 10386
rect 34524 10322 34580 10334
rect 34748 9604 34804 9614
rect 34748 9510 34804 9548
rect 35196 9492 35252 9502
rect 35084 9490 35252 9492
rect 35084 9438 35198 9490
rect 35250 9438 35252 9490
rect 35084 9436 35252 9438
rect 35084 8482 35140 9436
rect 35196 9426 35252 9436
rect 35196 9100 35460 9110
rect 35252 9044 35300 9100
rect 35356 9044 35404 9100
rect 35196 9034 35460 9044
rect 35532 8930 35588 11676
rect 35868 11666 35924 11676
rect 36092 9604 36148 9614
rect 36092 9510 36148 9548
rect 36540 9602 36596 9614
rect 36540 9550 36542 9602
rect 36594 9550 36596 9602
rect 35532 8878 35534 8930
rect 35586 8878 35588 8930
rect 35532 8866 35588 8878
rect 35644 9492 35700 9502
rect 35644 8708 35700 9436
rect 36540 9492 36596 9550
rect 36540 9426 36596 9436
rect 37212 9380 37268 14252
rect 37324 14644 37380 16606
rect 37548 15876 37604 18508
rect 37660 17554 37716 18620
rect 38332 18676 38388 20412
rect 38668 20356 38724 21422
rect 38668 19794 38724 20300
rect 38668 19742 38670 19794
rect 38722 19742 38724 19794
rect 38668 19730 38724 19742
rect 39116 21586 39172 21598
rect 39116 21534 39118 21586
rect 39170 21534 39172 21586
rect 39116 19684 39172 21534
rect 40012 21586 40068 21598
rect 40012 21534 40014 21586
rect 40066 21534 40068 21586
rect 40012 20356 40068 21534
rect 39116 19682 39508 19684
rect 39116 19630 39118 19682
rect 39170 19630 39508 19682
rect 39116 19628 39508 19630
rect 39116 19618 39172 19628
rect 38332 18610 38388 18620
rect 38892 19010 38948 19022
rect 38892 18958 38894 19010
rect 38946 18958 38948 19010
rect 38556 18564 38612 18574
rect 38892 18564 38948 18958
rect 38556 18470 38612 18508
rect 38668 18562 38948 18564
rect 38668 18510 38894 18562
rect 38946 18510 38948 18562
rect 38668 18508 38948 18510
rect 38108 18340 38164 18350
rect 38668 18340 38724 18508
rect 38892 18498 38948 18508
rect 39228 18898 39284 18910
rect 39228 18846 39230 18898
rect 39282 18846 39284 18898
rect 38108 17892 38164 18284
rect 38444 18284 38724 18340
rect 38444 17892 38500 18284
rect 38108 17890 38500 17892
rect 38108 17838 38110 17890
rect 38162 17838 38500 17890
rect 38108 17836 38500 17838
rect 38108 17826 38164 17836
rect 38444 17778 38500 17836
rect 38444 17726 38446 17778
rect 38498 17726 38500 17778
rect 38444 17714 38500 17726
rect 37660 17502 37662 17554
rect 37714 17502 37716 17554
rect 37660 16882 37716 17502
rect 39228 16996 39284 18846
rect 39340 18676 39396 18686
rect 39340 18582 39396 18620
rect 39452 18564 39508 19628
rect 40012 18898 40068 20300
rect 40348 20690 40404 20702
rect 40348 20638 40350 20690
rect 40402 20638 40404 20690
rect 40236 19460 40292 19470
rect 40236 19366 40292 19404
rect 40012 18846 40014 18898
rect 40066 18846 40068 18898
rect 40012 18834 40068 18846
rect 40236 19010 40292 19022
rect 40236 18958 40238 19010
rect 40290 18958 40292 19010
rect 40236 18788 40292 18958
rect 40348 18900 40404 20638
rect 40796 20468 40852 20478
rect 40908 20468 40964 22654
rect 41020 22596 41076 22606
rect 41020 21922 41076 22540
rect 41020 21870 41022 21922
rect 41074 21870 41076 21922
rect 41020 21858 41076 21870
rect 40796 20466 40964 20468
rect 40796 20414 40798 20466
rect 40850 20414 40964 20466
rect 40796 20412 40964 20414
rect 41020 21700 41076 21710
rect 40796 20356 40852 20412
rect 40796 20290 40852 20300
rect 40908 20244 40964 20254
rect 40908 19796 40964 20188
rect 40796 19794 40964 19796
rect 40796 19742 40910 19794
rect 40962 19742 40964 19794
rect 40796 19740 40964 19742
rect 40348 18844 40628 18900
rect 40236 18786 40404 18788
rect 40236 18734 40238 18786
rect 40290 18734 40404 18786
rect 40236 18732 40404 18734
rect 40236 18722 40292 18732
rect 39788 18564 39844 18574
rect 39452 18562 39844 18564
rect 39452 18510 39790 18562
rect 39842 18510 39844 18562
rect 39452 18508 39844 18510
rect 37660 16830 37662 16882
rect 37714 16830 37716 16882
rect 37660 16818 37716 16830
rect 38668 16940 39284 16996
rect 38668 16770 38724 16940
rect 38668 16718 38670 16770
rect 38722 16718 38724 16770
rect 38220 16660 38276 16670
rect 38220 16566 38276 16604
rect 37772 16548 37828 16558
rect 37828 16492 37940 16548
rect 37772 16454 37828 16492
rect 37772 15876 37828 15886
rect 37548 15874 37828 15876
rect 37548 15822 37774 15874
rect 37826 15822 37828 15874
rect 37548 15820 37828 15822
rect 37772 15810 37828 15820
rect 37436 15764 37492 15774
rect 37436 15670 37492 15708
rect 37884 15148 37940 16492
rect 37324 13860 37380 14588
rect 37772 15092 37940 15148
rect 37996 15764 38052 15774
rect 37772 14532 37828 15092
rect 37772 14466 37828 14476
rect 37884 14980 37940 14990
rect 37884 14642 37940 14924
rect 37884 14590 37886 14642
rect 37938 14590 37940 14642
rect 37324 13522 37380 13804
rect 37324 13470 37326 13522
rect 37378 13470 37380 13522
rect 37324 12628 37380 13470
rect 37884 12852 37940 14590
rect 37996 13970 38052 15708
rect 38332 15652 38388 15662
rect 38332 15558 38388 15596
rect 38668 14980 38724 16718
rect 39004 16770 39060 16782
rect 39004 16718 39006 16770
rect 39058 16718 39060 16770
rect 38668 14914 38724 14924
rect 38892 15650 38948 15662
rect 38892 15598 38894 15650
rect 38946 15598 38948 15650
rect 38220 14756 38276 14766
rect 38892 14756 38948 15598
rect 38276 14700 38948 14756
rect 38220 14662 38276 14700
rect 38556 14418 38612 14700
rect 39004 14532 39060 16718
rect 39228 16546 39284 16940
rect 39676 16772 39732 18508
rect 39788 18498 39844 18508
rect 39676 16706 39732 16716
rect 40348 18452 40404 18732
rect 40572 18674 40628 18844
rect 40572 18622 40574 18674
rect 40626 18622 40628 18674
rect 40572 18610 40628 18622
rect 40796 18452 40852 19740
rect 40908 19730 40964 19740
rect 40908 18564 40964 18574
rect 41020 18564 41076 21644
rect 41132 20188 41188 23436
rect 41244 22820 41300 23548
rect 41356 23714 41412 23884
rect 41356 23662 41358 23714
rect 41410 23662 41412 23714
rect 41356 23044 41412 23662
rect 41468 23716 41524 24108
rect 41468 23622 41524 23660
rect 41356 23042 41524 23044
rect 41356 22990 41358 23042
rect 41410 22990 41524 23042
rect 41356 22988 41524 22990
rect 41356 22978 41412 22988
rect 41356 22820 41412 22830
rect 41244 22818 41412 22820
rect 41244 22766 41358 22818
rect 41410 22766 41412 22818
rect 41244 22764 41412 22766
rect 41244 22596 41300 22764
rect 41244 22530 41300 22540
rect 41356 21924 41412 22764
rect 41356 20692 41412 21868
rect 41468 21922 41524 22988
rect 41468 21870 41470 21922
rect 41522 21870 41524 21922
rect 41468 21812 41524 21870
rect 41468 21746 41524 21756
rect 41580 21700 41636 33404
rect 41804 32564 41860 33628
rect 41916 33618 41972 33628
rect 42700 33684 42756 33694
rect 41692 32508 41804 32564
rect 41692 31890 41748 32508
rect 41804 32498 41860 32508
rect 41916 32900 41972 32910
rect 41916 32674 41972 32844
rect 41916 32622 41918 32674
rect 41970 32622 41972 32674
rect 41692 31838 41694 31890
rect 41746 31838 41748 31890
rect 41692 31108 41748 31838
rect 41692 31042 41748 31052
rect 41804 31892 41860 31902
rect 41804 30770 41860 31836
rect 41916 30884 41972 32622
rect 41916 30818 41972 30828
rect 42476 31442 42532 31454
rect 42476 31390 42478 31442
rect 42530 31390 42532 31442
rect 41804 30718 41806 30770
rect 41858 30718 41860 30770
rect 41804 30706 41860 30718
rect 41580 21634 41636 21644
rect 41692 29874 41748 29886
rect 41692 29822 41694 29874
rect 41746 29822 41748 29874
rect 41468 20692 41524 20702
rect 41356 20690 41524 20692
rect 41356 20638 41470 20690
rect 41522 20638 41524 20690
rect 41356 20636 41524 20638
rect 41468 20580 41524 20636
rect 41468 20514 41524 20524
rect 41580 20692 41636 20702
rect 41580 20244 41636 20636
rect 41132 20132 41524 20188
rect 41580 20178 41636 20188
rect 41356 19796 41412 19806
rect 41244 19460 41300 19470
rect 41244 18674 41300 19404
rect 41244 18622 41246 18674
rect 41298 18622 41300 18674
rect 41244 18610 41300 18622
rect 41356 18676 41412 19740
rect 41356 18610 41412 18620
rect 40964 18508 41076 18564
rect 40908 18470 40964 18508
rect 40348 18396 40796 18452
rect 40348 16658 40404 18396
rect 40796 18358 40852 18396
rect 40460 17332 40516 17342
rect 40460 17330 40852 17332
rect 40460 17278 40462 17330
rect 40514 17278 40852 17330
rect 40460 17276 40852 17278
rect 40460 17266 40516 17276
rect 40348 16606 40350 16658
rect 40402 16606 40404 16658
rect 39228 16494 39230 16546
rect 39282 16494 39284 16546
rect 39228 16482 39284 16494
rect 39452 16548 39508 16558
rect 39452 16454 39508 16492
rect 39900 16546 39956 16558
rect 39900 16494 39902 16546
rect 39954 16494 39956 16546
rect 39564 15764 39620 15774
rect 39564 15670 39620 15708
rect 39228 14756 39284 14766
rect 38556 14366 38558 14418
rect 38610 14366 38612 14418
rect 38556 14354 38612 14366
rect 38892 14530 39060 14532
rect 38892 14478 39006 14530
rect 39058 14478 39060 14530
rect 38892 14476 39060 14478
rect 37996 13918 37998 13970
rect 38050 13918 38052 13970
rect 37996 13906 38052 13918
rect 37884 12758 37940 12796
rect 38108 13636 38164 13646
rect 38108 12852 38164 13580
rect 38556 13524 38612 13534
rect 38892 13524 38948 14476
rect 39004 14466 39060 14476
rect 39116 14700 39228 14756
rect 39004 13860 39060 13870
rect 39116 13860 39172 14700
rect 39228 14690 39284 14700
rect 39676 14756 39732 14766
rect 39676 14642 39732 14700
rect 39676 14590 39678 14642
rect 39730 14590 39732 14642
rect 39676 14578 39732 14590
rect 39004 13858 39172 13860
rect 39004 13806 39006 13858
rect 39058 13806 39172 13858
rect 39004 13804 39172 13806
rect 39004 13794 39060 13804
rect 39004 13524 39060 13534
rect 38892 13468 39004 13524
rect 38556 13430 38612 13468
rect 39004 13458 39060 13468
rect 39900 13524 39956 16494
rect 40348 15874 40404 16606
rect 40796 15986 40852 17276
rect 40796 15934 40798 15986
rect 40850 15934 40852 15986
rect 40796 15922 40852 15934
rect 40348 15822 40350 15874
rect 40402 15822 40404 15874
rect 40236 14756 40292 14766
rect 40348 14756 40404 15822
rect 41020 15874 41076 18508
rect 41244 18452 41300 18462
rect 41300 18396 41412 18452
rect 41244 18386 41300 18396
rect 41356 17780 41412 18396
rect 41356 17686 41412 17724
rect 41132 15988 41188 15998
rect 41132 15986 41412 15988
rect 41132 15934 41134 15986
rect 41186 15934 41412 15986
rect 41132 15932 41412 15934
rect 41132 15922 41188 15932
rect 41020 15822 41022 15874
rect 41074 15822 41076 15874
rect 41020 15764 41076 15822
rect 41020 15698 41076 15708
rect 41356 15762 41412 15932
rect 41356 15710 41358 15762
rect 41410 15710 41412 15762
rect 41356 15698 41412 15710
rect 41468 15092 41524 20132
rect 41580 19348 41636 19358
rect 41580 18674 41636 19292
rect 41580 18622 41582 18674
rect 41634 18622 41636 18674
rect 41580 18610 41636 18622
rect 41692 15876 41748 29822
rect 42364 29876 42420 29886
rect 42476 29876 42532 31390
rect 42364 29874 42532 29876
rect 42364 29822 42366 29874
rect 42418 29822 42532 29874
rect 42364 29820 42532 29822
rect 42700 29876 42756 33628
rect 43148 33684 43204 33742
rect 43148 33618 43204 33628
rect 43260 32900 43316 34524
rect 43484 34578 43540 34590
rect 43484 34526 43486 34578
rect 43538 34526 43540 34578
rect 43484 33906 43540 34526
rect 43484 33854 43486 33906
rect 43538 33854 43540 33906
rect 43484 33842 43540 33854
rect 43260 32898 43428 32900
rect 43260 32846 43262 32898
rect 43314 32846 43428 32898
rect 43260 32844 43428 32846
rect 43260 32834 43316 32844
rect 42812 32786 42868 32798
rect 42812 32734 42814 32786
rect 42866 32734 42868 32786
rect 42812 32564 42868 32734
rect 42812 32498 42868 32508
rect 43260 32004 43316 32014
rect 42812 31892 42868 31902
rect 42812 31798 42868 31836
rect 43148 30548 43204 30558
rect 43036 30546 43204 30548
rect 43036 30494 43150 30546
rect 43202 30494 43204 30546
rect 43036 30492 43204 30494
rect 42700 29874 42868 29876
rect 42700 29822 42702 29874
rect 42754 29822 42868 29874
rect 42700 29820 42868 29822
rect 42364 29810 42420 29820
rect 42700 29810 42756 29820
rect 41804 27748 41860 27758
rect 42140 27748 42196 27758
rect 41804 27746 42196 27748
rect 41804 27694 41806 27746
rect 41858 27694 42142 27746
rect 42194 27694 42196 27746
rect 41804 27692 42196 27694
rect 41804 27682 41860 27692
rect 42140 26964 42196 27692
rect 42028 26852 42196 26908
rect 42700 27410 42756 27422
rect 42700 27358 42702 27410
rect 42754 27358 42756 27410
rect 42028 26850 42084 26852
rect 42028 26798 42030 26850
rect 42082 26798 42084 26850
rect 42028 26516 42084 26798
rect 42700 26738 42756 27358
rect 42700 26686 42702 26738
rect 42754 26686 42756 26738
rect 42700 26674 42756 26686
rect 42812 26740 42868 29820
rect 43036 29874 43092 30492
rect 43148 30482 43204 30492
rect 43036 29822 43038 29874
rect 43090 29822 43092 29874
rect 43036 29810 43092 29822
rect 42924 26740 42980 26750
rect 42812 26738 42980 26740
rect 42812 26686 42926 26738
rect 42978 26686 42980 26738
rect 42812 26684 42980 26686
rect 42924 26674 42980 26684
rect 42028 26450 42084 26460
rect 43148 26626 43204 26638
rect 43148 26574 43150 26626
rect 43202 26574 43204 26626
rect 42252 26402 42308 26414
rect 42252 26350 42254 26402
rect 42306 26350 42308 26402
rect 42252 25956 42308 26350
rect 43148 26066 43204 26574
rect 43148 26014 43150 26066
rect 43202 26014 43204 26066
rect 43148 26002 43204 26014
rect 42252 25890 42308 25900
rect 42364 24610 42420 24622
rect 42364 24558 42366 24610
rect 42418 24558 42420 24610
rect 42364 23940 42420 24558
rect 42028 23884 42420 23940
rect 41916 23604 41972 23614
rect 42028 23604 42084 23884
rect 42812 23828 42868 23838
rect 42812 23734 42868 23772
rect 42140 23716 42196 23726
rect 42196 23660 42308 23716
rect 42140 23650 42196 23660
rect 41916 23602 42084 23604
rect 41916 23550 41918 23602
rect 41970 23550 42084 23602
rect 41916 23548 42084 23550
rect 41804 23042 41860 23054
rect 41804 22990 41806 23042
rect 41858 22990 41860 23042
rect 41804 22818 41860 22990
rect 41916 22930 41972 23548
rect 41916 22878 41918 22930
rect 41970 22878 41972 22930
rect 41916 22866 41972 22878
rect 41804 22766 41806 22818
rect 41858 22766 41860 22818
rect 41804 22754 41860 22766
rect 42252 22820 42308 23660
rect 42700 22820 42756 22830
rect 42252 22818 42756 22820
rect 42252 22766 42254 22818
rect 42306 22766 42702 22818
rect 42754 22766 42756 22818
rect 42252 22764 42756 22766
rect 41916 21924 41972 21934
rect 41916 21830 41972 21868
rect 41804 21812 41860 21822
rect 41804 20578 41860 21756
rect 42252 20692 42308 22764
rect 42700 22754 42756 22764
rect 42364 21812 42420 21822
rect 42364 21718 42420 21756
rect 43036 21812 43092 21822
rect 43260 21812 43316 31948
rect 43372 31890 43428 32844
rect 43372 31838 43374 31890
rect 43426 31838 43428 31890
rect 43372 31826 43428 31838
rect 43484 32564 43540 32574
rect 43484 31778 43540 32508
rect 43484 31726 43486 31778
rect 43538 31726 43540 31778
rect 43484 31714 43540 31726
rect 43596 30884 43652 34860
rect 44268 34914 44324 36652
rect 44380 36036 44436 36046
rect 44380 35942 44436 35980
rect 44268 34862 44270 34914
rect 44322 34862 44324 34914
rect 44268 34804 44324 34862
rect 44268 34738 44324 34748
rect 44268 33906 44324 33918
rect 44268 33854 44270 33906
rect 44322 33854 44324 33906
rect 43820 33796 43876 33806
rect 43820 33702 43876 33740
rect 43708 32562 43764 32574
rect 43708 32510 43710 32562
rect 43762 32510 43764 32562
rect 43708 31892 43764 32510
rect 44156 32564 44212 32574
rect 44156 32470 44212 32508
rect 44044 31892 44100 31902
rect 43708 31836 44044 31892
rect 43820 31668 43876 31678
rect 43596 30882 43764 30884
rect 43596 30830 43598 30882
rect 43650 30830 43764 30882
rect 43596 30828 43764 30830
rect 43596 30818 43652 30828
rect 43708 30772 43764 30828
rect 43484 30100 43540 30110
rect 43372 29988 43428 29998
rect 43372 29894 43428 29932
rect 43372 28868 43428 28878
rect 43484 28868 43540 30044
rect 43372 28866 43540 28868
rect 43372 28814 43374 28866
rect 43426 28814 43540 28866
rect 43372 28812 43540 28814
rect 43708 28868 43764 30716
rect 43820 29874 43876 31612
rect 43932 30212 43988 31836
rect 44044 31798 44100 31836
rect 44268 31780 44324 33854
rect 44380 32004 44436 32014
rect 44492 32004 44548 37772
rect 44828 37828 44884 37884
rect 45948 37874 46004 37884
rect 46060 38498 46340 38500
rect 46060 38446 46286 38498
rect 46338 38446 46340 38498
rect 46060 38444 46340 38446
rect 44828 37762 44884 37772
rect 45276 37828 45332 37838
rect 45276 37734 45332 37772
rect 44940 37714 44996 37726
rect 44940 37662 44942 37714
rect 44994 37662 44996 37714
rect 44940 36820 44996 37662
rect 44940 36754 44996 36764
rect 45500 36706 45556 36718
rect 45500 36654 45502 36706
rect 45554 36654 45556 36706
rect 45052 36484 45108 36494
rect 45500 36484 45556 36654
rect 46060 36706 46116 38444
rect 46284 38434 46340 38444
rect 46844 37938 46900 39788
rect 47180 38724 47236 38734
rect 47180 38630 47236 38668
rect 47404 38722 47460 38734
rect 48300 38724 48356 38734
rect 47404 38670 47406 38722
rect 47458 38670 47460 38722
rect 47404 38668 47460 38670
rect 48188 38668 48300 38724
rect 47404 38612 47572 38668
rect 46844 37886 46846 37938
rect 46898 37886 46900 37938
rect 46844 37874 46900 37886
rect 47292 37940 47348 37950
rect 47292 37846 47348 37884
rect 47516 37714 47572 38612
rect 48188 38050 48244 38668
rect 48300 38658 48356 38668
rect 48188 37998 48190 38050
rect 48242 37998 48244 38050
rect 48188 37986 48244 37998
rect 47516 37662 47518 37714
rect 47570 37662 47572 37714
rect 46396 37492 46452 37502
rect 46284 37490 46452 37492
rect 46284 37438 46398 37490
rect 46450 37438 46452 37490
rect 46284 37436 46452 37438
rect 46172 36820 46228 36830
rect 46172 36726 46228 36764
rect 46060 36654 46062 36706
rect 46114 36654 46116 36706
rect 46060 36642 46116 36654
rect 46284 36484 46340 37436
rect 46396 37426 46452 37436
rect 47180 36820 47236 36830
rect 46732 36708 46788 36718
rect 47068 36708 47124 36718
rect 46788 36706 47124 36708
rect 46788 36654 47070 36706
rect 47122 36654 47124 36706
rect 46788 36652 47124 36654
rect 46732 36614 46788 36652
rect 47068 36642 47124 36652
rect 45052 36482 45220 36484
rect 45052 36430 45054 36482
rect 45106 36430 45220 36482
rect 45052 36428 45220 36430
rect 45500 36428 46340 36484
rect 45052 36418 45108 36428
rect 44828 36036 44884 36046
rect 44828 35942 44884 35980
rect 45052 34692 45108 34702
rect 45052 34598 45108 34636
rect 44436 31948 44548 32004
rect 44828 33908 44884 33918
rect 44380 31910 44436 31948
rect 44268 31714 44324 31724
rect 44044 30884 44100 30894
rect 44100 30828 44324 30884
rect 44044 30790 44100 30828
rect 43932 30146 43988 30156
rect 43820 29822 43822 29874
rect 43874 29822 43876 29874
rect 43820 29810 43876 29822
rect 43820 28868 43876 28878
rect 43708 28866 43876 28868
rect 43708 28814 43822 28866
rect 43874 28814 43876 28866
rect 43708 28812 43876 28814
rect 43372 28802 43428 28812
rect 43820 28802 43876 28812
rect 44268 28866 44324 30828
rect 44492 29764 44548 29774
rect 44492 29670 44548 29708
rect 44268 28814 44270 28866
rect 44322 28814 44324 28866
rect 44268 28802 44324 28814
rect 44828 28644 44884 33852
rect 44940 33794 44996 33806
rect 44940 33742 44942 33794
rect 44994 33742 44996 33794
rect 44940 33012 44996 33742
rect 45164 33124 45220 36428
rect 45612 36036 45668 36046
rect 45612 35942 45668 35980
rect 46732 36036 46788 36046
rect 46396 35812 46452 35822
rect 46396 34914 46452 35756
rect 46396 34862 46398 34914
rect 46450 34862 46452 34914
rect 46396 34850 46452 34862
rect 45164 33058 45220 33068
rect 45500 34804 45556 34814
rect 44940 32946 44996 32956
rect 45500 32900 45556 34748
rect 46620 34804 46676 34814
rect 46620 34130 46676 34748
rect 46620 34078 46622 34130
rect 46674 34078 46676 34130
rect 46620 34066 46676 34078
rect 45612 33908 45668 33918
rect 46284 33908 46340 33918
rect 45612 33906 45780 33908
rect 45612 33854 45614 33906
rect 45666 33854 45780 33906
rect 45612 33852 45780 33854
rect 45612 33842 45668 33852
rect 45612 32900 45668 32910
rect 45388 32898 45668 32900
rect 45388 32846 45614 32898
rect 45666 32846 45668 32898
rect 45388 32844 45668 32846
rect 45164 32564 45220 32574
rect 45164 31780 45220 32508
rect 45388 31892 45444 32844
rect 45612 32834 45668 32844
rect 45164 31714 45220 31724
rect 45276 31890 45444 31892
rect 45276 31838 45390 31890
rect 45442 31838 45444 31890
rect 45276 31836 45444 31838
rect 44940 31668 44996 31678
rect 44940 30770 44996 31612
rect 45276 31556 45332 31836
rect 45388 31826 45444 31836
rect 45388 31668 45444 31678
rect 45388 31574 45444 31612
rect 44940 30718 44942 30770
rect 44994 30718 44996 30770
rect 44940 30706 44996 30718
rect 45164 31500 45332 31556
rect 45724 31554 45780 33852
rect 46284 33814 46340 33852
rect 46060 33012 46116 33022
rect 46060 32918 46116 32956
rect 46620 32788 46676 32798
rect 46732 32788 46788 35980
rect 47068 33908 47124 33918
rect 47068 33814 47124 33852
rect 47180 33684 47236 36764
rect 47516 34804 47572 37662
rect 48188 36820 48244 36830
rect 47516 34738 47572 34748
rect 47740 36708 47796 36718
rect 47740 36036 47796 36652
rect 47740 34802 47796 35980
rect 47740 34750 47742 34802
rect 47794 34750 47796 34802
rect 47740 34738 47796 34750
rect 47516 33908 47572 33918
rect 48188 33908 48244 36764
rect 48300 36036 48356 36046
rect 48748 36036 48804 39900
rect 49196 39956 49252 39966
rect 49196 39862 49252 39900
rect 49308 38162 49364 42028
rect 49420 41858 49476 42588
rect 49532 42578 49588 42588
rect 50876 42642 50932 42654
rect 50876 42590 50878 42642
rect 50930 42590 50932 42642
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 49420 41806 49422 41858
rect 49474 41806 49476 41858
rect 49420 41636 49476 41806
rect 49420 41570 49476 41580
rect 49756 42196 49812 42206
rect 49756 41858 49812 42140
rect 49756 41806 49758 41858
rect 49810 41806 49812 41858
rect 49420 40516 49476 40526
rect 49420 40514 49588 40516
rect 49420 40462 49422 40514
rect 49474 40462 49588 40514
rect 49420 40460 49588 40462
rect 49420 40450 49476 40460
rect 49532 39954 49588 40460
rect 49532 39902 49534 39954
rect 49586 39902 49588 39954
rect 49532 39890 49588 39902
rect 49756 38612 49812 41806
rect 49868 42084 49924 42094
rect 49868 41858 49924 42028
rect 50876 41972 50932 42590
rect 51212 42642 51268 42654
rect 51212 42590 51214 42642
rect 51266 42590 51268 42642
rect 50932 41916 51044 41972
rect 50876 41906 50932 41916
rect 49868 41806 49870 41858
rect 49922 41806 49924 41858
rect 49868 41794 49924 41806
rect 50876 41748 50932 41758
rect 50316 41636 50372 41646
rect 50204 41634 50372 41636
rect 50204 41582 50318 41634
rect 50370 41582 50372 41634
rect 50204 41580 50372 41582
rect 49868 39956 49924 39966
rect 49868 39862 49924 39900
rect 50204 39954 50260 41580
rect 50316 41570 50372 41580
rect 50556 40348 50820 40358
rect 50612 40292 50660 40348
rect 50716 40292 50764 40348
rect 50556 40282 50820 40292
rect 50204 39902 50206 39954
rect 50258 39902 50260 39954
rect 50204 39890 50260 39902
rect 50540 39844 50596 39854
rect 50540 39750 50596 39788
rect 50876 38948 50932 41692
rect 50988 39956 51044 41916
rect 50988 39890 51044 39900
rect 51100 41860 51156 41870
rect 51100 39956 51156 41804
rect 51212 41748 51268 42590
rect 51660 42644 51716 42654
rect 51660 42084 51716 42588
rect 51660 42018 51716 42028
rect 51548 41748 51604 41758
rect 51268 41746 51604 41748
rect 51268 41694 51550 41746
rect 51602 41694 51604 41746
rect 51268 41692 51604 41694
rect 51212 41682 51268 41692
rect 51548 41682 51604 41692
rect 51660 39956 51716 39966
rect 51772 39956 51828 43710
rect 54124 43708 54180 43822
rect 54124 43652 54292 43708
rect 52108 42642 52164 42654
rect 52108 42590 52110 42642
rect 52162 42590 52164 42642
rect 52108 42196 52164 42590
rect 52108 42130 52164 42140
rect 52780 42642 52836 42654
rect 53340 42644 53396 42654
rect 52780 42590 52782 42642
rect 52834 42590 52836 42642
rect 51100 39954 51268 39956
rect 51100 39902 51102 39954
rect 51154 39902 51268 39954
rect 51100 39900 51268 39902
rect 51100 39890 51156 39900
rect 50428 38946 50932 38948
rect 50428 38894 50878 38946
rect 50930 38894 50932 38946
rect 50428 38892 50932 38894
rect 50428 38836 50484 38892
rect 50876 38882 50932 38892
rect 50316 38780 50484 38836
rect 49980 38612 50036 38622
rect 49756 38610 50036 38612
rect 49756 38558 49982 38610
rect 50034 38558 50036 38610
rect 49756 38556 50036 38558
rect 49308 38110 49310 38162
rect 49362 38110 49364 38162
rect 49308 38050 49364 38110
rect 49308 37998 49310 38050
rect 49362 37998 49364 38050
rect 49308 37986 49364 37998
rect 49644 38162 49700 38174
rect 49644 38110 49646 38162
rect 49698 38110 49700 38162
rect 48860 37716 48916 37726
rect 48860 37622 48916 37660
rect 49644 36818 49700 38110
rect 49756 37716 49812 38556
rect 49980 38498 50036 38556
rect 49980 38446 49982 38498
rect 50034 38446 50036 38498
rect 49980 38434 50036 38446
rect 50204 38052 50260 38062
rect 50316 38052 50372 38780
rect 50540 38724 50596 38734
rect 50204 38050 50372 38052
rect 50204 37998 50206 38050
rect 50258 37998 50372 38050
rect 50204 37996 50372 37998
rect 50428 38668 50540 38724
rect 50428 38610 50484 38668
rect 50540 38658 50596 38668
rect 50428 38558 50430 38610
rect 50482 38558 50484 38610
rect 50092 37716 50148 37726
rect 49756 37714 49924 37716
rect 49756 37662 49758 37714
rect 49810 37662 49924 37714
rect 49756 37660 49924 37662
rect 49756 37650 49812 37660
rect 49644 36766 49646 36818
rect 49698 36766 49700 36818
rect 49644 36754 49700 36766
rect 49756 37490 49812 37502
rect 49756 37438 49758 37490
rect 49810 37438 49812 37490
rect 49756 36708 49812 37438
rect 49868 36818 49924 37660
rect 49868 36766 49870 36818
rect 49922 36766 49924 36818
rect 49868 36754 49924 36766
rect 50092 36818 50148 37660
rect 50204 37490 50260 37996
rect 50204 37438 50206 37490
rect 50258 37438 50260 37490
rect 50204 37426 50260 37438
rect 50428 37156 50484 38558
rect 50556 38332 50820 38342
rect 50612 38276 50660 38332
rect 50716 38276 50764 38332
rect 50556 38266 50820 38276
rect 50652 38162 50708 38174
rect 50652 38110 50654 38162
rect 50706 38110 50708 38162
rect 50652 38050 50708 38110
rect 50652 37998 50654 38050
rect 50706 37998 50708 38050
rect 50652 37986 50708 37998
rect 51100 37714 51156 37726
rect 51100 37662 51102 37714
rect 51154 37662 51156 37714
rect 51100 37602 51156 37662
rect 51100 37550 51102 37602
rect 51154 37550 51156 37602
rect 51100 37538 51156 37550
rect 50316 37100 50484 37156
rect 50092 36766 50094 36818
rect 50146 36766 50148 36818
rect 49756 36642 49812 36652
rect 48860 36484 48916 36494
rect 48860 36482 49476 36484
rect 48860 36430 48862 36482
rect 48914 36430 49476 36482
rect 48860 36428 49476 36430
rect 48860 36418 48916 36428
rect 48300 36034 49140 36036
rect 48300 35982 48302 36034
rect 48354 35982 49140 36034
rect 48300 35980 49140 35982
rect 48300 35970 48356 35980
rect 49084 35922 49140 35980
rect 49084 35870 49086 35922
rect 49138 35870 49140 35922
rect 49084 35858 49140 35870
rect 49420 35922 49476 36428
rect 49420 35870 49422 35922
rect 49474 35870 49476 35922
rect 49420 35858 49476 35870
rect 48748 35812 48804 35822
rect 48748 35718 48804 35756
rect 49756 35810 49812 35822
rect 49756 35758 49758 35810
rect 49810 35758 49812 35810
rect 49644 34804 49700 34842
rect 49644 34738 49700 34748
rect 48524 34690 48580 34702
rect 48524 34638 48526 34690
rect 48578 34638 48580 34690
rect 48524 33908 48580 34638
rect 49308 34692 49364 34702
rect 47516 33906 48580 33908
rect 47516 33854 47518 33906
rect 47570 33854 48580 33906
rect 47516 33852 48580 33854
rect 47516 33842 47572 33852
rect 47180 33618 47236 33628
rect 48188 33684 48244 33694
rect 48524 33684 48580 33852
rect 49084 34468 49140 34478
rect 49084 33906 49140 34412
rect 49084 33854 49086 33906
rect 49138 33854 49140 33906
rect 49084 33842 49140 33854
rect 48524 33628 48804 33684
rect 46620 32786 46788 32788
rect 46620 32734 46622 32786
rect 46674 32734 46788 32786
rect 46620 32732 46788 32734
rect 46620 32722 46676 32732
rect 46620 31890 46676 31902
rect 46620 31838 46622 31890
rect 46674 31838 46676 31890
rect 45724 31502 45726 31554
rect 45778 31502 45780 31554
rect 45164 30770 45220 31500
rect 45724 31490 45780 31502
rect 46396 31780 46452 31790
rect 45276 30884 45332 30894
rect 45332 30828 45444 30884
rect 45276 30818 45332 30828
rect 45164 30718 45166 30770
rect 45218 30718 45220 30770
rect 45164 30706 45220 30718
rect 45388 30770 45444 30828
rect 45388 30718 45390 30770
rect 45442 30718 45444 30770
rect 45388 30706 45444 30718
rect 45612 30882 45668 30894
rect 45612 30830 45614 30882
rect 45666 30830 45668 30882
rect 45612 30658 45668 30830
rect 46396 30882 46452 31724
rect 46396 30830 46398 30882
rect 46450 30830 46452 30882
rect 46396 30818 46452 30830
rect 46620 30884 46676 31838
rect 46620 30818 46676 30828
rect 46732 31668 46788 32732
rect 46956 32674 47012 32686
rect 46956 32622 46958 32674
rect 47010 32622 47012 32674
rect 46956 31780 47012 32622
rect 47180 31892 47236 31902
rect 47180 31798 47236 31836
rect 47516 31892 47572 31902
rect 46956 31714 47012 31724
rect 45948 30772 46004 30782
rect 46172 30772 46228 30782
rect 45948 30678 46004 30716
rect 46060 30770 46228 30772
rect 46060 30718 46174 30770
rect 46226 30718 46228 30770
rect 46060 30716 46228 30718
rect 45612 30606 45614 30658
rect 45666 30606 45668 30658
rect 45052 30548 45108 30558
rect 45052 30546 45220 30548
rect 45052 30494 45054 30546
rect 45106 30494 45220 30546
rect 45052 30492 45220 30494
rect 45052 30482 45108 30492
rect 45164 29986 45220 30492
rect 45164 29934 45166 29986
rect 45218 29934 45220 29986
rect 45164 29922 45220 29934
rect 45612 28756 45668 30606
rect 46060 30100 46116 30716
rect 46172 30706 46228 30716
rect 46620 30660 46676 30670
rect 46732 30660 46788 31612
rect 46844 31666 46900 31678
rect 46844 31614 46846 31666
rect 46898 31614 46900 31666
rect 46844 30772 46900 31614
rect 47516 31666 47572 31836
rect 47964 31780 48020 31790
rect 47964 31686 48020 31724
rect 47516 31614 47518 31666
rect 47570 31614 47572 31666
rect 47516 31602 47572 31614
rect 46844 30706 46900 30716
rect 44828 28642 45108 28644
rect 44828 28590 44830 28642
rect 44882 28590 45108 28642
rect 44828 28588 45108 28590
rect 44828 28578 44884 28588
rect 45052 27972 45108 28588
rect 45164 28532 45220 28542
rect 45220 28476 45332 28532
rect 45164 28438 45220 28476
rect 45164 27972 45220 27982
rect 45052 27970 45220 27972
rect 45052 27918 45166 27970
rect 45218 27918 45220 27970
rect 45052 27916 45220 27918
rect 45164 27906 45220 27916
rect 45276 27860 45332 28476
rect 45612 27970 45668 28700
rect 45948 29650 46004 29662
rect 45948 29598 45950 29650
rect 46002 29598 46004 29650
rect 45948 28756 46004 29598
rect 45948 28690 46004 28700
rect 46060 28644 46116 30044
rect 46396 30658 46788 30660
rect 46396 30606 46622 30658
rect 46674 30606 46788 30658
rect 46396 30604 46788 30606
rect 46396 29986 46452 30604
rect 46620 30594 46676 30604
rect 46396 29934 46398 29986
rect 46450 29934 46452 29986
rect 46396 29922 46452 29934
rect 46172 29764 46228 29774
rect 46172 28866 46228 29708
rect 46172 28814 46174 28866
rect 46226 28814 46228 28866
rect 46172 28802 46228 28814
rect 46508 28980 46564 28990
rect 46060 28588 46228 28644
rect 45612 27918 45614 27970
rect 45666 27918 45668 27970
rect 45612 27906 45668 27918
rect 45276 27794 45332 27804
rect 46060 27636 46116 27646
rect 43932 26514 43988 26526
rect 43932 26462 43934 26514
rect 43986 26462 43988 26514
rect 43932 26404 43988 26462
rect 43596 24610 43652 24622
rect 43596 24558 43598 24610
rect 43650 24558 43652 24610
rect 43596 23604 43652 24558
rect 43932 23940 43988 26348
rect 43932 23874 43988 23884
rect 44828 26516 44884 26526
rect 44828 25730 44884 26460
rect 45500 26516 45556 26526
rect 45500 26422 45556 26460
rect 45836 26180 45892 26190
rect 45836 26066 45892 26124
rect 45836 26014 45838 26066
rect 45890 26014 45892 26066
rect 45836 26002 45892 26014
rect 44828 25678 44830 25730
rect 44882 25678 44884 25730
rect 44828 23940 44884 25678
rect 45948 25620 46004 25630
rect 45724 25564 45948 25620
rect 45724 24834 45780 25564
rect 45948 25554 46004 25564
rect 45724 24782 45726 24834
rect 45778 24782 45780 24834
rect 45724 24770 45780 24782
rect 44828 23846 44884 23884
rect 45276 24052 45332 24062
rect 45276 23938 45332 23996
rect 45276 23886 45278 23938
rect 45330 23886 45332 23938
rect 43596 23538 43652 23548
rect 45276 23604 45332 23886
rect 45724 23828 45780 23838
rect 45724 23734 45780 23772
rect 46060 23828 46116 27580
rect 46172 25956 46228 28588
rect 46172 25890 46228 25900
rect 46284 25732 46340 25742
rect 46284 25638 46340 25676
rect 46508 25730 46564 28924
rect 46732 28756 46788 30604
rect 47068 30546 47124 30558
rect 47068 30494 47070 30546
rect 47122 30494 47124 30546
rect 46844 28756 46900 28766
rect 46732 28754 46900 28756
rect 46732 28702 46846 28754
rect 46898 28702 46900 28754
rect 46732 28700 46900 28702
rect 46844 28690 46900 28700
rect 47068 28532 47124 30494
rect 48188 29652 48244 33628
rect 48636 33458 48692 33470
rect 48636 33406 48638 33458
rect 48690 33406 48692 33458
rect 48636 32788 48692 33406
rect 48748 32788 48804 33628
rect 48972 32788 49028 32798
rect 48748 32786 49028 32788
rect 48748 32734 48974 32786
rect 49026 32734 49028 32786
rect 48748 32732 49028 32734
rect 48636 32722 48692 32732
rect 48748 31556 48804 31566
rect 48804 31500 48916 31556
rect 48748 31490 48804 31500
rect 48748 30660 48804 30670
rect 48300 30548 48356 30558
rect 48300 30454 48356 30492
rect 48748 30546 48804 30604
rect 48748 30494 48750 30546
rect 48802 30494 48804 30546
rect 48636 30436 48692 30446
rect 48636 30098 48692 30380
rect 48636 30046 48638 30098
rect 48690 30046 48692 30098
rect 48636 30034 48692 30046
rect 48188 29558 48244 29596
rect 48188 28756 48244 28766
rect 48188 28642 48244 28700
rect 48188 28590 48190 28642
rect 48242 28590 48244 28642
rect 48188 28578 48244 28590
rect 48748 28644 48804 30494
rect 48748 28578 48804 28588
rect 47068 28466 47124 28476
rect 47740 28532 47796 28542
rect 46620 27860 46676 27870
rect 46620 27766 46676 27804
rect 47740 27636 47796 28476
rect 48300 27860 48356 27870
rect 48748 27860 48804 27870
rect 48860 27860 48916 31500
rect 48972 30660 49028 32732
rect 49308 32786 49364 34636
rect 49756 34690 49812 35758
rect 50092 35812 50148 36766
rect 50204 36932 50260 36942
rect 50204 35924 50260 36876
rect 50316 36820 50372 37100
rect 50428 36932 50484 36942
rect 51212 36932 51268 39900
rect 51660 39954 51828 39956
rect 51660 39902 51662 39954
rect 51714 39902 51828 39954
rect 51660 39900 51828 39902
rect 51996 42084 52052 42094
rect 51996 41746 52052 42028
rect 51996 41694 51998 41746
rect 52050 41694 52052 41746
rect 51996 41636 52052 41694
rect 51660 39890 51716 39900
rect 51996 39844 52052 41580
rect 52332 42082 52388 42094
rect 52332 42030 52334 42082
rect 52386 42030 52388 42082
rect 52332 40066 52388 42030
rect 52780 42084 52836 42590
rect 52780 42018 52836 42028
rect 53228 42588 53340 42644
rect 53116 41972 53172 41982
rect 53116 41878 53172 41916
rect 52332 40014 52334 40066
rect 52386 40014 52388 40066
rect 52332 40002 52388 40014
rect 52780 41858 52836 41870
rect 52780 41806 52782 41858
rect 52834 41806 52836 41858
rect 52780 40068 52836 41806
rect 53228 40850 53284 42588
rect 53340 42550 53396 42588
rect 53788 42642 53844 42654
rect 53788 42590 53790 42642
rect 53842 42590 53844 42642
rect 53788 42196 53844 42590
rect 53788 42130 53844 42140
rect 54236 42642 54292 43652
rect 54236 42590 54238 42642
rect 54290 42590 54292 42642
rect 53452 41860 53508 41870
rect 53340 41858 53508 41860
rect 53340 41806 53454 41858
rect 53506 41806 53508 41858
rect 53340 41804 53508 41806
rect 53340 41186 53396 41804
rect 53452 41794 53508 41804
rect 53788 41858 53844 41870
rect 53788 41806 53790 41858
rect 53842 41806 53844 41858
rect 53340 41134 53342 41186
rect 53394 41134 53396 41186
rect 53340 41122 53396 41134
rect 53228 40798 53230 40850
rect 53282 40798 53284 40850
rect 53228 40786 53284 40798
rect 53788 40180 53844 41806
rect 54236 41076 54292 42590
rect 55580 41970 55636 41982
rect 55580 41918 55582 41970
rect 55634 41918 55636 41970
rect 54348 41860 54404 41870
rect 54348 41766 54404 41804
rect 54908 41858 54964 41870
rect 54908 41806 54910 41858
rect 54962 41806 54964 41858
rect 54236 41020 54628 41076
rect 53788 40114 53844 40124
rect 54460 40850 54516 40862
rect 54460 40798 54462 40850
rect 54514 40798 54516 40850
rect 53116 40068 53172 40078
rect 52780 40066 53172 40068
rect 52780 40014 53118 40066
rect 53170 40014 53172 40066
rect 52780 40012 53172 40014
rect 53116 40002 53172 40012
rect 53228 39956 53284 39966
rect 53004 39844 53060 39854
rect 51772 39788 51996 39844
rect 51772 38946 51828 39788
rect 51996 39778 52052 39788
rect 52780 39788 53004 39844
rect 51772 38894 51774 38946
rect 51826 38894 51828 38946
rect 51772 38724 51828 38894
rect 51772 38658 51828 38668
rect 52780 38946 52836 39788
rect 53004 39750 53060 39788
rect 52780 38894 52782 38946
rect 52834 38894 52836 38946
rect 51324 38610 51380 38622
rect 51324 38558 51326 38610
rect 51378 38558 51380 38610
rect 51324 38498 51380 38558
rect 51324 38446 51326 38498
rect 51378 38446 51380 38498
rect 51324 37602 51380 38446
rect 52556 38498 52612 38510
rect 52556 38446 52558 38498
rect 52610 38446 52612 38498
rect 51660 38162 51716 38174
rect 51660 38110 51662 38162
rect 51714 38110 51716 38162
rect 51548 37828 51604 37838
rect 51548 37734 51604 37772
rect 51324 37550 51326 37602
rect 51378 37550 51380 37602
rect 51324 37044 51380 37550
rect 51436 37044 51492 37054
rect 51324 36988 51436 37044
rect 50428 36930 50708 36932
rect 50428 36878 50430 36930
rect 50482 36878 50708 36930
rect 50428 36876 50708 36878
rect 50428 36866 50484 36876
rect 50316 36726 50372 36764
rect 50652 36818 50708 36876
rect 51212 36866 51268 36876
rect 50652 36766 50654 36818
rect 50706 36766 50708 36818
rect 50652 36754 50708 36766
rect 51324 36820 51380 36830
rect 50540 36708 50596 36718
rect 50540 36614 50596 36652
rect 50876 36708 50932 36718
rect 51212 36708 51268 36718
rect 51324 36708 51380 36764
rect 51436 36818 51492 36988
rect 51436 36766 51438 36818
rect 51490 36766 51492 36818
rect 51436 36754 51492 36766
rect 51548 36930 51604 36942
rect 51548 36878 51550 36930
rect 51602 36878 51604 36930
rect 50932 36652 51156 36708
rect 50876 36614 50932 36652
rect 50556 36316 50820 36326
rect 50612 36260 50660 36316
rect 50716 36260 50764 36316
rect 50556 36250 50820 36260
rect 50316 35924 50372 35934
rect 50204 35922 50484 35924
rect 50204 35870 50318 35922
rect 50370 35870 50484 35922
rect 50204 35868 50484 35870
rect 50316 35830 50372 35868
rect 50092 35746 50148 35756
rect 49756 34638 49758 34690
rect 49810 34638 49812 34690
rect 49756 34626 49812 34638
rect 50316 34690 50372 34702
rect 50316 34638 50318 34690
rect 50370 34638 50372 34690
rect 49644 34580 49700 34590
rect 49644 33906 49700 34524
rect 49644 33854 49646 33906
rect 49698 33854 49700 33906
rect 49644 33842 49700 33854
rect 49420 33794 49476 33806
rect 49420 33742 49422 33794
rect 49474 33742 49476 33794
rect 49420 33684 49476 33742
rect 49420 33618 49476 33628
rect 50204 33794 50260 33806
rect 50204 33742 50206 33794
rect 50258 33742 50260 33794
rect 49308 32734 49310 32786
rect 49362 32734 49364 32786
rect 49308 32722 49364 32734
rect 49420 31892 49476 31902
rect 48972 30594 49028 30604
rect 49308 30660 49364 30670
rect 49308 30566 49364 30604
rect 49084 29764 49140 29774
rect 49084 29762 49252 29764
rect 49084 29710 49086 29762
rect 49138 29710 49252 29762
rect 49084 29708 49252 29710
rect 49084 29698 49140 29708
rect 49084 28754 49140 28766
rect 49084 28702 49086 28754
rect 49138 28702 49140 28754
rect 49084 28644 49140 28702
rect 49084 28578 49140 28588
rect 48300 27858 48916 27860
rect 48300 27806 48302 27858
rect 48354 27806 48750 27858
rect 48802 27806 48916 27858
rect 48300 27804 48916 27806
rect 48300 27794 48356 27804
rect 48748 27794 48804 27804
rect 47740 27542 47796 27580
rect 49084 27636 49140 27646
rect 46956 27524 47012 27534
rect 46956 27430 47012 27468
rect 48412 27524 48468 27534
rect 46508 25678 46510 25730
rect 46562 25678 46564 25730
rect 46508 25620 46564 25678
rect 46508 25554 46564 25564
rect 46732 27412 46788 27422
rect 46060 23762 46116 23772
rect 45276 23538 45332 23548
rect 46620 23378 46676 23390
rect 46620 23326 46622 23378
rect 46674 23326 46676 23378
rect 46620 22706 46676 23326
rect 46620 22654 46622 22706
rect 46674 22654 46676 22706
rect 46620 22642 46676 22654
rect 46732 22708 46788 27356
rect 46844 25842 46900 25854
rect 46844 25790 46846 25842
rect 46898 25790 46900 25842
rect 46844 25172 46900 25790
rect 46844 25116 47460 25172
rect 47404 25058 47460 25116
rect 47404 25006 47406 25058
rect 47458 25006 47460 25058
rect 47404 24994 47460 25006
rect 48412 24836 48468 27468
rect 49084 27522 49140 27580
rect 49084 27470 49086 27522
rect 49138 27470 49140 27522
rect 49084 27412 49140 27470
rect 49084 27346 49140 27356
rect 48860 27074 48916 27086
rect 48860 27022 48862 27074
rect 48914 27022 48916 27074
rect 48860 26738 48916 27022
rect 48860 26686 48862 26738
rect 48914 26686 48916 26738
rect 48860 26674 48916 26686
rect 48412 24722 48468 24780
rect 48412 24670 48414 24722
rect 48466 24670 48468 24722
rect 48412 24658 48468 24670
rect 48524 26404 48580 26414
rect 47852 24612 47908 24622
rect 48300 24612 48356 24622
rect 47404 24610 47908 24612
rect 47404 24558 47854 24610
rect 47906 24558 47908 24610
rect 47404 24556 47908 24558
rect 46844 23828 46900 23838
rect 47068 23828 47124 23838
rect 46900 23826 47124 23828
rect 46900 23774 47070 23826
rect 47122 23774 47124 23826
rect 46900 23772 47124 23774
rect 46844 23762 46900 23772
rect 47068 23762 47124 23772
rect 46956 22708 47012 22718
rect 46732 22706 47012 22708
rect 46732 22654 46958 22706
rect 47010 22654 47012 22706
rect 46732 22652 47012 22654
rect 46956 22642 47012 22652
rect 47292 22594 47348 22606
rect 47292 22542 47294 22594
rect 47346 22542 47348 22594
rect 47292 21922 47348 22542
rect 47292 21870 47294 21922
rect 47346 21870 47348 21922
rect 47292 21858 47348 21870
rect 43596 21812 43652 21822
rect 43036 21810 43652 21812
rect 43036 21758 43038 21810
rect 43090 21758 43598 21810
rect 43650 21758 43652 21810
rect 43036 21756 43652 21758
rect 43036 21746 43092 21756
rect 43596 21746 43652 21756
rect 45052 21810 45108 21822
rect 45052 21758 45054 21810
rect 45106 21758 45108 21810
rect 44604 21700 44660 21710
rect 44604 21606 44660 21644
rect 45052 21700 45108 21758
rect 45052 21634 45108 21644
rect 45164 21698 45220 21710
rect 45388 21700 45444 21710
rect 45164 21646 45166 21698
rect 45218 21646 45220 21698
rect 44156 21588 44212 21598
rect 42700 21476 42756 21486
rect 42252 20626 42308 20636
rect 42476 21474 42756 21476
rect 42476 21422 42702 21474
rect 42754 21422 42756 21474
rect 42476 21420 42756 21422
rect 41804 20526 41806 20578
rect 41858 20526 41860 20578
rect 41804 19796 41860 20526
rect 41804 19730 41860 19740
rect 42140 18564 42196 18574
rect 42476 18564 42532 21420
rect 42700 21410 42756 21420
rect 42700 20578 42756 20590
rect 42700 20526 42702 20578
rect 42754 20526 42756 20578
rect 42700 20356 42756 20526
rect 43484 20580 43540 20590
rect 42700 20290 42756 20300
rect 43372 20468 43428 20478
rect 42700 19460 42756 19470
rect 42700 18674 42756 19404
rect 42700 18622 42702 18674
rect 42754 18622 42756 18674
rect 42700 18610 42756 18622
rect 42140 18562 42532 18564
rect 42140 18510 42142 18562
rect 42194 18510 42532 18562
rect 42140 18508 42532 18510
rect 43372 18562 43428 20412
rect 43484 20244 43540 20524
rect 43596 20468 43652 20478
rect 43708 20468 43764 20478
rect 43652 20466 43764 20468
rect 43652 20414 43710 20466
rect 43762 20414 43764 20466
rect 43652 20412 43764 20414
rect 43596 20402 43652 20412
rect 43708 20402 43764 20412
rect 43484 19794 43540 20188
rect 44156 20244 44212 21532
rect 45164 21588 45220 21646
rect 45164 21522 45220 21532
rect 45276 21698 45444 21700
rect 45276 21646 45390 21698
rect 45442 21646 45444 21698
rect 45276 21644 45444 21646
rect 45276 20916 45332 21644
rect 45388 21634 45444 21644
rect 45724 21700 45780 21710
rect 44940 20860 45332 20916
rect 44940 20802 44996 20860
rect 44940 20750 44942 20802
rect 44994 20750 44996 20802
rect 44940 20738 44996 20750
rect 44156 20178 44212 20188
rect 45276 20188 45332 20860
rect 45500 21588 45556 21598
rect 45500 20802 45556 21532
rect 45500 20750 45502 20802
rect 45554 20750 45556 20802
rect 45500 20738 45556 20750
rect 45724 20468 45780 21644
rect 46396 20692 46452 20702
rect 46284 20636 46396 20692
rect 45948 20580 46004 20590
rect 45948 20486 46004 20524
rect 45724 20188 45780 20412
rect 45276 20132 45668 20188
rect 45724 20132 46116 20188
rect 43484 19742 43486 19794
rect 43538 19742 43540 19794
rect 43484 19730 43540 19742
rect 45612 19570 45668 20132
rect 45612 19518 45614 19570
rect 45666 19518 45668 19570
rect 44268 19460 44324 19470
rect 44268 19366 44324 19404
rect 43372 18510 43374 18562
rect 43426 18510 43428 18562
rect 42140 18498 42196 18508
rect 41692 15810 41748 15820
rect 42140 17554 42196 17566
rect 42140 17502 42142 17554
rect 42194 17502 42196 17554
rect 41580 15764 41636 15774
rect 41580 15652 41636 15708
rect 42028 15764 42084 15774
rect 42140 15764 42196 17502
rect 42028 15762 42196 15764
rect 42028 15710 42030 15762
rect 42082 15710 42196 15762
rect 42028 15708 42196 15710
rect 42028 15698 42084 15708
rect 41692 15652 41748 15662
rect 41580 15650 41748 15652
rect 41580 15598 41694 15650
rect 41746 15598 41748 15650
rect 41580 15596 41748 15598
rect 42252 15652 42308 18508
rect 43372 18498 43428 18510
rect 45612 18564 45668 19518
rect 45612 18498 45668 18508
rect 46060 19570 46116 20132
rect 46060 19518 46062 19570
rect 46114 19518 46116 19570
rect 43484 18452 43540 18462
rect 43484 17892 43540 18396
rect 43036 17890 43540 17892
rect 43036 17838 43486 17890
rect 43538 17838 43540 17890
rect 43036 17836 43540 17838
rect 42924 17780 42980 17790
rect 42924 16884 42980 17724
rect 42924 16818 42980 16828
rect 43036 16660 43092 17836
rect 43484 17826 43540 17836
rect 45276 18450 45332 18462
rect 45276 18398 45278 18450
rect 45330 18398 45332 18450
rect 43932 17668 43988 17678
rect 43092 16604 43316 16660
rect 43036 16566 43092 16604
rect 42364 15876 42420 15886
rect 42364 15782 42420 15820
rect 42924 15652 42980 15662
rect 42252 15650 42980 15652
rect 42252 15598 42926 15650
rect 42978 15598 42980 15650
rect 42252 15596 42980 15598
rect 41692 15428 41748 15596
rect 41692 15362 41748 15372
rect 42364 15428 42420 15438
rect 41468 15026 41524 15036
rect 40292 14700 40628 14756
rect 40236 14662 40292 14700
rect 40348 13858 40404 14700
rect 40572 14530 40628 14700
rect 40572 14478 40574 14530
rect 40626 14478 40628 14530
rect 40572 14466 40628 14478
rect 41692 14754 41748 14766
rect 42364 14756 42420 15372
rect 41692 14702 41694 14754
rect 41746 14702 41748 14754
rect 40348 13806 40350 13858
rect 40402 13806 40404 13858
rect 40348 13748 40404 13806
rect 41356 13860 41412 13870
rect 41356 13766 41412 13804
rect 41020 13748 41076 13758
rect 40404 13692 40628 13748
rect 40348 13682 40404 13692
rect 38108 12738 38164 12796
rect 38108 12686 38110 12738
rect 38162 12686 38164 12738
rect 38108 12674 38164 12686
rect 38556 12850 38612 12862
rect 38556 12798 38558 12850
rect 38610 12798 38612 12850
rect 38556 12738 38612 12798
rect 39116 12852 39172 12862
rect 39676 12852 39732 12862
rect 39116 12850 39396 12852
rect 39116 12798 39118 12850
rect 39170 12798 39396 12850
rect 39116 12796 39396 12798
rect 39116 12786 39172 12796
rect 38556 12686 38558 12738
rect 38610 12686 38612 12738
rect 38556 12674 38612 12686
rect 37324 12562 37380 12572
rect 38668 12628 38724 12638
rect 38668 10724 38724 12572
rect 39004 12628 39060 12638
rect 39004 12534 39060 12572
rect 39340 12628 39396 12796
rect 39340 12534 39396 12572
rect 39676 12626 39732 12796
rect 39676 12574 39678 12626
rect 39730 12574 39732 12626
rect 39676 12562 39732 12574
rect 39900 12626 39956 13468
rect 39900 12574 39902 12626
rect 39954 12574 39956 12626
rect 39900 12562 39956 12574
rect 40012 12628 40068 12638
rect 38780 11508 38836 11518
rect 38780 11506 38948 11508
rect 38780 11454 38782 11506
rect 38834 11454 38948 11506
rect 38780 11452 38948 11454
rect 38780 11442 38836 11452
rect 38780 10724 38836 10734
rect 38668 10722 38836 10724
rect 38668 10670 38782 10722
rect 38834 10670 38836 10722
rect 38668 10668 38836 10670
rect 37212 9314 37268 9324
rect 37324 10612 37380 10622
rect 37324 9604 37380 10556
rect 38332 10612 38388 10622
rect 38332 10518 38388 10556
rect 35644 8642 35700 8652
rect 36204 8708 36260 8718
rect 36204 8614 36260 8652
rect 37324 8596 37380 9548
rect 38780 9602 38836 10668
rect 38892 10388 38948 11452
rect 39228 11506 39284 11518
rect 39228 11454 39230 11506
rect 39282 11454 39284 11506
rect 39228 10612 39284 11454
rect 39228 10546 39284 10556
rect 39676 10612 39732 10622
rect 39676 10518 39732 10556
rect 39452 10500 39508 10510
rect 39340 10444 39452 10500
rect 39228 10388 39284 10398
rect 39340 10388 39396 10444
rect 39452 10434 39508 10444
rect 38892 10386 39396 10388
rect 38892 10334 39230 10386
rect 39282 10334 39396 10386
rect 38892 10332 39396 10334
rect 39228 10322 39284 10332
rect 38780 9550 38782 9602
rect 38834 9550 38836 9602
rect 37660 9492 37716 9502
rect 37324 8594 37604 8596
rect 37324 8542 37326 8594
rect 37378 8542 37604 8594
rect 37324 8540 37604 8542
rect 37324 8530 37380 8540
rect 35084 8430 35086 8482
rect 35138 8430 35140 8482
rect 35084 8428 35140 8430
rect 35084 8372 35364 8428
rect 35308 8148 35364 8372
rect 35308 8082 35364 8092
rect 36652 8148 36708 8158
rect 36652 7810 36708 8092
rect 36652 7758 36654 7810
rect 36706 7758 36708 7810
rect 36652 7746 36708 7758
rect 37100 7922 37156 7934
rect 37100 7870 37102 7922
rect 37154 7870 37156 7922
rect 37100 7810 37156 7870
rect 37100 7758 37102 7810
rect 37154 7758 37156 7810
rect 37100 7746 37156 7758
rect 37548 7810 37604 8540
rect 37660 8594 37716 9436
rect 37660 8542 37662 8594
rect 37714 8542 37716 8594
rect 37660 8372 37716 8542
rect 37660 7922 37716 8316
rect 38780 8484 38836 9550
rect 38780 8148 38836 8428
rect 40012 8708 40068 12572
rect 40572 12626 40628 13692
rect 41020 13654 41076 13692
rect 41692 13746 41748 14702
rect 41692 13694 41694 13746
rect 41746 13694 41748 13746
rect 41692 13682 41748 13694
rect 42028 14754 42420 14756
rect 42028 14702 42366 14754
rect 42418 14702 42420 14754
rect 42028 14700 42420 14702
rect 42028 13746 42084 14700
rect 42364 14690 42420 14700
rect 42700 15092 42756 15102
rect 42028 13694 42030 13746
rect 42082 13694 42084 13746
rect 42028 13682 42084 13694
rect 42364 13860 42420 13870
rect 42364 13746 42420 13804
rect 42700 13858 42756 15036
rect 42700 13806 42702 13858
rect 42754 13806 42756 13858
rect 42700 13794 42756 13806
rect 42364 13694 42366 13746
rect 42418 13694 42420 13746
rect 42364 13682 42420 13694
rect 42924 13412 42980 15596
rect 43148 13746 43204 13758
rect 43148 13694 43150 13746
rect 43202 13694 43204 13746
rect 43148 13412 43204 13694
rect 40572 12574 40574 12626
rect 40626 12574 40628 12626
rect 40572 12562 40628 12574
rect 42476 13356 43204 13412
rect 42140 12516 42196 12526
rect 40012 8482 40068 8652
rect 40012 8430 40014 8482
rect 40066 8430 40068 8482
rect 40012 8418 40068 8430
rect 40124 10610 40180 10622
rect 40124 10558 40126 10610
rect 40178 10558 40180 10610
rect 40124 10500 40180 10558
rect 40348 10612 40404 10622
rect 40404 10556 40516 10612
rect 40348 10546 40404 10556
rect 40124 8372 40180 10444
rect 40236 9604 40292 9614
rect 40236 9510 40292 9548
rect 40460 8708 40516 10556
rect 42140 10388 42196 12460
rect 42028 10386 42196 10388
rect 42028 10334 42142 10386
rect 42194 10334 42196 10386
rect 42028 10332 42196 10334
rect 42028 10052 42084 10332
rect 42140 10322 42196 10332
rect 41804 9996 42084 10052
rect 40908 9604 40964 9614
rect 40908 9510 40964 9548
rect 41244 9602 41300 9614
rect 41580 9604 41636 9614
rect 41244 9550 41246 9602
rect 41298 9550 41300 9602
rect 41244 9380 41300 9550
rect 41244 9314 41300 9324
rect 41356 9602 41636 9604
rect 41356 9550 41582 9602
rect 41634 9550 41636 9602
rect 41356 9548 41636 9550
rect 41356 9044 41412 9548
rect 41580 9538 41636 9548
rect 41132 8988 41412 9044
rect 41132 8818 41188 8988
rect 41132 8766 41134 8818
rect 41186 8766 41188 8818
rect 41132 8754 41188 8766
rect 40348 8596 40404 8606
rect 40236 8594 40404 8596
rect 40236 8542 40350 8594
rect 40402 8542 40404 8594
rect 40236 8540 40404 8542
rect 40236 8484 40292 8540
rect 40348 8530 40404 8540
rect 40460 8428 40516 8652
rect 40236 8418 40292 8428
rect 40124 8306 40180 8316
rect 40348 8372 40516 8428
rect 41020 8596 41076 8606
rect 38780 8082 38836 8092
rect 37660 7870 37662 7922
rect 37714 7870 37716 7922
rect 37660 7858 37716 7870
rect 37548 7758 37550 7810
rect 37602 7758 37604 7810
rect 37548 7746 37604 7758
rect 40348 7810 40404 8372
rect 40348 7758 40350 7810
rect 40402 7758 40404 7810
rect 40348 7746 40404 7758
rect 41020 7810 41076 8540
rect 41804 8594 41860 9996
rect 41916 9828 41972 9838
rect 41916 9734 41972 9772
rect 42476 9714 42532 13356
rect 43260 12852 43316 16604
rect 43372 16546 43428 16558
rect 43372 16494 43374 16546
rect 43426 16494 43428 16546
rect 43372 15204 43428 16494
rect 43932 16548 43988 17612
rect 45276 17668 45332 18398
rect 45724 18452 45780 18462
rect 45724 18358 45780 18396
rect 45276 17602 45332 17612
rect 45948 17668 46004 17678
rect 45948 17574 46004 17612
rect 43932 16482 43988 16492
rect 44716 17442 44772 17454
rect 44716 17390 44718 17442
rect 44770 17390 44772 17442
rect 44716 16436 44772 17390
rect 44828 16772 44884 16782
rect 44828 16546 44884 16716
rect 46060 16660 46116 19518
rect 46284 18452 46340 20636
rect 46396 20598 46452 20636
rect 46844 20468 46900 20478
rect 46732 20466 46900 20468
rect 46732 20414 46846 20466
rect 46898 20414 46900 20466
rect 46732 20412 46900 20414
rect 46284 18386 46340 18396
rect 46396 20244 46452 20254
rect 46396 18786 46452 20188
rect 46732 20132 46788 20412
rect 46844 20402 46900 20412
rect 46732 20066 46788 20076
rect 46396 18734 46398 18786
rect 46450 18734 46452 18786
rect 46284 16660 46340 16670
rect 46060 16658 46340 16660
rect 46060 16606 46286 16658
rect 46338 16606 46340 16658
rect 46060 16604 46340 16606
rect 46284 16594 46340 16604
rect 44828 16494 44830 16546
rect 44882 16494 44884 16546
rect 44828 16436 44884 16494
rect 46060 16436 46116 16446
rect 44828 16380 45108 16436
rect 44156 16322 44212 16334
rect 44156 16270 44158 16322
rect 44210 16270 44212 16322
rect 44156 15874 44212 16270
rect 44156 15822 44158 15874
rect 44210 15822 44212 15874
rect 44156 15810 44212 15822
rect 44716 15876 44772 16380
rect 44940 15876 44996 15886
rect 44716 15874 44996 15876
rect 44716 15822 44942 15874
rect 44994 15822 44996 15874
rect 44716 15820 44996 15822
rect 43484 15764 43540 15774
rect 43484 15670 43540 15708
rect 44940 15764 44996 15820
rect 44940 15698 44996 15708
rect 43372 15148 43540 15204
rect 43260 12786 43316 12796
rect 43484 14532 43540 15148
rect 43820 14756 43876 14766
rect 43820 14662 43876 14700
rect 42924 12516 42980 12526
rect 42924 12422 42980 12460
rect 43484 12516 43540 14476
rect 44940 14532 44996 14542
rect 45052 14532 45108 16380
rect 46060 16342 46116 16380
rect 46172 15764 46228 15774
rect 46396 15764 46452 18734
rect 46620 19906 46676 19918
rect 46620 19854 46622 19906
rect 46674 19854 46676 19906
rect 46620 17892 46676 19854
rect 46956 19796 47012 19806
rect 46620 17826 46676 17836
rect 46732 18452 46788 18462
rect 46732 17780 46788 18396
rect 46844 17780 46900 17790
rect 46732 17778 46900 17780
rect 46732 17726 46846 17778
rect 46898 17726 46900 17778
rect 46732 17724 46900 17726
rect 46732 16658 46788 17724
rect 46844 17714 46900 17724
rect 46956 17668 47012 19740
rect 47068 18564 47124 18574
rect 47068 18470 47124 18508
rect 47404 18004 47460 24556
rect 47852 24546 47908 24556
rect 47964 24610 48356 24612
rect 47964 24558 48302 24610
rect 48354 24558 48356 24610
rect 47964 24556 48356 24558
rect 47740 24052 47796 24062
rect 47516 23940 47572 23950
rect 47516 23846 47572 23884
rect 47740 23826 47796 23996
rect 47740 23774 47742 23826
rect 47794 23774 47796 23826
rect 47740 23762 47796 23774
rect 47964 23492 48020 24556
rect 48300 24546 48356 24556
rect 47628 23436 48020 23492
rect 48188 24388 48244 24398
rect 47628 22706 47684 23436
rect 47628 22654 47630 22706
rect 47682 22654 47684 22706
rect 47628 22642 47684 22654
rect 48188 22706 48244 24332
rect 48188 22654 48190 22706
rect 48242 22654 48244 22706
rect 48188 22642 48244 22654
rect 48524 21700 48580 26348
rect 49196 25058 49252 29708
rect 49308 29762 49364 29774
rect 49308 29710 49310 29762
rect 49362 29710 49364 29762
rect 49308 29652 49364 29710
rect 49308 29586 49364 29596
rect 49420 27858 49476 31836
rect 50204 31892 50260 33742
rect 50316 33572 50372 34638
rect 50428 34132 50484 35868
rect 50876 35810 50932 35822
rect 50876 35758 50878 35810
rect 50930 35758 50932 35810
rect 50876 34692 50932 35758
rect 50876 34626 50932 34636
rect 51100 34804 51156 36652
rect 51212 36706 51380 36708
rect 51212 36654 51214 36706
rect 51266 36654 51380 36706
rect 51212 36652 51380 36654
rect 51212 36642 51268 36652
rect 51548 36034 51604 36878
rect 51660 36594 51716 38110
rect 52556 37938 52612 38446
rect 52556 37886 52558 37938
rect 52610 37886 52612 37938
rect 52556 37874 52612 37886
rect 52780 37838 52836 38894
rect 53228 38610 53284 39900
rect 53452 39848 53508 39860
rect 53452 39796 53454 39848
rect 53506 39844 53508 39848
rect 53564 39844 53620 39854
rect 53506 39796 53564 39844
rect 53452 39788 53564 39796
rect 53452 39784 53508 39788
rect 53564 39778 53620 39788
rect 54012 39844 54068 39854
rect 54012 39750 54068 39788
rect 54348 39844 54404 39854
rect 54460 39844 54516 40798
rect 54572 40738 54628 41020
rect 54572 40686 54574 40738
rect 54626 40686 54628 40738
rect 54572 39956 54628 40686
rect 54572 39862 54628 39900
rect 54684 40404 54740 40414
rect 54348 39842 54516 39844
rect 54348 39790 54350 39842
rect 54402 39790 54516 39842
rect 54348 39788 54516 39790
rect 54348 39732 54404 39788
rect 54348 39666 54404 39676
rect 54684 38946 54740 40348
rect 54908 40066 54964 41806
rect 55580 40404 55636 41918
rect 55580 40338 55636 40348
rect 56140 40738 56196 40750
rect 56140 40686 56142 40738
rect 56194 40686 56196 40738
rect 54908 40014 54910 40066
rect 54962 40014 54964 40066
rect 54908 40002 54964 40014
rect 55580 39956 55636 39966
rect 55580 39954 56084 39956
rect 55580 39902 55582 39954
rect 55634 39902 56084 39954
rect 55580 39900 56084 39902
rect 55580 39890 55636 39900
rect 54684 38894 54686 38946
rect 54738 38894 54740 38946
rect 54684 38882 54740 38894
rect 55356 39844 55412 39854
rect 53228 38558 53230 38610
rect 53282 38558 53284 38610
rect 53228 38498 53284 38558
rect 53228 38446 53230 38498
rect 53282 38446 53284 38498
rect 53228 38434 53284 38446
rect 53676 38836 53732 38846
rect 53676 38610 53732 38780
rect 53676 38558 53678 38610
rect 53730 38558 53732 38610
rect 53676 38498 53732 38558
rect 53676 38446 53678 38498
rect 53730 38446 53732 38498
rect 53676 38434 53732 38446
rect 55356 38834 55412 39788
rect 55356 38782 55358 38834
rect 55410 38782 55412 38834
rect 52724 37826 52836 37838
rect 52724 37774 52726 37826
rect 52778 37774 52836 37826
rect 52724 37772 52836 37774
rect 53788 37826 53844 37838
rect 53788 37774 53790 37826
rect 53842 37774 53844 37826
rect 52724 37762 52780 37772
rect 53676 37492 53732 37502
rect 51996 36820 52052 36830
rect 51660 36542 51662 36594
rect 51714 36542 51716 36594
rect 51660 36484 51716 36542
rect 51660 36418 51716 36428
rect 51884 36596 51940 36606
rect 51548 35982 51550 36034
rect 51602 35982 51604 36034
rect 51548 35970 51604 35982
rect 50764 34580 50820 34590
rect 50764 34486 50820 34524
rect 50876 34468 50932 34478
rect 50876 34374 50932 34412
rect 50556 34300 50820 34310
rect 50612 34244 50660 34300
rect 50716 34244 50764 34300
rect 50556 34234 50820 34244
rect 50540 34132 50596 34142
rect 50428 34130 50596 34132
rect 50428 34078 50542 34130
rect 50594 34078 50596 34130
rect 50428 34076 50596 34078
rect 50540 34066 50596 34076
rect 50316 33506 50372 33516
rect 51100 33794 51156 34748
rect 51548 34916 51604 34926
rect 51548 34802 51604 34860
rect 51548 34750 51550 34802
rect 51602 34750 51604 34802
rect 51548 34738 51604 34750
rect 51324 34692 51380 34702
rect 51324 34598 51380 34636
rect 51884 34690 51940 36540
rect 51996 36036 52052 36764
rect 53676 36818 53732 37436
rect 53676 36766 53678 36818
rect 53730 36766 53732 36818
rect 53676 36754 53732 36766
rect 53788 37044 53844 37774
rect 54348 37492 54404 37502
rect 54348 37398 54404 37436
rect 52108 36708 52164 36718
rect 53004 36708 53060 36718
rect 53340 36708 53396 36718
rect 52108 36706 53060 36708
rect 52108 36654 52110 36706
rect 52162 36654 53006 36706
rect 53058 36654 53060 36706
rect 52108 36652 53060 36654
rect 52108 36642 52164 36652
rect 53004 36642 53060 36652
rect 53116 36706 53396 36708
rect 53116 36654 53342 36706
rect 53394 36654 53396 36706
rect 53116 36652 53396 36654
rect 53116 36260 53172 36652
rect 53340 36642 53396 36652
rect 52556 36204 53172 36260
rect 53452 36484 53508 36494
rect 52332 36036 52388 36046
rect 51996 35980 52332 36036
rect 52332 35942 52388 35980
rect 51884 34638 51886 34690
rect 51938 34638 51940 34690
rect 51884 34626 51940 34638
rect 52556 33908 52612 36204
rect 52780 36036 52836 36046
rect 52780 34802 52836 35980
rect 53452 36036 53508 36428
rect 53788 36372 53844 36988
rect 55356 37044 55412 38782
rect 56028 38052 56084 39900
rect 56140 39844 56196 40686
rect 56140 39778 56196 39788
rect 56476 39732 56532 39742
rect 56476 38834 56532 39676
rect 56476 38782 56478 38834
rect 56530 38782 56532 38834
rect 56476 38770 56532 38782
rect 56700 39730 56756 39742
rect 56700 39678 56702 39730
rect 56754 39678 56756 39730
rect 56700 38612 56756 39678
rect 57148 39732 57204 39742
rect 57148 39638 57204 39676
rect 56700 38546 56756 38556
rect 57036 38612 57092 38622
rect 55356 36978 55412 36988
rect 55468 38050 56084 38052
rect 55468 37998 56030 38050
rect 56082 37998 56084 38050
rect 55468 37996 56084 37998
rect 54460 36932 54516 36942
rect 54460 36706 54516 36876
rect 54460 36654 54462 36706
rect 54514 36654 54516 36706
rect 54460 36642 54516 36654
rect 55132 36708 55188 36718
rect 55356 36708 55412 36718
rect 55468 36708 55524 37996
rect 56028 37986 56084 37996
rect 55132 36614 55188 36652
rect 55244 36652 55356 36708
rect 55412 36652 55524 36708
rect 55580 37716 55636 37726
rect 54012 36596 54068 36606
rect 54012 36502 54068 36540
rect 55244 36484 55300 36652
rect 55356 36614 55412 36652
rect 55244 36418 55300 36428
rect 53788 36316 54068 36372
rect 53452 35980 53956 36036
rect 53452 35810 53508 35980
rect 53452 35758 53454 35810
rect 53506 35758 53508 35810
rect 53452 35746 53508 35758
rect 53676 35812 53732 35822
rect 53564 35586 53620 35598
rect 53564 35534 53566 35586
rect 53618 35534 53620 35586
rect 53452 35364 53508 35374
rect 52780 34750 52782 34802
rect 52834 34750 52836 34802
rect 52780 34738 52836 34750
rect 53004 34804 53060 34814
rect 53004 34710 53060 34748
rect 53452 34804 53508 35308
rect 53452 34710 53508 34748
rect 53228 34692 53284 34702
rect 52892 34578 52948 34590
rect 52892 34526 52894 34578
rect 52946 34526 52948 34578
rect 52556 33906 52836 33908
rect 52556 33854 52558 33906
rect 52610 33854 52836 33906
rect 52556 33852 52836 33854
rect 52556 33842 52612 33852
rect 51100 33742 51102 33794
rect 51154 33742 51156 33794
rect 50652 33010 50708 33022
rect 50652 32958 50654 33010
rect 50706 32958 50708 33010
rect 50652 32900 50708 32958
rect 50428 32898 50708 32900
rect 50428 32846 50654 32898
rect 50706 32846 50708 32898
rect 50428 32844 50708 32846
rect 50428 31948 50484 32844
rect 50652 32834 50708 32844
rect 51100 32898 51156 33742
rect 51324 33794 51380 33806
rect 51324 33742 51326 33794
rect 51378 33742 51380 33794
rect 51212 33012 51268 33022
rect 51324 33012 51380 33742
rect 51772 33796 51828 33806
rect 52220 33796 52276 33806
rect 51772 33794 52276 33796
rect 51772 33742 51774 33794
rect 51826 33742 52222 33794
rect 52274 33742 52276 33794
rect 51772 33740 52276 33742
rect 51772 33730 51828 33740
rect 52220 33730 52276 33740
rect 51212 33010 51380 33012
rect 51212 32958 51214 33010
rect 51266 32958 51380 33010
rect 51212 32956 51380 32958
rect 52780 33684 52836 33852
rect 52892 33906 52948 34526
rect 53228 34018 53284 34636
rect 53228 33966 53230 34018
rect 53282 33966 53284 34018
rect 53228 33954 53284 33966
rect 52892 33854 52894 33906
rect 52946 33854 52948 33906
rect 52892 33842 52948 33854
rect 52780 33628 53284 33684
rect 51212 32946 51268 32956
rect 51100 32846 51102 32898
rect 51154 32846 51156 32898
rect 51100 32788 51156 32846
rect 51100 32732 51604 32788
rect 50556 32284 50820 32294
rect 50612 32228 50660 32284
rect 50716 32228 50764 32284
rect 50556 32218 50820 32228
rect 50204 31826 50260 31836
rect 50316 31892 50484 31948
rect 51548 32002 51604 32732
rect 51548 31950 51550 32002
rect 51602 31950 51604 32002
rect 49868 31778 49924 31790
rect 49868 31726 49870 31778
rect 49922 31726 49924 31778
rect 49532 31668 49588 31678
rect 49868 31668 49924 31726
rect 49532 31666 49924 31668
rect 49532 31614 49534 31666
rect 49586 31614 49924 31666
rect 49532 31612 49924 31614
rect 50204 31668 50260 31678
rect 49532 31556 49588 31612
rect 50204 31574 50260 31612
rect 49532 31490 49588 31500
rect 50316 30772 50372 31892
rect 50316 30706 50372 30716
rect 51100 31666 51156 31678
rect 51100 31614 51102 31666
rect 51154 31614 51156 31666
rect 49980 30548 50036 30558
rect 50036 30492 50372 30548
rect 49980 30454 50036 30492
rect 50316 30436 50372 30492
rect 50316 30380 50484 30436
rect 49644 29876 49700 29886
rect 49644 29782 49700 29820
rect 49868 29764 49924 29774
rect 49420 27806 49422 27858
rect 49474 27806 49476 27858
rect 49420 27074 49476 27806
rect 49420 27022 49422 27074
rect 49474 27022 49476 27074
rect 49420 27010 49476 27022
rect 49756 28868 49812 28878
rect 49756 28082 49812 28812
rect 49868 28866 49924 29708
rect 49868 28814 49870 28866
rect 49922 28814 49924 28866
rect 49868 28802 49924 28814
rect 49756 28030 49758 28082
rect 49810 28030 49812 28082
rect 49756 26908 49812 28030
rect 50316 28756 50372 28766
rect 50316 27748 50372 28700
rect 50428 28532 50484 30380
rect 50988 30324 51044 30334
rect 50556 30268 50820 30278
rect 50612 30212 50660 30268
rect 50716 30212 50764 30268
rect 50556 30202 50820 30212
rect 50540 30098 50596 30110
rect 50540 30046 50542 30098
rect 50594 30046 50596 30098
rect 50540 29650 50596 30046
rect 50540 29598 50542 29650
rect 50594 29598 50596 29650
rect 50540 28756 50596 29598
rect 50876 29876 50932 29886
rect 50876 29090 50932 29820
rect 50876 29038 50878 29090
rect 50930 29038 50932 29090
rect 50876 29026 50932 29038
rect 50988 29650 51044 30268
rect 51100 30098 51156 31614
rect 51548 31556 51604 31950
rect 52108 32562 52164 32574
rect 52108 32510 52110 32562
rect 52162 32510 52164 32562
rect 51996 31892 52052 31902
rect 52108 31892 52164 32510
rect 51996 31890 52108 31892
rect 51996 31838 51998 31890
rect 52050 31838 52108 31890
rect 51996 31836 52108 31838
rect 51996 31826 52052 31836
rect 52108 31826 52164 31836
rect 52444 31780 52500 31790
rect 51548 31490 51604 31500
rect 51660 31668 51716 31678
rect 51100 30046 51102 30098
rect 51154 30046 51156 30098
rect 51100 30034 51156 30046
rect 51324 30436 51380 30446
rect 51324 29874 51380 30380
rect 51324 29822 51326 29874
rect 51378 29822 51380 29874
rect 51324 29810 51380 29822
rect 51660 29874 51716 31612
rect 52444 31666 52500 31724
rect 52444 31614 52446 31666
rect 52498 31614 52500 31666
rect 51884 30436 51940 30446
rect 51884 30434 52052 30436
rect 51884 30382 51886 30434
rect 51938 30382 52052 30434
rect 51884 30380 52052 30382
rect 51884 30370 51940 30380
rect 51660 29822 51662 29874
rect 51714 29822 51716 29874
rect 51660 29810 51716 29822
rect 51996 29874 52052 30380
rect 52444 30324 52500 31614
rect 52780 31668 52836 33628
rect 53228 32786 53284 33628
rect 53228 32734 53230 32786
rect 53282 32734 53284 32786
rect 53228 32722 53284 32734
rect 53564 32786 53620 35534
rect 53564 32734 53566 32786
rect 53618 32734 53620 32786
rect 53564 32722 53620 32734
rect 53676 32788 53732 35756
rect 53900 34914 53956 35980
rect 54012 35810 54068 36316
rect 54236 36036 54292 36046
rect 54236 35922 54292 35980
rect 54236 35870 54238 35922
rect 54290 35870 54292 35922
rect 54236 35858 54292 35870
rect 54012 35758 54014 35810
rect 54066 35758 54068 35810
rect 54012 35746 54068 35758
rect 54572 35812 54628 35822
rect 54572 35718 54628 35756
rect 55580 35812 55636 37660
rect 56700 37714 56756 37726
rect 56700 37662 56702 37714
rect 56754 37662 56756 37714
rect 56700 37044 56756 37662
rect 57036 37716 57092 38556
rect 57036 37650 57092 37660
rect 57148 37714 57204 37726
rect 57148 37662 57150 37714
rect 57202 37662 57204 37714
rect 57148 37044 57204 37662
rect 57596 37716 57652 37726
rect 57596 37622 57652 37660
rect 56700 36988 57092 37044
rect 56924 36818 56980 36830
rect 56924 36766 56926 36818
rect 56978 36766 56980 36818
rect 56700 36708 56756 36718
rect 55580 35746 55636 35756
rect 55804 36594 55860 36606
rect 55804 36542 55806 36594
rect 55858 36542 55860 36594
rect 53900 34862 53902 34914
rect 53954 34862 53956 34914
rect 53900 34850 53956 34862
rect 55020 35476 55076 35486
rect 54348 34020 54404 34030
rect 54348 33906 54404 33964
rect 55020 34018 55076 35420
rect 55580 35476 55636 35486
rect 55580 35382 55636 35420
rect 55468 35140 55524 35150
rect 55804 35140 55860 36542
rect 56588 36596 56644 36606
rect 56588 36502 56644 36540
rect 56700 36034 56756 36652
rect 56700 35982 56702 36034
rect 56754 35982 56756 36034
rect 55468 35138 55860 35140
rect 55468 35086 55470 35138
rect 55522 35086 55860 35138
rect 55468 35084 55860 35086
rect 55916 35810 55972 35822
rect 55916 35758 55918 35810
rect 55970 35758 55972 35810
rect 55916 35364 55972 35758
rect 56700 35474 56756 35982
rect 56924 35812 56980 36766
rect 57036 36708 57092 36988
rect 57148 36978 57204 36988
rect 57484 37044 57540 37054
rect 57484 36820 57540 36988
rect 57484 36818 57764 36820
rect 57484 36766 57486 36818
rect 57538 36766 57764 36818
rect 57484 36764 57764 36766
rect 57484 36754 57540 36764
rect 57148 36708 57204 36718
rect 57036 36706 57204 36708
rect 57036 36654 57150 36706
rect 57202 36654 57204 36706
rect 57036 36652 57204 36654
rect 56924 35746 56980 35756
rect 56700 35422 56702 35474
rect 56754 35422 56756 35474
rect 56700 35410 56756 35422
rect 57148 35700 57204 36652
rect 57596 35700 57652 35710
rect 57148 35698 57652 35700
rect 57148 35646 57150 35698
rect 57202 35646 57598 35698
rect 57650 35646 57652 35698
rect 57148 35644 57652 35646
rect 57148 35364 57204 35644
rect 57596 35634 57652 35644
rect 55468 35074 55524 35084
rect 55020 33966 55022 34018
rect 55074 33966 55076 34018
rect 55020 33954 55076 33966
rect 55468 34802 55524 34814
rect 55468 34750 55470 34802
rect 55522 34750 55524 34802
rect 54348 33854 54350 33906
rect 54402 33854 54404 33906
rect 54348 33842 54404 33854
rect 53788 33796 53844 33806
rect 55468 33796 55524 34750
rect 55804 34692 55860 34702
rect 55916 34692 55972 35308
rect 55804 34690 55972 34692
rect 55804 34638 55806 34690
rect 55858 34638 55972 34690
rect 55804 34636 55972 34638
rect 55804 34626 55860 34636
rect 55804 34020 55860 34030
rect 55804 33926 55860 33964
rect 55580 33796 55636 33806
rect 53788 33794 54292 33796
rect 53788 33742 53790 33794
rect 53842 33742 54292 33794
rect 53788 33740 54292 33742
rect 55468 33740 55580 33796
rect 55916 33796 55972 34636
rect 56812 35308 57204 35364
rect 57372 35474 57428 35486
rect 57372 35422 57374 35474
rect 57426 35422 57428 35474
rect 56028 33796 56084 33806
rect 55916 33794 56084 33796
rect 55916 33742 56030 33794
rect 56082 33742 56084 33794
rect 55916 33740 56084 33742
rect 53788 33730 53844 33740
rect 53676 32722 53732 32732
rect 53900 33572 53956 33582
rect 53900 32786 53956 33516
rect 53900 32734 53902 32786
rect 53954 32734 53956 32786
rect 53900 32722 53956 32734
rect 52892 32674 52948 32686
rect 52892 32622 52894 32674
rect 52946 32622 52948 32674
rect 52892 32002 52948 32622
rect 54236 32676 54292 33740
rect 55580 33730 55636 33740
rect 55692 33684 55748 33694
rect 55132 32788 55188 32798
rect 54348 32676 54404 32686
rect 54236 32674 54404 32676
rect 54236 32622 54350 32674
rect 54402 32622 54404 32674
rect 54236 32620 54404 32622
rect 52892 31950 52894 32002
rect 52946 31950 52948 32002
rect 52892 31938 52948 31950
rect 52780 31602 52836 31612
rect 53340 31890 53396 31902
rect 53340 31838 53342 31890
rect 53394 31838 53396 31890
rect 53340 31556 53396 31838
rect 53676 31892 53732 31902
rect 53452 31780 53508 31790
rect 53452 31686 53508 31724
rect 53004 30658 53060 30670
rect 53004 30606 53006 30658
rect 53058 30606 53060 30658
rect 52556 30436 52612 30446
rect 52556 30342 52612 30380
rect 52444 30258 52500 30268
rect 53004 30324 53060 30606
rect 53340 30660 53396 31500
rect 53676 30882 53732 31836
rect 53676 30830 53678 30882
rect 53730 30830 53732 30882
rect 53676 30818 53732 30830
rect 53564 30660 53620 30670
rect 53340 30604 53564 30660
rect 53564 30566 53620 30604
rect 54236 30660 54292 30670
rect 54236 30566 54292 30604
rect 53004 30258 53060 30268
rect 54236 30324 54292 30334
rect 51996 29822 51998 29874
rect 52050 29822 52052 29874
rect 51996 29810 52052 29822
rect 52780 29876 52836 29886
rect 52332 29764 52388 29774
rect 50988 29598 50990 29650
rect 51042 29598 51044 29650
rect 50540 28690 50596 28700
rect 50988 28644 51044 29598
rect 52108 29762 52388 29764
rect 52108 29710 52334 29762
rect 52386 29710 52388 29762
rect 52108 29708 52388 29710
rect 52108 29204 52164 29708
rect 52332 29698 52388 29708
rect 51884 29148 52164 29204
rect 51548 28756 51604 28766
rect 51436 28754 51604 28756
rect 51436 28702 51550 28754
rect 51602 28702 51604 28754
rect 51436 28700 51604 28702
rect 50988 28578 51044 28588
rect 51324 28642 51380 28654
rect 51324 28590 51326 28642
rect 51378 28590 51380 28642
rect 50652 28532 50708 28542
rect 50428 28530 50708 28532
rect 50428 28478 50654 28530
rect 50706 28478 50708 28530
rect 50428 28476 50708 28478
rect 50652 28420 50708 28476
rect 50652 28364 50932 28420
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 49644 26852 49812 26908
rect 49980 27746 50372 27748
rect 49980 27694 50318 27746
rect 50370 27694 50372 27746
rect 49980 27692 50372 27694
rect 49308 26516 49364 26526
rect 49308 26422 49364 26460
rect 49308 25956 49364 25966
rect 49308 25862 49364 25900
rect 49196 25006 49198 25058
rect 49250 25006 49252 25058
rect 49196 24994 49252 25006
rect 49084 24498 49140 24510
rect 49084 24446 49086 24498
rect 49138 24446 49140 24498
rect 49084 24386 49140 24446
rect 49084 24334 49086 24386
rect 49138 24334 49140 24386
rect 48748 24052 48804 24062
rect 48636 23940 48692 23950
rect 48636 23602 48692 23884
rect 48748 23826 48804 23996
rect 48748 23774 48750 23826
rect 48802 23774 48804 23826
rect 48748 23762 48804 23774
rect 48972 23828 49028 23838
rect 49084 23828 49140 24334
rect 49532 24498 49588 24510
rect 49532 24446 49534 24498
rect 49586 24446 49588 24498
rect 49532 23940 49588 24446
rect 49644 24388 49700 26852
rect 49756 26516 49812 26526
rect 49980 26516 50036 27692
rect 50316 27682 50372 27692
rect 50540 27746 50596 27758
rect 50540 27694 50542 27746
rect 50594 27694 50596 27746
rect 50092 27074 50148 27086
rect 50092 27022 50094 27074
rect 50146 27022 50148 27074
rect 50092 26738 50148 27022
rect 50092 26686 50094 26738
rect 50146 26686 50148 26738
rect 50092 26674 50148 26686
rect 50428 26964 50484 26974
rect 49756 26514 50036 26516
rect 49756 26462 49758 26514
rect 49810 26462 50036 26514
rect 49756 26460 50036 26462
rect 50204 26516 50260 26526
rect 49756 26450 49812 26460
rect 49756 26066 49812 26078
rect 49756 26014 49758 26066
rect 49810 26014 49812 26066
rect 49756 25954 49812 26014
rect 49756 25902 49758 25954
rect 49810 25902 49812 25954
rect 49756 25890 49812 25902
rect 49644 24322 49700 24332
rect 49868 25506 49924 26460
rect 50204 25620 50260 26460
rect 50428 26402 50484 26908
rect 50540 26516 50596 27694
rect 50876 27748 50932 28364
rect 51324 27972 51380 28590
rect 51324 27906 51380 27916
rect 51212 27748 51268 27758
rect 50876 27746 51268 27748
rect 50876 27694 51214 27746
rect 51266 27694 51268 27746
rect 50876 27692 51268 27694
rect 51212 27300 51268 27692
rect 51324 27524 51380 27534
rect 51436 27524 51492 28700
rect 51548 28690 51604 28700
rect 51884 28642 51940 29148
rect 52780 28868 52836 29820
rect 54124 29874 54180 29886
rect 54124 29822 54126 29874
rect 54178 29822 54180 29874
rect 53452 29764 53508 29774
rect 53452 29670 53508 29708
rect 54012 29092 54068 29102
rect 54124 29092 54180 29822
rect 54012 29090 54180 29092
rect 54012 29038 54014 29090
rect 54066 29038 54180 29090
rect 54012 29036 54180 29038
rect 54012 29026 54068 29036
rect 52780 28802 52836 28812
rect 54012 28868 54068 28878
rect 52780 28644 52836 28654
rect 51884 28590 51886 28642
rect 51938 28590 51940 28642
rect 51884 28578 51940 28590
rect 52668 28588 52780 28644
rect 51548 27972 51604 27982
rect 51548 27970 52164 27972
rect 51548 27918 51550 27970
rect 51602 27918 52164 27970
rect 51548 27916 52164 27918
rect 51548 27906 51604 27916
rect 52108 27858 52164 27916
rect 52108 27806 52110 27858
rect 52162 27806 52164 27858
rect 52108 27794 52164 27806
rect 51380 27468 51492 27524
rect 51548 27746 51604 27758
rect 51548 27694 51550 27746
rect 51602 27694 51604 27746
rect 51324 27458 51380 27468
rect 51212 27244 51492 27300
rect 50764 26740 50820 26750
rect 50764 26738 50932 26740
rect 50764 26686 50766 26738
rect 50818 26686 50932 26738
rect 50764 26684 50932 26686
rect 50764 26674 50820 26684
rect 50540 26450 50596 26460
rect 50428 26350 50430 26402
rect 50482 26350 50484 26402
rect 50204 25618 50372 25620
rect 50204 25566 50206 25618
rect 50258 25566 50372 25618
rect 50204 25564 50372 25566
rect 50204 25554 50260 25564
rect 49868 25454 49870 25506
rect 49922 25454 49924 25506
rect 49868 24052 49924 25454
rect 50092 25060 50148 25070
rect 50092 25058 50260 25060
rect 50092 25006 50094 25058
rect 50146 25006 50260 25058
rect 50092 25004 50260 25006
rect 50092 24994 50148 25004
rect 50204 24946 50260 25004
rect 50204 24894 50206 24946
rect 50258 24894 50260 24946
rect 50204 24882 50260 24894
rect 49980 24498 50036 24510
rect 49980 24446 49982 24498
rect 50034 24446 50036 24498
rect 49980 24386 50036 24446
rect 49980 24334 49982 24386
rect 50034 24334 50036 24386
rect 49980 24322 50036 24334
rect 49980 24052 50036 24062
rect 49868 23996 49980 24052
rect 49588 23884 49700 23940
rect 49532 23874 49588 23884
rect 49028 23772 49140 23828
rect 48636 23550 48638 23602
rect 48690 23550 48692 23602
rect 48636 23538 48692 23550
rect 48972 23602 49028 23772
rect 48972 23550 48974 23602
rect 49026 23550 49028 23602
rect 48972 23538 49028 23550
rect 49644 23604 49700 23884
rect 49980 23938 50036 23996
rect 49980 23886 49982 23938
rect 50034 23886 50036 23938
rect 49980 23874 50036 23886
rect 49644 23538 49700 23548
rect 50204 23716 50260 23726
rect 50316 23716 50372 25564
rect 50428 25394 50484 26350
rect 50556 26236 50820 26246
rect 50612 26180 50660 26236
rect 50716 26180 50764 26236
rect 50556 26170 50820 26180
rect 50764 25956 50820 25966
rect 50876 25956 50932 26684
rect 50988 26738 51044 26750
rect 50988 26686 50990 26738
rect 51042 26686 51044 26738
rect 50988 26066 51044 26686
rect 51212 26738 51268 26750
rect 51212 26686 51214 26738
rect 51266 26686 51268 26738
rect 51100 26516 51156 26526
rect 51212 26516 51268 26686
rect 51156 26460 51268 26516
rect 51436 26740 51492 27244
rect 51548 26740 51604 27694
rect 51996 27748 52052 27758
rect 51660 26740 51716 26750
rect 51548 26738 51716 26740
rect 51548 26686 51662 26738
rect 51714 26686 51716 26738
rect 51548 26684 51716 26686
rect 51436 26626 51492 26684
rect 51436 26574 51438 26626
rect 51490 26574 51492 26626
rect 51100 26450 51156 26460
rect 50988 26014 50990 26066
rect 51042 26014 51044 26066
rect 50988 26002 51044 26014
rect 50820 25900 50932 25956
rect 51436 25956 51492 26574
rect 51548 25956 51604 25966
rect 51436 25954 51604 25956
rect 51436 25902 51550 25954
rect 51602 25902 51604 25954
rect 51436 25900 51604 25902
rect 50764 25890 50820 25900
rect 50876 25732 50932 25742
rect 50652 25618 50708 25630
rect 50652 25566 50654 25618
rect 50706 25566 50708 25618
rect 50652 25506 50708 25566
rect 50652 25454 50654 25506
rect 50706 25454 50708 25506
rect 50652 25442 50708 25454
rect 50428 25342 50430 25394
rect 50482 25342 50484 25394
rect 50428 25330 50484 25342
rect 50652 24612 50708 24622
rect 50428 24610 50708 24612
rect 50428 24558 50654 24610
rect 50706 24558 50708 24610
rect 50428 24556 50708 24558
rect 50428 23828 50484 24556
rect 50652 24546 50708 24556
rect 50556 24220 50820 24230
rect 50612 24164 50660 24220
rect 50716 24164 50764 24220
rect 50556 24154 50820 24164
rect 50652 24050 50708 24062
rect 50652 23998 50654 24050
rect 50706 23998 50708 24050
rect 50428 23772 50596 23828
rect 50260 23660 50372 23716
rect 49532 23490 49588 23502
rect 49532 23438 49534 23490
rect 49586 23438 49588 23490
rect 48524 21634 48580 21644
rect 48748 22594 48804 22606
rect 48748 22542 48750 22594
rect 48802 22542 48804 22594
rect 47852 21586 47908 21598
rect 47852 21534 47854 21586
rect 47906 21534 47908 21586
rect 47628 20580 47684 20590
rect 47516 20244 47572 20254
rect 47516 18676 47572 20188
rect 47628 19796 47684 20524
rect 47628 19730 47684 19740
rect 47740 20468 47796 20478
rect 47852 20468 47908 21534
rect 48076 20692 48132 20702
rect 48076 20598 48132 20636
rect 48636 20690 48692 20702
rect 48636 20638 48638 20690
rect 48690 20638 48692 20690
rect 47796 20412 47908 20468
rect 47740 19684 47796 20412
rect 48636 20356 48692 20638
rect 48636 20290 48692 20300
rect 48748 20188 48804 22542
rect 49420 22484 49476 22494
rect 49196 22482 49476 22484
rect 49196 22430 49422 22482
rect 49474 22430 49476 22482
rect 49196 22428 49476 22430
rect 49084 21812 49140 21822
rect 48860 21700 48916 21710
rect 48860 21606 48916 21644
rect 49084 20802 49140 21756
rect 49196 21026 49252 22428
rect 49420 22418 49476 22428
rect 49420 21812 49476 21822
rect 49532 21812 49588 23438
rect 49420 21810 49588 21812
rect 49420 21758 49422 21810
rect 49474 21758 49588 21810
rect 49420 21756 49588 21758
rect 50204 22482 50260 23660
rect 50428 23604 50484 23614
rect 50428 23510 50484 23548
rect 50540 23156 50596 23772
rect 50204 22430 50206 22482
rect 50258 22430 50260 22482
rect 49420 21746 49476 21756
rect 49756 21698 49812 21710
rect 49756 21646 49758 21698
rect 49810 21646 49812 21698
rect 49756 21476 49812 21646
rect 50092 21698 50148 21710
rect 50092 21646 50094 21698
rect 50146 21646 50148 21698
rect 49812 21420 49924 21476
rect 49756 21410 49812 21420
rect 49196 20974 49198 21026
rect 49250 20974 49252 21026
rect 49196 20962 49252 20974
rect 49084 20750 49086 20802
rect 49138 20750 49140 20802
rect 49084 20738 49140 20750
rect 49532 20690 49588 20702
rect 49532 20638 49534 20690
rect 49586 20638 49588 20690
rect 49532 20468 49588 20638
rect 49532 20188 49588 20412
rect 48300 20132 48804 20188
rect 49084 20132 49588 20188
rect 49756 20690 49812 20702
rect 49756 20638 49758 20690
rect 49810 20638 49812 20690
rect 48300 19906 48356 20132
rect 48300 19854 48302 19906
rect 48354 19854 48356 19906
rect 48300 19842 48356 19854
rect 49084 19794 49140 20132
rect 49084 19742 49086 19794
rect 49138 19742 49140 19794
rect 47740 19682 47908 19684
rect 47740 19630 47742 19682
rect 47794 19630 47908 19682
rect 47740 19628 47908 19630
rect 47740 19618 47796 19628
rect 47628 19570 47684 19582
rect 47628 19518 47630 19570
rect 47682 19518 47684 19570
rect 47628 18788 47684 19518
rect 47628 18732 47796 18788
rect 47516 18620 47684 18676
rect 47516 18450 47572 18462
rect 47516 18398 47518 18450
rect 47570 18398 47572 18450
rect 47516 18338 47572 18398
rect 47516 18286 47518 18338
rect 47570 18286 47572 18338
rect 47516 18274 47572 18286
rect 47404 17938 47460 17948
rect 47628 17892 47684 18620
rect 47516 17836 47684 17892
rect 47740 18564 47796 18732
rect 47404 17780 47460 17790
rect 47516 17780 47572 17836
rect 47404 17778 47572 17780
rect 47404 17726 47406 17778
rect 47458 17726 47572 17778
rect 47404 17724 47572 17726
rect 47404 17714 47460 17724
rect 47180 17668 47236 17678
rect 46956 17612 47180 17668
rect 46732 16606 46734 16658
rect 46786 16606 46788 16658
rect 46732 16594 46788 16606
rect 45836 15762 46452 15764
rect 45836 15710 46174 15762
rect 46226 15710 46452 15762
rect 45836 15708 46452 15710
rect 47180 16546 47236 17612
rect 47516 16660 47572 17724
rect 47628 17668 47684 17678
rect 47740 17668 47796 18508
rect 47852 17778 47908 19628
rect 49084 18788 49140 19742
rect 49756 19684 49812 20638
rect 48860 18676 48916 18686
rect 47964 18564 48020 18574
rect 47964 18470 48020 18508
rect 48748 18564 48804 18574
rect 48860 18564 48916 18620
rect 48748 18562 48916 18564
rect 48748 18510 48750 18562
rect 48802 18510 48916 18562
rect 48748 18508 48916 18510
rect 48748 18498 48804 18508
rect 48412 18450 48468 18462
rect 48412 18398 48414 18450
rect 48466 18398 48468 18450
rect 48076 18338 48132 18350
rect 48076 18286 48078 18338
rect 48130 18286 48132 18338
rect 48076 17780 48132 18286
rect 48188 17892 48244 17902
rect 48188 17798 48244 17836
rect 47852 17726 47854 17778
rect 47906 17726 47908 17778
rect 47852 17714 47908 17726
rect 47964 17778 48132 17780
rect 47964 17726 48078 17778
rect 48130 17726 48132 17778
rect 47964 17724 48132 17726
rect 47628 17666 47796 17668
rect 47628 17614 47630 17666
rect 47682 17614 47796 17666
rect 47628 17612 47796 17614
rect 47628 17602 47684 17612
rect 47740 16772 47796 17612
rect 47516 16594 47572 16604
rect 47628 16716 47740 16772
rect 47180 16494 47182 16546
rect 47234 16494 47236 16546
rect 47180 15876 47236 16494
rect 45388 14866 45444 14878
rect 45388 14814 45390 14866
rect 45442 14814 45444 14866
rect 45388 14644 45444 14814
rect 45836 14756 45892 15708
rect 46172 15698 46228 15708
rect 47068 15652 47124 15662
rect 46956 15596 47068 15652
rect 45836 14662 45892 14700
rect 46284 14866 46340 14878
rect 46284 14814 46286 14866
rect 46338 14814 46340 14866
rect 46284 14754 46340 14814
rect 46956 14866 47012 15596
rect 47068 15558 47124 15596
rect 47180 15428 47236 15820
rect 47516 15876 47572 15886
rect 47628 15876 47684 16716
rect 47740 16706 47796 16716
rect 47516 15874 47684 15876
rect 47516 15822 47518 15874
rect 47570 15822 47684 15874
rect 47516 15820 47684 15822
rect 47516 15810 47572 15820
rect 46956 14814 46958 14866
rect 47010 14814 47012 14866
rect 46956 14802 47012 14814
rect 47068 15372 47236 15428
rect 46284 14702 46286 14754
rect 46338 14702 46340 14754
rect 46284 14690 46340 14702
rect 45388 14550 45444 14588
rect 44996 14476 45108 14532
rect 46396 14532 46452 14542
rect 44940 14438 44996 14476
rect 44268 14420 44324 14430
rect 44268 14326 44324 14364
rect 45612 14420 45668 14430
rect 45612 13858 45668 14364
rect 45612 13806 45614 13858
rect 45666 13806 45668 13858
rect 45612 13794 45668 13806
rect 44492 13746 44548 13758
rect 44492 13694 44494 13746
rect 44546 13694 44548 13746
rect 43820 13634 43876 13646
rect 43820 13582 43822 13634
rect 43874 13582 43876 13634
rect 43820 12852 43876 13582
rect 44044 12964 44100 12974
rect 44492 12964 44548 13694
rect 46396 13634 46452 14476
rect 46732 14420 46788 14430
rect 46732 14306 46788 14364
rect 46732 14254 46734 14306
rect 46786 14254 46788 14306
rect 46732 14242 46788 14254
rect 46396 13582 46398 13634
rect 46450 13582 46452 13634
rect 46396 13570 46452 13582
rect 44044 12962 44548 12964
rect 44044 12910 44046 12962
rect 44098 12910 44548 12962
rect 44044 12908 44548 12910
rect 44044 12898 44100 12908
rect 43820 12786 43876 12796
rect 46284 12852 46340 12862
rect 43484 11844 43540 12460
rect 44492 12628 44548 12638
rect 43596 11844 43652 11854
rect 43484 11842 43652 11844
rect 43484 11790 43598 11842
rect 43650 11790 43652 11842
rect 43484 11788 43652 11790
rect 42588 10836 42644 10846
rect 42588 10834 43092 10836
rect 42588 10782 42590 10834
rect 42642 10782 43092 10834
rect 42588 10780 43092 10782
rect 42588 10770 42644 10780
rect 42476 9662 42478 9714
rect 42530 9662 42532 9714
rect 42476 9650 42532 9662
rect 43036 9714 43092 10780
rect 43596 10500 43652 11788
rect 43596 10434 43652 10444
rect 44044 11732 44100 11742
rect 44044 10164 44100 11676
rect 44492 11730 44548 12572
rect 44940 12516 44996 12526
rect 44940 12422 44996 12460
rect 46284 11842 46340 12796
rect 47068 12516 47124 15372
rect 47180 14756 47236 14766
rect 47628 14756 47684 15820
rect 47964 15652 48020 17724
rect 48076 17714 48132 17724
rect 48412 17556 48468 18398
rect 49084 18450 49140 18732
rect 49420 19628 49756 19684
rect 49420 18564 49476 19628
rect 49756 19618 49812 19628
rect 49868 20692 49924 21420
rect 49420 18470 49476 18508
rect 49084 18398 49086 18450
rect 49138 18398 49140 18450
rect 48860 17556 48916 17566
rect 49084 17556 49140 18398
rect 49532 17892 49588 17902
rect 49532 17778 49588 17836
rect 49532 17726 49534 17778
rect 49586 17726 49588 17778
rect 49532 17714 49588 17726
rect 48412 17554 49140 17556
rect 48412 17502 48862 17554
rect 48914 17502 49140 17554
rect 48412 17500 49140 17502
rect 49868 17666 49924 20636
rect 49980 19684 50036 19694
rect 49980 19590 50036 19628
rect 50092 19458 50148 21646
rect 50204 20356 50260 22430
rect 50428 23100 50596 23156
rect 50428 21698 50484 23100
rect 50652 22484 50708 23998
rect 50876 23042 50932 25676
rect 51100 25620 51156 25630
rect 51100 25618 51380 25620
rect 51100 25566 51102 25618
rect 51154 25566 51380 25618
rect 51100 25564 51380 25566
rect 51100 25554 51156 25564
rect 51100 25394 51156 25406
rect 51100 25342 51102 25394
rect 51154 25342 51156 25394
rect 50988 24836 51044 24846
rect 50988 24722 51044 24780
rect 50988 24670 50990 24722
rect 51042 24670 51044 24722
rect 50988 24658 51044 24670
rect 50876 22990 50878 23042
rect 50930 22990 50932 23042
rect 50876 22978 50932 22990
rect 51100 23604 51156 25342
rect 51324 25394 51380 25564
rect 51324 25342 51326 25394
rect 51378 25342 51380 25394
rect 51212 24610 51268 24622
rect 51212 24558 51214 24610
rect 51266 24558 51268 24610
rect 51212 24500 51268 24558
rect 51212 24434 51268 24444
rect 51324 23828 51380 25342
rect 51324 23762 51380 23772
rect 50652 22482 50932 22484
rect 50652 22430 50654 22482
rect 50706 22430 50932 22482
rect 50652 22428 50932 22430
rect 50652 22418 50708 22428
rect 50556 22204 50820 22214
rect 50612 22148 50660 22204
rect 50716 22148 50764 22204
rect 50556 22138 50820 22148
rect 50876 21812 50932 22428
rect 50876 21746 50932 21756
rect 50428 21646 50430 21698
rect 50482 21646 50484 21698
rect 50428 21634 50484 21646
rect 50988 21700 51044 21710
rect 50540 20692 50596 20702
rect 50540 20598 50596 20636
rect 50876 20690 50932 20702
rect 50876 20638 50878 20690
rect 50930 20638 50932 20690
rect 50204 20290 50260 20300
rect 50556 20188 50820 20198
rect 50612 20132 50660 20188
rect 50716 20132 50764 20188
rect 50556 20122 50820 20132
rect 50876 19684 50932 20638
rect 50988 20468 51044 21644
rect 50988 20402 51044 20412
rect 50092 19406 50094 19458
rect 50146 19406 50148 19458
rect 50092 19394 50148 19406
rect 50652 19628 50876 19684
rect 49980 18900 50036 18910
rect 49980 18786 50036 18844
rect 49980 18734 49982 18786
rect 50034 18734 50036 18786
rect 49980 18722 50036 18734
rect 50092 18676 50148 18686
rect 50092 18582 50148 18620
rect 50652 18562 50708 19628
rect 50876 19618 50932 19628
rect 50652 18510 50654 18562
rect 50706 18510 50708 18562
rect 50652 18498 50708 18510
rect 50876 18788 50932 18798
rect 50876 18562 50932 18732
rect 50876 18510 50878 18562
rect 50930 18510 50932 18562
rect 50876 18498 50932 18510
rect 50556 18172 50820 18182
rect 50612 18116 50660 18172
rect 50716 18116 50764 18172
rect 50556 18106 50820 18116
rect 50540 18004 50596 18014
rect 50540 17890 50596 17948
rect 50540 17838 50542 17890
rect 50594 17838 50596 17890
rect 50540 17826 50596 17838
rect 51100 17778 51156 23548
rect 51212 23716 51268 23726
rect 51212 23602 51268 23660
rect 51212 23550 51214 23602
rect 51266 23550 51268 23602
rect 51212 23538 51268 23550
rect 51436 23492 51492 25900
rect 51548 25890 51604 25900
rect 51660 25394 51716 26684
rect 51660 25342 51662 25394
rect 51714 25342 51716 25394
rect 51660 25330 51716 25342
rect 51884 26738 51940 26750
rect 51884 26686 51886 26738
rect 51938 26686 51940 26738
rect 51436 23426 51492 23436
rect 51548 24836 51604 24846
rect 51548 22706 51604 24780
rect 51884 24500 51940 26686
rect 51996 26514 52052 27692
rect 52444 27746 52500 27758
rect 52444 27694 52446 27746
rect 52498 27694 52500 27746
rect 52444 27636 52500 27694
rect 52444 27570 52500 27580
rect 51996 26462 51998 26514
rect 52050 26462 52052 26514
rect 51996 26450 52052 26462
rect 52668 26852 52724 28588
rect 52780 28550 52836 28588
rect 53116 27972 53172 27982
rect 53116 27878 53172 27916
rect 53564 27858 53620 27870
rect 53564 27806 53566 27858
rect 53618 27806 53620 27858
rect 52780 27748 52836 27758
rect 52780 27654 52836 27692
rect 53116 27636 53172 27646
rect 53172 27580 53284 27636
rect 53116 27570 53172 27580
rect 52108 26066 52164 26078
rect 52108 26014 52110 26066
rect 52162 26014 52164 26066
rect 52108 25954 52164 26014
rect 52668 26066 52724 26796
rect 52668 26014 52670 26066
rect 52722 26014 52724 26066
rect 52668 26002 52724 26014
rect 52780 26516 52836 26526
rect 52108 25902 52110 25954
rect 52162 25902 52164 25954
rect 52108 25890 52164 25902
rect 52556 25618 52612 25630
rect 52556 25566 52558 25618
rect 52610 25566 52612 25618
rect 52556 25394 52612 25566
rect 52556 25342 52558 25394
rect 52610 25342 52612 25394
rect 52556 25330 52612 25342
rect 52108 24500 52164 24510
rect 51884 24498 52164 24500
rect 51884 24446 52110 24498
rect 52162 24446 52164 24498
rect 51884 24444 52164 24446
rect 51660 23828 51716 23838
rect 51660 23714 51716 23772
rect 51660 23662 51662 23714
rect 51714 23662 51716 23714
rect 51660 23650 51716 23662
rect 51772 23714 51828 23726
rect 52108 23716 52164 24444
rect 52780 24498 52836 26460
rect 53228 25060 53284 27580
rect 53564 26964 53620 27806
rect 53788 26964 53844 26974
rect 53564 26898 53620 26908
rect 53676 26908 53788 26964
rect 53564 26740 53620 26750
rect 53564 26646 53620 26684
rect 53676 26516 53732 26908
rect 53788 26898 53844 26908
rect 53676 26450 53732 26460
rect 54012 26740 54068 28812
rect 54236 28644 54292 30268
rect 54348 29876 54404 32620
rect 55020 32676 55076 32686
rect 55020 32582 55076 32620
rect 55020 31892 55076 31902
rect 55020 31805 55076 31836
rect 55020 31753 55022 31805
rect 55074 31753 55076 31805
rect 55020 31741 55076 31753
rect 54684 30660 54740 30670
rect 54684 30436 54740 30604
rect 55132 30546 55188 32732
rect 55692 32674 55748 33628
rect 56028 32900 56084 33740
rect 56700 33796 56756 33806
rect 56812 33796 56868 35308
rect 57372 34692 57428 35422
rect 57596 34804 57652 34814
rect 57708 34804 57764 36764
rect 57932 36708 57988 36718
rect 57932 36614 57988 36652
rect 58044 34804 58100 34814
rect 57596 34802 58212 34804
rect 57596 34750 57598 34802
rect 57650 34750 58046 34802
rect 58098 34750 58212 34802
rect 57596 34748 58212 34750
rect 57596 34738 57652 34748
rect 57260 34690 57428 34692
rect 57260 34638 57374 34690
rect 57426 34638 57428 34690
rect 57260 34636 57428 34638
rect 56756 33740 56868 33796
rect 56924 33906 56980 33918
rect 56924 33854 56926 33906
rect 56978 33854 56980 33906
rect 56364 32900 56420 32910
rect 56028 32844 56364 32900
rect 56364 32806 56420 32844
rect 55692 32622 55694 32674
rect 55746 32622 55748 32674
rect 55692 32610 55748 32622
rect 56700 32786 56756 33740
rect 56924 32900 56980 33854
rect 56924 32834 56980 32844
rect 57148 33908 57204 33918
rect 56700 32734 56702 32786
rect 56754 32734 56756 32786
rect 56252 32564 56308 32574
rect 56252 32470 56308 32508
rect 55580 32004 55636 32014
rect 55580 30882 55636 31948
rect 56028 31892 56084 31902
rect 55580 30830 55582 30882
rect 55634 30830 55636 30882
rect 55580 30818 55636 30830
rect 55804 31666 55860 31678
rect 55804 31614 55806 31666
rect 55858 31614 55860 31666
rect 55132 30494 55134 30546
rect 55186 30494 55188 30546
rect 54908 30436 54964 30446
rect 54684 30434 54964 30436
rect 54684 30382 54910 30434
rect 54962 30382 54964 30434
rect 54684 30380 54964 30382
rect 54348 29810 54404 29820
rect 54908 29650 54964 30380
rect 54908 29598 54910 29650
rect 54962 29598 54964 29650
rect 54796 28868 54852 28878
rect 54908 28868 54964 29598
rect 54852 28812 54964 28868
rect 54796 28802 54852 28812
rect 53340 25956 53396 25966
rect 53340 25954 53732 25956
rect 53340 25902 53342 25954
rect 53394 25902 53732 25954
rect 53340 25900 53732 25902
rect 53340 25890 53396 25900
rect 53228 25004 53508 25060
rect 53452 24724 53508 25004
rect 53676 24724 53732 25900
rect 54012 25844 54068 26684
rect 54124 28642 54292 28644
rect 54124 28590 54238 28642
rect 54290 28590 54292 28642
rect 54124 28588 54292 28590
rect 54124 26738 54180 28588
rect 54236 28578 54292 28588
rect 55132 28754 55188 30494
rect 55804 30434 55860 31614
rect 55804 30382 55806 30434
rect 55858 30382 55860 30434
rect 55804 30370 55860 30382
rect 56028 30546 56084 31836
rect 56028 30494 56030 30546
rect 56082 30494 56084 30546
rect 55132 28702 55134 28754
rect 55186 28702 55188 28754
rect 55132 28644 55188 28702
rect 55132 28578 55188 28588
rect 55804 29652 55860 29662
rect 56028 29652 56084 30494
rect 56700 31668 56756 32734
rect 56812 32676 56868 32686
rect 56812 32582 56868 32620
rect 57148 32674 57204 33852
rect 57148 32622 57150 32674
rect 57202 32622 57204 32674
rect 57148 32228 57204 32622
rect 56924 32172 57204 32228
rect 57260 32786 57316 34636
rect 57372 34626 57428 34636
rect 57708 33908 57764 34748
rect 58044 34738 58100 34748
rect 58156 34018 58212 34748
rect 58156 33966 58158 34018
rect 58210 33966 58212 34018
rect 58156 33954 58212 33966
rect 57708 33814 57764 33852
rect 57372 33684 57428 33694
rect 57372 33590 57428 33628
rect 57708 32900 57764 32910
rect 58156 32900 58212 32910
rect 57764 32898 58212 32900
rect 57764 32846 58158 32898
rect 58210 32846 58212 32898
rect 57764 32844 58212 32846
rect 57708 32806 57764 32844
rect 58156 32834 58212 32844
rect 57260 32734 57262 32786
rect 57314 32734 57316 32786
rect 56924 31892 56980 32172
rect 56924 31826 56980 31836
rect 57036 32004 57092 32014
rect 57260 31948 57316 32734
rect 57036 31892 57316 31948
rect 56700 30324 56756 31612
rect 56700 30258 56756 30268
rect 55804 29650 56084 29652
rect 55804 29598 55806 29650
rect 55858 29598 56084 29650
rect 55804 29596 56084 29598
rect 55804 28532 55860 29596
rect 55804 28466 55860 28476
rect 56924 28754 56980 28766
rect 56924 28702 56926 28754
rect 56978 28702 56980 28754
rect 56924 28532 56980 28702
rect 57036 28642 57092 31892
rect 57148 31668 57204 31678
rect 57148 31574 57204 31612
rect 57036 28590 57038 28642
rect 57090 28590 57092 28642
rect 57036 28532 57092 28590
rect 57036 28476 57316 28532
rect 56924 28420 56980 28476
rect 56924 28364 57092 28420
rect 54908 27860 54964 27870
rect 54908 27766 54964 27804
rect 56700 27858 56756 27870
rect 56700 27806 56702 27858
rect 56754 27806 56756 27858
rect 54236 27748 54292 27758
rect 55692 27748 55748 27758
rect 54236 27746 54404 27748
rect 54236 27694 54238 27746
rect 54290 27694 54404 27746
rect 54236 27692 54404 27694
rect 54236 27682 54292 27692
rect 54124 26686 54126 26738
rect 54178 26686 54180 26738
rect 54124 26292 54180 26686
rect 54348 26514 54404 27692
rect 55468 27692 55692 27748
rect 55468 27524 55524 27692
rect 55692 27654 55748 27692
rect 56588 27748 56644 27758
rect 56588 27654 56644 27692
rect 54348 26462 54350 26514
rect 54402 26462 54404 26514
rect 54348 26450 54404 26462
rect 55356 27468 55524 27524
rect 54124 26236 54516 26292
rect 54012 25750 54068 25788
rect 54460 25956 54516 26236
rect 54460 25730 54516 25900
rect 55020 25956 55076 25966
rect 55356 25956 55412 27468
rect 55804 26740 55860 26750
rect 55804 26646 55860 26684
rect 55020 25954 55300 25956
rect 55020 25902 55022 25954
rect 55074 25902 55300 25954
rect 55020 25900 55300 25902
rect 55020 25890 55076 25900
rect 54572 25844 54628 25854
rect 54628 25788 54740 25844
rect 54572 25778 54628 25788
rect 54460 25678 54462 25730
rect 54514 25678 54516 25730
rect 54460 25666 54516 25678
rect 53788 24724 53844 24734
rect 53452 24722 53620 24724
rect 53452 24670 53454 24722
rect 53506 24670 53620 24722
rect 53452 24668 53620 24670
rect 53676 24722 53844 24724
rect 53676 24670 53790 24722
rect 53842 24670 53844 24722
rect 53676 24668 53844 24670
rect 53452 24658 53508 24668
rect 53116 24612 53172 24622
rect 53116 24610 53284 24612
rect 53116 24558 53118 24610
rect 53170 24558 53284 24610
rect 53116 24556 53284 24558
rect 53116 24546 53172 24556
rect 52780 24446 52782 24498
rect 52834 24446 52836 24498
rect 52332 23826 52388 23838
rect 52332 23774 52334 23826
rect 52386 23774 52388 23826
rect 52332 23716 52388 23774
rect 51772 23662 51774 23714
rect 51826 23662 51828 23714
rect 51660 23492 51716 23502
rect 51772 23492 51828 23662
rect 51716 23436 51828 23492
rect 51996 23660 52388 23716
rect 52668 23828 52724 23838
rect 51660 23426 51716 23436
rect 51996 23380 52052 23660
rect 51548 22654 51550 22706
rect 51602 22654 51604 22706
rect 51548 22642 51604 22654
rect 51772 23324 52052 23380
rect 51324 22594 51380 22606
rect 51324 22542 51326 22594
rect 51378 22542 51380 22594
rect 51324 21364 51380 22542
rect 51324 21298 51380 21308
rect 51548 21698 51604 21710
rect 51548 21646 51550 21698
rect 51602 21646 51604 21698
rect 51548 20188 51604 21646
rect 51772 21700 51828 23324
rect 52668 22820 52724 23772
rect 52780 23716 52836 24446
rect 53228 23826 53284 24556
rect 53228 23774 53230 23826
rect 53282 23774 53284 23826
rect 53228 23762 53284 23774
rect 52780 23650 52836 23660
rect 53564 23492 53620 24668
rect 53788 24658 53844 24668
rect 54572 24612 54628 24622
rect 54460 24610 54628 24612
rect 54460 24558 54574 24610
rect 54626 24558 54628 24610
rect 54460 24556 54628 24558
rect 54124 24500 54180 24510
rect 54124 24406 54180 24444
rect 54460 23604 54516 24556
rect 54572 24546 54628 24556
rect 54684 24388 54740 25788
rect 55244 24722 55300 25900
rect 55244 24670 55246 24722
rect 55298 24670 55300 24722
rect 55244 24658 55300 24670
rect 55356 24612 55412 25900
rect 55580 25620 55636 25630
rect 55580 25526 55636 25564
rect 56028 25620 56084 25630
rect 56028 25526 56084 25564
rect 56700 25620 56756 27806
rect 56924 27860 56980 27870
rect 56924 27766 56980 27804
rect 57036 27860 57092 28364
rect 57260 27972 57316 28476
rect 57708 27972 57764 27982
rect 57260 27970 57764 27972
rect 57260 27918 57710 27970
rect 57762 27918 57764 27970
rect 57260 27916 57764 27918
rect 57148 27860 57204 27870
rect 57036 27858 57204 27860
rect 57036 27806 57150 27858
rect 57202 27806 57204 27858
rect 57036 27804 57204 27806
rect 56924 26628 56980 26638
rect 57036 26628 57092 27804
rect 57148 27794 57204 27804
rect 57260 27746 57316 27916
rect 57708 27906 57764 27916
rect 57260 27694 57262 27746
rect 57314 27694 57316 27746
rect 57260 26964 57316 27694
rect 58156 27748 58212 27758
rect 58156 27654 58212 27692
rect 57260 26738 57316 26908
rect 57260 26686 57262 26738
rect 57314 26686 57316 26738
rect 57260 26674 57316 26686
rect 56924 26626 57092 26628
rect 56924 26574 56926 26626
rect 56978 26574 57092 26626
rect 56924 26572 57092 26574
rect 56924 26562 56980 26572
rect 56700 25506 56756 25564
rect 56700 25454 56702 25506
rect 56754 25454 56756 25506
rect 56700 25442 56756 25454
rect 57148 25618 57204 25630
rect 57148 25566 57150 25618
rect 57202 25566 57204 25618
rect 57148 24948 57204 25566
rect 57036 24892 57204 24948
rect 57596 25618 57652 25630
rect 57596 25566 57598 25618
rect 57650 25566 57652 25618
rect 57596 25506 57652 25566
rect 57596 25454 57598 25506
rect 57650 25454 57652 25506
rect 55356 24546 55412 24556
rect 56812 24612 56868 24622
rect 57036 24612 57092 24892
rect 56868 24556 57092 24612
rect 57148 24724 57204 24734
rect 57596 24724 57652 25454
rect 57148 24722 57652 24724
rect 57148 24670 57150 24722
rect 57202 24670 57652 24722
rect 57148 24668 57652 24670
rect 55916 24500 55972 24510
rect 56700 24500 56756 24510
rect 55916 24498 56756 24500
rect 55916 24446 55918 24498
rect 55970 24446 56702 24498
rect 56754 24446 56756 24498
rect 55916 24444 56756 24446
rect 55916 24434 55972 24444
rect 56700 24434 56756 24444
rect 54572 24332 54740 24388
rect 54572 23714 54628 24332
rect 56700 24052 56756 24062
rect 56812 24052 56868 24556
rect 56700 24050 56868 24052
rect 56700 23998 56702 24050
rect 56754 23998 56868 24050
rect 56700 23996 56868 23998
rect 55692 23940 55748 23950
rect 55692 23938 55860 23940
rect 55692 23886 55694 23938
rect 55746 23886 55860 23938
rect 55692 23884 55860 23886
rect 55692 23874 55748 23884
rect 54572 23662 54574 23714
rect 54626 23662 54628 23714
rect 54572 23650 54628 23662
rect 54684 23828 54740 23838
rect 54684 23714 54740 23772
rect 54684 23662 54686 23714
rect 54738 23662 54740 23714
rect 54684 23650 54740 23662
rect 54460 23538 54516 23548
rect 55132 23604 55188 23614
rect 53564 23436 54068 23492
rect 52780 22820 52836 22830
rect 52668 22818 52836 22820
rect 52668 22766 52782 22818
rect 52834 22766 52836 22818
rect 52668 22764 52836 22766
rect 52780 22754 52836 22764
rect 54012 22706 54068 23436
rect 54012 22654 54014 22706
rect 54066 22654 54068 22706
rect 54012 22642 54068 22654
rect 51884 22594 51940 22606
rect 51884 22542 51886 22594
rect 51938 22542 51940 22594
rect 51884 22484 51940 22542
rect 53452 22596 53508 22606
rect 53228 22484 53284 22494
rect 51884 22418 51940 22428
rect 53004 22482 53284 22484
rect 53004 22430 53230 22482
rect 53282 22430 53284 22482
rect 53004 22428 53284 22430
rect 53004 21922 53060 22428
rect 53004 21870 53006 21922
rect 53058 21870 53060 21922
rect 53004 21858 53060 21870
rect 52220 21812 52276 21822
rect 51772 21634 51828 21644
rect 51884 21810 52276 21812
rect 51884 21758 52222 21810
rect 52274 21758 52276 21810
rect 51884 21756 52276 21758
rect 51884 21026 51940 21756
rect 52220 21746 52276 21756
rect 53228 21812 53284 22428
rect 51884 20974 51886 21026
rect 51938 20974 51940 21026
rect 51884 20962 51940 20974
rect 52892 21364 52948 21374
rect 51436 20132 51604 20188
rect 52220 20692 52276 20702
rect 51436 20018 51492 20132
rect 51436 19966 51438 20018
rect 51490 19966 51492 20018
rect 51436 19954 51492 19966
rect 52220 19794 52276 20636
rect 52892 19906 52948 21308
rect 52892 19854 52894 19906
rect 52946 19854 52948 19906
rect 52892 19842 52948 19854
rect 53116 20692 53172 20702
rect 52220 19742 52222 19794
rect 52274 19742 52276 19794
rect 52220 19730 52276 19742
rect 51548 19684 51604 19694
rect 51548 19590 51604 19628
rect 51884 19682 51940 19694
rect 51884 19630 51886 19682
rect 51938 19630 51940 19682
rect 51884 18786 51940 19630
rect 52556 19682 52612 19694
rect 52556 19630 52558 19682
rect 52610 19630 52612 19682
rect 52556 18900 52612 19630
rect 52556 18834 52612 18844
rect 52780 18898 52836 18910
rect 52780 18846 52782 18898
rect 52834 18846 52836 18898
rect 51884 18734 51886 18786
rect 51938 18734 51940 18786
rect 51884 18722 51940 18734
rect 52780 18786 52836 18846
rect 52780 18734 52782 18786
rect 52834 18734 52836 18786
rect 52780 18722 52836 18734
rect 53116 17890 53172 20636
rect 53228 20692 53284 21756
rect 53452 21586 53508 22540
rect 53452 21534 53454 21586
rect 53506 21534 53508 21586
rect 53452 21522 53508 21534
rect 53676 22594 53732 22606
rect 53676 22542 53678 22594
rect 53730 22542 53732 22594
rect 53564 20692 53620 20702
rect 53228 20690 53620 20692
rect 53228 20638 53566 20690
rect 53618 20638 53620 20690
rect 53228 20636 53620 20638
rect 53228 19684 53284 20636
rect 53564 20626 53620 20636
rect 53340 20468 53396 20478
rect 53676 20468 53732 22542
rect 54348 22596 54404 22606
rect 54348 22502 54404 22540
rect 55132 22594 55188 23548
rect 55804 22706 55860 23884
rect 56700 23938 56756 23996
rect 56700 23886 56702 23938
rect 56754 23886 56756 23938
rect 56700 23874 56756 23886
rect 57148 23602 57204 24668
rect 57820 24498 57876 24510
rect 57820 24446 57822 24498
rect 57874 24446 57876 24498
rect 57148 23550 57150 23602
rect 57202 23550 57204 23602
rect 57148 23490 57204 23550
rect 57148 23438 57150 23490
rect 57202 23438 57204 23490
rect 57148 23426 57204 23438
rect 57484 24052 57540 24062
rect 57820 24052 57876 24446
rect 57484 24050 57876 24052
rect 57484 23998 57486 24050
rect 57538 23998 57876 24050
rect 57484 23996 57876 23998
rect 55804 22654 55806 22706
rect 55858 22654 55860 22706
rect 55804 22642 55860 22654
rect 57484 22706 57540 23996
rect 57596 23604 57652 23614
rect 57596 23602 57876 23604
rect 57596 23550 57598 23602
rect 57650 23550 57876 23602
rect 57596 23548 57876 23550
rect 57596 23490 57652 23548
rect 57596 23438 57598 23490
rect 57650 23438 57652 23490
rect 57596 23426 57652 23438
rect 57820 22820 57876 23548
rect 58156 22820 58212 22830
rect 57820 22818 58212 22820
rect 57820 22766 58158 22818
rect 58210 22766 58212 22818
rect 57820 22764 58212 22766
rect 58156 22754 58212 22764
rect 57484 22654 57486 22706
rect 57538 22654 57540 22706
rect 55132 22542 55134 22594
rect 55186 22542 55188 22594
rect 55132 22530 55188 22542
rect 57260 22594 57316 22606
rect 57260 22542 57262 22594
rect 57314 22542 57316 22594
rect 54684 22484 54740 22494
rect 54684 22390 54740 22428
rect 56476 22484 56532 22494
rect 56476 22390 56532 22428
rect 57148 22484 57204 22494
rect 57148 22390 57204 22428
rect 54908 21924 54964 21934
rect 57260 21924 57316 22542
rect 54124 21700 54180 21710
rect 54124 20804 54180 21644
rect 54124 20738 54180 20748
rect 54908 20804 54964 21868
rect 57148 21868 57316 21924
rect 55244 21812 55300 21822
rect 55244 20804 55300 21756
rect 56700 21812 56756 21822
rect 57148 21812 57204 21868
rect 56700 21718 56756 21756
rect 57036 21756 57204 21812
rect 55468 21588 55524 21598
rect 56028 21588 56084 21598
rect 55468 21586 56084 21588
rect 55468 21534 55470 21586
rect 55522 21534 56030 21586
rect 56082 21534 56084 21586
rect 55468 21532 56084 21534
rect 55468 21522 55524 21532
rect 55356 20804 55412 20814
rect 55244 20802 55524 20804
rect 55244 20750 55358 20802
rect 55410 20750 55524 20802
rect 55244 20748 55524 20750
rect 54908 20710 54964 20748
rect 55356 20738 55412 20748
rect 53788 20692 53844 20702
rect 53788 20598 53844 20636
rect 54236 20468 54292 20478
rect 53676 20466 54292 20468
rect 53676 20414 54238 20466
rect 54290 20414 54292 20466
rect 53676 20412 54292 20414
rect 53340 20188 53396 20412
rect 54236 20402 54292 20412
rect 53340 20132 53508 20188
rect 53228 18898 53284 19628
rect 53228 18846 53230 18898
rect 53282 18846 53284 18898
rect 53228 18786 53284 18846
rect 53228 18734 53230 18786
rect 53282 18734 53284 18786
rect 53228 18722 53284 18734
rect 53452 19682 53508 20132
rect 54684 19794 54740 19806
rect 54684 19742 54686 19794
rect 54738 19742 54740 19794
rect 53452 19630 53454 19682
rect 53506 19630 53508 19682
rect 53452 18788 53508 19630
rect 54012 19682 54068 19694
rect 54012 19630 54014 19682
rect 54066 19630 54068 19682
rect 53676 18788 53732 18798
rect 53452 18786 53732 18788
rect 53452 18734 53678 18786
rect 53730 18734 53732 18786
rect 53452 18732 53732 18734
rect 53676 18722 53732 18732
rect 54012 18002 54068 19630
rect 54684 19010 54740 19742
rect 54684 18958 54686 19010
rect 54738 18958 54740 19010
rect 54684 18946 54740 18958
rect 55468 19570 55524 20748
rect 55804 20692 55860 21532
rect 56028 21476 56084 21532
rect 56028 21410 56084 21420
rect 57036 21588 57092 21756
rect 56252 20804 56308 20814
rect 56252 20710 56308 20748
rect 57036 20804 57092 21532
rect 57148 21588 57204 21598
rect 57484 21588 57540 22654
rect 57708 22706 57764 22718
rect 57708 22654 57710 22706
rect 57762 22654 57764 22706
rect 57708 21812 57764 22654
rect 57708 21746 57764 21756
rect 57148 21586 57540 21588
rect 57148 21534 57150 21586
rect 57202 21534 57540 21586
rect 57148 21532 57540 21534
rect 57148 21476 57204 21532
rect 57148 21410 57204 21420
rect 55804 20598 55860 20636
rect 55468 19518 55470 19570
rect 55522 19518 55524 19570
rect 55468 18564 55524 19518
rect 57036 18674 57092 20748
rect 57036 18622 57038 18674
rect 57090 18622 57092 18674
rect 57036 18610 57092 18622
rect 54012 17950 54014 18002
rect 54066 17950 54068 18002
rect 54012 17938 54068 17950
rect 55356 18508 55524 18564
rect 53116 17838 53118 17890
rect 53170 17838 53172 17890
rect 53116 17826 53172 17838
rect 51100 17726 51102 17778
rect 51154 17726 51156 17778
rect 51100 17714 51156 17726
rect 52332 17778 52388 17790
rect 52332 17726 52334 17778
rect 52386 17726 52388 17778
rect 49868 17614 49870 17666
rect 49922 17614 49924 17666
rect 47964 15558 48020 15596
rect 47180 14754 47684 14756
rect 47180 14702 47182 14754
rect 47234 14702 47630 14754
rect 47682 14702 47684 14754
rect 47180 14700 47684 14702
rect 47180 14532 47236 14700
rect 47628 14690 47684 14700
rect 48860 15538 48916 17500
rect 49308 16772 49364 16782
rect 48972 16660 49028 16670
rect 48972 16566 49028 16604
rect 49308 15874 49364 16716
rect 49756 16772 49812 16782
rect 49756 16658 49812 16716
rect 49756 16606 49758 16658
rect 49810 16606 49812 16658
rect 49756 16594 49812 16606
rect 49308 15822 49310 15874
rect 49362 15822 49364 15874
rect 49308 15810 49364 15822
rect 49756 15652 49812 15662
rect 49756 15558 49812 15596
rect 48860 15486 48862 15538
rect 48914 15486 48916 15538
rect 47180 14466 47236 14476
rect 48860 14420 48916 15486
rect 49308 14756 49364 14766
rect 49868 14756 49924 17614
rect 50204 17666 50260 17678
rect 50204 17614 50206 17666
rect 50258 17614 50260 17666
rect 50204 16770 50260 17614
rect 50204 16718 50206 16770
rect 50258 16718 50260 16770
rect 50204 16706 50260 16718
rect 51660 17666 51716 17678
rect 51660 17614 51662 17666
rect 51714 17614 51716 17666
rect 50316 16660 50372 16670
rect 50204 16324 50260 16334
rect 50204 15538 50260 16268
rect 50316 15988 50372 16604
rect 50764 16658 50820 16670
rect 50764 16606 50766 16658
rect 50818 16606 50820 16658
rect 50764 16324 50820 16606
rect 50764 16258 50820 16268
rect 50876 16660 50932 16670
rect 50556 16156 50820 16166
rect 50612 16100 50660 16156
rect 50716 16100 50764 16156
rect 50556 16090 50820 16100
rect 50316 15932 50596 15988
rect 50204 15486 50206 15538
rect 50258 15486 50260 15538
rect 49308 14754 49924 14756
rect 49308 14702 49310 14754
rect 49362 14702 49924 14754
rect 49308 14700 49924 14702
rect 49980 15204 50036 15214
rect 49308 14690 49364 14700
rect 48860 14354 48916 14364
rect 47180 14306 47236 14318
rect 47180 14254 47182 14306
rect 47234 14254 47236 14306
rect 47180 13746 47236 14254
rect 47180 13694 47182 13746
rect 47234 13694 47236 13746
rect 47180 13682 47236 13694
rect 47852 13524 47908 13534
rect 47740 13522 47908 13524
rect 47740 13470 47854 13522
rect 47906 13470 47908 13522
rect 47740 13468 47908 13470
rect 47740 12852 47796 13468
rect 47852 13458 47908 13468
rect 47740 12758 47796 12796
rect 49980 12628 50036 15148
rect 50092 14420 50148 14430
rect 50204 14420 50260 15486
rect 50540 15316 50596 15932
rect 50540 14754 50596 15260
rect 50764 15876 50820 15886
rect 50876 15876 50932 16604
rect 51212 16548 51268 16558
rect 50764 15874 50932 15876
rect 50764 15822 50766 15874
rect 50818 15822 50932 15874
rect 50764 15820 50932 15822
rect 51100 16546 51268 16548
rect 51100 16494 51214 16546
rect 51266 16494 51268 16546
rect 51100 16492 51268 16494
rect 50764 15204 50820 15820
rect 50764 15138 50820 15148
rect 50988 15652 51044 15662
rect 51100 15652 51156 16492
rect 51212 16482 51268 16492
rect 51660 16436 51716 17614
rect 51660 16370 51716 16380
rect 51772 16324 51828 16334
rect 51772 15986 51828 16268
rect 51772 15934 51774 15986
rect 51826 15934 51828 15986
rect 51212 15876 51268 15886
rect 51212 15782 51268 15820
rect 51772 15764 51828 15934
rect 52332 15988 52388 17726
rect 53340 17668 53396 17678
rect 53228 17666 53396 17668
rect 53228 17614 53342 17666
rect 53394 17614 53396 17666
rect 53228 17612 53396 17614
rect 52556 16660 52612 16698
rect 52556 16594 52612 16604
rect 52892 16546 52948 16558
rect 52892 16494 52894 16546
rect 52946 16494 52948 16546
rect 52556 16436 52612 16446
rect 52556 16342 52612 16380
rect 52780 15988 52836 15998
rect 52332 15986 52836 15988
rect 52332 15934 52782 15986
rect 52834 15934 52836 15986
rect 52332 15932 52836 15934
rect 52780 15922 52836 15932
rect 52892 15876 52948 16494
rect 52892 15810 52948 15820
rect 53228 16436 53284 17612
rect 53340 17602 53396 17612
rect 55356 16772 55412 18508
rect 55580 16772 55636 16782
rect 55356 16770 55636 16772
rect 55356 16718 55582 16770
rect 55634 16718 55636 16770
rect 55356 16716 55636 16718
rect 51772 15698 51828 15708
rect 52780 15764 52836 15774
rect 51044 15596 51156 15652
rect 52556 15650 52612 15662
rect 52556 15598 52558 15650
rect 52610 15598 52612 15650
rect 50540 14702 50542 14754
rect 50594 14702 50596 14754
rect 50540 14690 50596 14702
rect 50988 14756 51044 15596
rect 50988 14662 51044 14700
rect 51660 15316 51716 15326
rect 51660 14754 51716 15260
rect 51660 14702 51662 14754
rect 51714 14702 51716 14754
rect 51660 14690 51716 14702
rect 52108 14756 52164 14766
rect 52108 14662 52164 14700
rect 50148 14364 50260 14420
rect 52556 14644 52612 15598
rect 52780 14754 52836 15708
rect 52780 14702 52782 14754
rect 52834 14702 52836 14754
rect 52780 14690 52836 14702
rect 50092 14326 50148 14364
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 51212 13860 51268 13870
rect 51212 13766 51268 13804
rect 52444 13860 52500 13870
rect 52556 13860 52612 14588
rect 53228 14644 53284 16380
rect 53564 16546 53620 16558
rect 53564 16494 53566 16546
rect 53618 16494 53620 16546
rect 53340 15652 53396 15662
rect 53564 15652 53620 16494
rect 53340 15650 53620 15652
rect 53340 15598 53342 15650
rect 53394 15598 53620 15650
rect 53340 15596 53620 15598
rect 54236 16546 54292 16558
rect 54236 16494 54238 16546
rect 54290 16494 54292 16546
rect 54236 15652 54292 16494
rect 54572 16434 54628 16446
rect 54572 16382 54574 16434
rect 54626 16382 54628 16434
rect 54572 15764 54628 16382
rect 54908 16436 54964 16446
rect 55356 16436 55412 16716
rect 55580 16706 55636 16716
rect 54964 16380 55412 16436
rect 54908 16342 54964 16380
rect 54572 15698 54628 15708
rect 53340 15316 53396 15596
rect 54236 15558 54292 15596
rect 53340 15250 53396 15260
rect 53228 14550 53284 14588
rect 52500 13804 52612 13860
rect 52444 13794 52500 13804
rect 49980 12534 50036 12572
rect 47068 12450 47124 12460
rect 47964 12516 48020 12526
rect 48188 12516 48244 12526
rect 48020 12514 48244 12516
rect 48020 12462 48190 12514
rect 48242 12462 48244 12514
rect 48020 12460 48244 12462
rect 47964 12450 48020 12460
rect 48188 12450 48244 12460
rect 50556 12124 50820 12134
rect 50612 12068 50660 12124
rect 50716 12068 50764 12124
rect 50556 12058 50820 12068
rect 46284 11790 46286 11842
rect 46338 11790 46340 11842
rect 46284 11778 46340 11790
rect 44492 11678 44494 11730
rect 44546 11678 44548 11730
rect 44492 11666 44548 11678
rect 46620 11732 46676 11742
rect 46620 11638 46676 11676
rect 48076 11618 48132 11630
rect 48076 11566 48078 11618
rect 48130 11566 48132 11618
rect 48076 10500 48132 11566
rect 48076 10434 48132 10444
rect 43036 9662 43038 9714
rect 43090 9662 43092 9714
rect 43036 9650 43092 9662
rect 43596 10108 44100 10164
rect 50556 10108 50820 10118
rect 42028 8708 42084 8718
rect 42028 8614 42084 8652
rect 41804 8542 41806 8594
rect 41858 8542 41860 8594
rect 41020 7758 41022 7810
rect 41074 7758 41076 7810
rect 41020 7746 41076 7758
rect 41468 8484 41524 8494
rect 41804 8484 41860 8542
rect 43260 8596 43316 8606
rect 43596 8596 43652 10108
rect 50612 10052 50660 10108
rect 50716 10052 50764 10108
rect 50556 10042 50820 10052
rect 43708 9716 43764 9726
rect 43708 9714 44100 9716
rect 43708 9662 43710 9714
rect 43762 9662 44100 9714
rect 43708 9660 44100 9662
rect 43708 9650 43764 9660
rect 44044 8930 44100 9660
rect 44044 8878 44046 8930
rect 44098 8878 44100 8930
rect 44044 8866 44100 8878
rect 43316 8540 43652 8596
rect 43260 8502 43316 8540
rect 41524 8428 41860 8484
rect 42252 8482 42308 8494
rect 42252 8430 42254 8482
rect 42306 8430 42308 8482
rect 42252 8428 42308 8430
rect 41468 7810 41524 8428
rect 41468 7758 41470 7810
rect 41522 7758 41524 7810
rect 41468 7746 41524 7758
rect 41916 8372 42308 8428
rect 41916 7810 41972 8316
rect 50556 8092 50820 8102
rect 50612 8036 50660 8092
rect 50716 8036 50764 8092
rect 50556 8026 50820 8036
rect 41916 7758 41918 7810
rect 41970 7758 41972 7810
rect 41916 7746 41972 7758
rect 34524 7700 34580 7710
rect 34412 7698 34580 7700
rect 34412 7646 34526 7698
rect 34578 7646 34580 7698
rect 34412 7644 34580 7646
rect 34524 7634 34580 7644
rect 35868 7698 35924 7710
rect 35868 7646 35870 7698
rect 35922 7646 35924 7698
rect 33740 7588 33796 7598
rect 35196 7588 35252 7598
rect 33740 7494 33796 7532
rect 35084 7586 35252 7588
rect 35084 7534 35198 7586
rect 35250 7534 35252 7586
rect 35084 7532 35252 7534
rect 33852 6692 33908 6702
rect 33516 6636 33684 6692
rect 33628 6580 33684 6636
rect 33628 6486 33684 6524
rect 33852 6578 33908 6636
rect 33852 6526 33854 6578
rect 33906 6526 33908 6578
rect 33852 6514 33908 6526
rect 34972 6468 35028 6478
rect 34972 6374 35028 6412
rect 33628 6356 33684 6366
rect 33292 6354 33684 6356
rect 33292 6302 33630 6354
rect 33682 6302 33684 6354
rect 33292 6300 33684 6302
rect 33628 5572 33684 6300
rect 33068 5570 33348 5572
rect 33068 5518 33070 5570
rect 33122 5518 33348 5570
rect 33068 5516 33348 5518
rect 33068 5506 33124 5516
rect 31500 5406 31502 5458
rect 31554 5406 31556 5458
rect 31500 5394 31556 5406
rect 28924 4622 28926 4674
rect 28978 4622 28980 4674
rect 28924 4610 28980 4622
rect 32396 4898 32452 4910
rect 32396 4846 32398 4898
rect 32450 4846 32452 4898
rect 32396 4674 32452 4846
rect 32396 4622 32398 4674
rect 32450 4622 32452 4674
rect 32396 4610 32452 4622
rect 32844 4898 32900 4910
rect 32844 4846 32846 4898
rect 32898 4846 32900 4898
rect 32844 4674 32900 4846
rect 32844 4622 32846 4674
rect 32898 4622 32900 4674
rect 32844 4610 32900 4622
rect 33292 4676 33348 5516
rect 33516 5570 33684 5572
rect 33516 5518 33630 5570
rect 33682 5518 33684 5570
rect 33516 5516 33684 5518
rect 33516 4898 33572 5516
rect 33628 5506 33684 5516
rect 35084 5460 35140 7532
rect 35196 7522 35252 7532
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35756 6916 35812 6926
rect 35868 6916 35924 7646
rect 35756 6914 35924 6916
rect 35756 6862 35758 6914
rect 35810 6862 35924 6914
rect 35756 6860 35924 6862
rect 35756 6850 35812 6860
rect 50556 6076 50820 6086
rect 50612 6020 50660 6076
rect 50716 6020 50764 6076
rect 50556 6010 50820 6020
rect 35196 5460 35252 5470
rect 35084 5404 35196 5460
rect 35196 5394 35252 5404
rect 36092 5460 36148 5470
rect 36092 5366 36148 5404
rect 35196 5068 35460 5078
rect 35252 5012 35300 5068
rect 35356 5012 35404 5068
rect 35196 5002 35460 5012
rect 33516 4846 33518 4898
rect 33570 4846 33572 4898
rect 33516 4834 33572 4846
rect 33740 4676 33796 4686
rect 33292 4674 33796 4676
rect 33292 4622 33294 4674
rect 33346 4622 33742 4674
rect 33794 4622 33796 4674
rect 33292 4620 33796 4622
rect 33292 4610 33348 4620
rect 33740 4610 33796 4620
rect 19836 4060 20100 4070
rect 19892 4004 19940 4060
rect 19996 4004 20044 4060
rect 19836 3994 20100 4004
rect 50556 4060 50820 4070
rect 50612 4004 50660 4060
rect 50716 4004 50764 4060
rect 50556 3994 50820 4004
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
<< via2 >>
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 4476 55466 4532 55468
rect 4476 55414 4478 55466
rect 4478 55414 4530 55466
rect 4530 55414 4532 55466
rect 4476 55412 4532 55414
rect 4580 55466 4636 55468
rect 4580 55414 4582 55466
rect 4582 55414 4634 55466
rect 4634 55414 4636 55466
rect 4580 55412 4636 55414
rect 4684 55466 4740 55468
rect 4684 55414 4686 55466
rect 4686 55414 4738 55466
rect 4738 55414 4740 55466
rect 4684 55412 4740 55414
rect 19836 54458 19892 54460
rect 19836 54406 19838 54458
rect 19838 54406 19890 54458
rect 19890 54406 19892 54458
rect 19836 54404 19892 54406
rect 19940 54458 19996 54460
rect 19940 54406 19942 54458
rect 19942 54406 19994 54458
rect 19994 54406 19996 54458
rect 19940 54404 19996 54406
rect 20044 54458 20100 54460
rect 20044 54406 20046 54458
rect 20046 54406 20098 54458
rect 20098 54406 20100 54458
rect 20044 54404 20100 54406
rect 4476 53450 4532 53452
rect 4476 53398 4478 53450
rect 4478 53398 4530 53450
rect 4530 53398 4532 53450
rect 4476 53396 4532 53398
rect 4580 53450 4636 53452
rect 4580 53398 4582 53450
rect 4582 53398 4634 53450
rect 4634 53398 4636 53450
rect 4580 53396 4636 53398
rect 4684 53450 4740 53452
rect 4684 53398 4686 53450
rect 4686 53398 4738 53450
rect 4738 53398 4740 53450
rect 4684 53396 4740 53398
rect 19836 52442 19892 52444
rect 19836 52390 19838 52442
rect 19838 52390 19890 52442
rect 19890 52390 19892 52442
rect 19836 52388 19892 52390
rect 19940 52442 19996 52444
rect 19940 52390 19942 52442
rect 19942 52390 19994 52442
rect 19994 52390 19996 52442
rect 19940 52388 19996 52390
rect 20044 52442 20100 52444
rect 20044 52390 20046 52442
rect 20046 52390 20098 52442
rect 20098 52390 20100 52442
rect 20044 52388 20100 52390
rect 5852 52162 5908 52164
rect 5852 52110 5854 52162
rect 5854 52110 5906 52162
rect 5906 52110 5908 52162
rect 5852 52108 5908 52110
rect 4476 51434 4532 51436
rect 4476 51382 4478 51434
rect 4478 51382 4530 51434
rect 4530 51382 4532 51434
rect 4476 51380 4532 51382
rect 4580 51434 4636 51436
rect 4580 51382 4582 51434
rect 4582 51382 4634 51434
rect 4634 51382 4636 51434
rect 4580 51380 4636 51382
rect 4684 51434 4740 51436
rect 4684 51382 4686 51434
rect 4686 51382 4738 51434
rect 4738 51382 4740 51434
rect 4684 51380 4740 51382
rect 19836 50426 19892 50428
rect 19836 50374 19838 50426
rect 19838 50374 19890 50426
rect 19890 50374 19892 50426
rect 19836 50372 19892 50374
rect 19940 50426 19996 50428
rect 19940 50374 19942 50426
rect 19942 50374 19994 50426
rect 19994 50374 19996 50426
rect 19940 50372 19996 50374
rect 20044 50426 20100 50428
rect 20044 50374 20046 50426
rect 20046 50374 20098 50426
rect 20098 50374 20100 50426
rect 20044 50372 20100 50374
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 19836 48410 19892 48412
rect 19836 48358 19838 48410
rect 19838 48358 19890 48410
rect 19890 48358 19892 48410
rect 19836 48356 19892 48358
rect 19940 48410 19996 48412
rect 19940 48358 19942 48410
rect 19942 48358 19994 48410
rect 19994 48358 19996 48410
rect 19940 48356 19996 48358
rect 20044 48410 20100 48412
rect 20044 48358 20046 48410
rect 20046 48358 20098 48410
rect 20098 48358 20100 48410
rect 20044 48356 20100 48358
rect 1708 45276 1764 45332
rect 3052 45276 3108 45332
rect 1820 44380 1876 44436
rect 2380 44604 2436 44660
rect 4476 47402 4532 47404
rect 4476 47350 4478 47402
rect 4478 47350 4530 47402
rect 4530 47350 4532 47402
rect 4476 47348 4532 47350
rect 4580 47402 4636 47404
rect 4580 47350 4582 47402
rect 4582 47350 4634 47402
rect 4634 47350 4636 47402
rect 4580 47348 4636 47350
rect 4684 47402 4740 47404
rect 4684 47350 4686 47402
rect 4686 47350 4738 47402
rect 4738 47350 4740 47402
rect 4684 47348 4740 47350
rect 3948 46956 4004 47012
rect 4508 46956 4564 47012
rect 5628 47010 5684 47012
rect 5628 46958 5630 47010
rect 5630 46958 5682 47010
rect 5682 46958 5684 47010
rect 5628 46956 5684 46958
rect 24668 47794 24724 47796
rect 24668 47742 24670 47794
rect 24670 47742 24722 47794
rect 24722 47742 24724 47794
rect 24668 47740 24724 47742
rect 4172 45778 4228 45780
rect 4172 45726 4174 45778
rect 4174 45726 4226 45778
rect 4226 45726 4228 45778
rect 4172 45724 4228 45726
rect 4476 45386 4532 45388
rect 4476 45334 4478 45386
rect 4478 45334 4530 45386
rect 4530 45334 4532 45386
rect 4476 45332 4532 45334
rect 4580 45386 4636 45388
rect 4580 45334 4582 45386
rect 4582 45334 4634 45386
rect 4634 45334 4636 45386
rect 4580 45332 4636 45334
rect 4684 45386 4740 45388
rect 4684 45334 4686 45386
rect 4686 45334 4738 45386
rect 4738 45334 4740 45386
rect 4684 45332 4740 45334
rect 4172 45276 4228 45332
rect 19836 46394 19892 46396
rect 19836 46342 19838 46394
rect 19838 46342 19890 46394
rect 19890 46342 19892 46394
rect 19836 46340 19892 46342
rect 19940 46394 19996 46396
rect 19940 46342 19942 46394
rect 19942 46342 19994 46394
rect 19994 46342 19996 46394
rect 19940 46340 19996 46342
rect 20044 46394 20100 46396
rect 20044 46342 20046 46394
rect 20046 46342 20098 46394
rect 20098 46342 20100 46394
rect 20044 46340 20100 46342
rect 6188 45724 6244 45780
rect 7196 45724 7252 45780
rect 3388 44604 3444 44660
rect 1932 43148 1988 43204
rect 4476 43370 4532 43372
rect 4476 43318 4478 43370
rect 4478 43318 4530 43370
rect 4530 43318 4532 43370
rect 4476 43316 4532 43318
rect 4580 43370 4636 43372
rect 4580 43318 4582 43370
rect 4582 43318 4634 43370
rect 4634 43318 4636 43370
rect 4580 43316 4636 43318
rect 4684 43370 4740 43372
rect 4684 43318 4686 43370
rect 4686 43318 4738 43370
rect 4738 43318 4740 43370
rect 4684 43316 4740 43318
rect 2716 43148 2772 43204
rect 5740 45612 5796 45668
rect 7644 45666 7700 45668
rect 7644 45614 7646 45666
rect 7646 45614 7698 45666
rect 7698 45614 7700 45666
rect 7644 45612 7700 45614
rect 8764 45612 8820 45668
rect 6076 45500 6132 45556
rect 8316 45554 8372 45556
rect 8316 45502 8318 45554
rect 8318 45502 8370 45554
rect 8370 45502 8372 45554
rect 8316 45500 8372 45502
rect 6076 44604 6132 44660
rect 4956 42812 5012 42868
rect 5628 43202 5684 43204
rect 5628 43150 5630 43202
rect 5630 43150 5682 43202
rect 5682 43150 5684 43202
rect 5628 43148 5684 43150
rect 6636 44882 6692 44884
rect 6636 44830 6638 44882
rect 6638 44830 6690 44882
rect 6690 44830 6692 44882
rect 6636 44828 6692 44830
rect 8540 44098 8596 44100
rect 8540 44046 8542 44098
rect 8542 44046 8594 44098
rect 8594 44046 8596 44098
rect 8540 44044 8596 44046
rect 9660 45778 9716 45780
rect 9660 45726 9662 45778
rect 9662 45726 9714 45778
rect 9714 45726 9716 45778
rect 9660 45724 9716 45726
rect 9548 44940 9604 44996
rect 9212 44658 9268 44660
rect 9212 44606 9214 44658
rect 9214 44606 9266 44658
rect 9266 44606 9268 44658
rect 9212 44604 9268 44606
rect 10220 44940 10276 44996
rect 9660 44882 9716 44884
rect 9660 44830 9662 44882
rect 9662 44830 9714 44882
rect 9714 44830 9716 44882
rect 9660 44828 9716 44830
rect 11676 45052 11732 45108
rect 12796 45106 12852 45108
rect 12796 45054 12798 45106
rect 12798 45054 12850 45106
rect 12850 45054 12852 45106
rect 12796 45052 12852 45054
rect 11564 44940 11620 44996
rect 10332 44604 10388 44660
rect 9884 44098 9940 44100
rect 9884 44046 9886 44098
rect 9886 44046 9938 44098
rect 9938 44046 9940 44098
rect 9884 44044 9940 44046
rect 6188 42866 6244 42868
rect 6188 42814 6190 42866
rect 6190 42814 6242 42866
rect 6242 42814 6244 42866
rect 6188 42812 6244 42814
rect 2380 41916 2436 41972
rect 3388 41970 3444 41972
rect 3388 41918 3390 41970
rect 3390 41918 3442 41970
rect 3442 41918 3444 41970
rect 3388 41916 3444 41918
rect 1708 40908 1764 40964
rect 1820 41468 1876 41524
rect 2380 40908 2436 40964
rect 1820 40348 1876 40404
rect 3052 40348 3108 40404
rect 5740 41580 5796 41636
rect 4396 41468 4452 41524
rect 5628 41468 5684 41524
rect 4476 41354 4532 41356
rect 4476 41302 4478 41354
rect 4478 41302 4530 41354
rect 4530 41302 4532 41354
rect 4476 41300 4532 41302
rect 4580 41354 4636 41356
rect 4580 41302 4582 41354
rect 4582 41302 4634 41354
rect 4634 41302 4636 41354
rect 4580 41300 4636 41302
rect 4684 41354 4740 41356
rect 4684 41302 4686 41354
rect 4686 41302 4738 41354
rect 4738 41302 4740 41354
rect 4684 41300 4740 41302
rect 6076 40962 6132 40964
rect 6076 40910 6078 40962
rect 6078 40910 6130 40962
rect 6130 40910 6132 40962
rect 6076 40908 6132 40910
rect 3836 39900 3892 39956
rect 4060 40348 4116 40404
rect 4956 40626 5012 40628
rect 4956 40574 4958 40626
rect 4958 40574 5010 40626
rect 5010 40574 5012 40626
rect 4956 40572 5012 40574
rect 6188 40626 6244 40628
rect 6188 40574 6190 40626
rect 6190 40574 6242 40626
rect 6242 40574 6244 40626
rect 6188 40572 6244 40574
rect 19836 44378 19892 44380
rect 19836 44326 19838 44378
rect 19838 44326 19890 44378
rect 19890 44326 19892 44378
rect 19836 44324 19892 44326
rect 19940 44378 19996 44380
rect 19940 44326 19942 44378
rect 19942 44326 19994 44378
rect 19994 44326 19996 44378
rect 19940 44324 19996 44326
rect 20044 44378 20100 44380
rect 20044 44326 20046 44378
rect 20046 44326 20098 44378
rect 20098 44326 20100 44378
rect 20044 44324 20100 44326
rect 12348 44044 12404 44100
rect 10892 43932 10948 43988
rect 10780 43148 10836 43204
rect 6972 41634 7028 41636
rect 6972 41582 6974 41634
rect 6974 41582 7026 41634
rect 7026 41582 7028 41634
rect 6972 41580 7028 41582
rect 11452 43148 11508 43204
rect 12348 43596 12404 43652
rect 12796 43820 12852 43876
rect 14476 43986 14532 43988
rect 14476 43934 14478 43986
rect 14478 43934 14530 43986
rect 14530 43934 14532 43986
rect 14476 43932 14532 43934
rect 14588 43874 14644 43876
rect 14588 43822 14590 43874
rect 14590 43822 14642 43874
rect 14642 43822 14644 43874
rect 14588 43820 14644 43822
rect 13468 43596 13524 43652
rect 9660 41580 9716 41636
rect 10220 40684 10276 40740
rect 9324 40626 9380 40628
rect 9324 40574 9326 40626
rect 9326 40574 9378 40626
rect 9378 40574 9380 40626
rect 9324 40572 9380 40574
rect 11340 41580 11396 41636
rect 10444 40572 10500 40628
rect 6860 40236 6916 40292
rect 4956 39900 5012 39956
rect 3836 38668 3892 38724
rect 2716 36034 2772 36036
rect 2716 35982 2718 36034
rect 2718 35982 2770 36034
rect 2770 35982 2772 36034
rect 2716 35980 2772 35982
rect 3164 35980 3220 36036
rect 4284 39676 4340 39732
rect 4476 39338 4532 39340
rect 4476 39286 4478 39338
rect 4478 39286 4530 39338
rect 4530 39286 4532 39338
rect 4476 39284 4532 39286
rect 4580 39338 4636 39340
rect 4580 39286 4582 39338
rect 4582 39286 4634 39338
rect 4634 39286 4636 39338
rect 4580 39284 4636 39286
rect 4684 39338 4740 39340
rect 4684 39286 4686 39338
rect 4686 39286 4738 39338
rect 4738 39286 4740 39338
rect 4684 39284 4740 39286
rect 4620 38722 4676 38724
rect 4620 38670 4622 38722
rect 4622 38670 4674 38722
rect 4674 38670 4676 38722
rect 4620 38668 4676 38670
rect 4956 39170 5012 39172
rect 4956 39118 4958 39170
rect 4958 39118 5010 39170
rect 5010 39118 5012 39170
rect 4956 39116 5012 39118
rect 6076 38668 6132 38724
rect 10780 40684 10836 40740
rect 13468 43202 13524 43204
rect 13468 43150 13470 43202
rect 13470 43150 13522 43202
rect 13522 43150 13524 43202
rect 13468 43148 13524 43150
rect 20188 43762 20244 43764
rect 20188 43710 20190 43762
rect 20190 43710 20242 43762
rect 20242 43710 20244 43762
rect 20188 43708 20244 43710
rect 21644 43708 21700 43764
rect 22204 44994 22260 44996
rect 22204 44942 22206 44994
rect 22206 44942 22258 44994
rect 22258 44942 22260 44994
rect 22204 44940 22260 44942
rect 22764 44828 22820 44884
rect 25004 45724 25060 45780
rect 22204 43820 22260 43876
rect 13356 42588 13412 42644
rect 16716 42642 16772 42644
rect 16716 42590 16718 42642
rect 16718 42590 16770 42642
rect 16770 42590 16772 42642
rect 16716 42588 16772 42590
rect 12796 40626 12852 40628
rect 12796 40574 12798 40626
rect 12798 40574 12850 40626
rect 12850 40574 12852 40626
rect 12796 40572 12852 40574
rect 14364 41634 14420 41636
rect 14364 41582 14366 41634
rect 14366 41582 14418 41634
rect 14418 41582 14420 41634
rect 14364 41580 14420 41582
rect 13468 40738 13524 40740
rect 13468 40686 13470 40738
rect 13470 40686 13522 40738
rect 13522 40686 13524 40738
rect 13468 40684 13524 40686
rect 13580 40626 13636 40628
rect 13580 40574 13582 40626
rect 13582 40574 13634 40626
rect 13634 40574 13636 40626
rect 13580 40572 13636 40574
rect 17836 42364 17892 42420
rect 17612 40796 17668 40852
rect 11340 39842 11396 39844
rect 11340 39790 11342 39842
rect 11342 39790 11394 39842
rect 11394 39790 11396 39842
rect 11340 39788 11396 39790
rect 11676 39788 11732 39844
rect 6860 38668 6916 38724
rect 4844 38220 4900 38276
rect 5516 38220 5572 38276
rect 4284 37772 4340 37828
rect 4476 37322 4532 37324
rect 4476 37270 4478 37322
rect 4478 37270 4530 37322
rect 4530 37270 4532 37322
rect 4476 37268 4532 37270
rect 4580 37322 4636 37324
rect 4580 37270 4582 37322
rect 4582 37270 4634 37322
rect 4634 37270 4636 37322
rect 4580 37268 4636 37270
rect 4684 37322 4740 37324
rect 4684 37270 4686 37322
rect 4686 37270 4738 37322
rect 4738 37270 4740 37322
rect 4684 37268 4740 37270
rect 4508 37100 4564 37156
rect 7084 38220 7140 38276
rect 6300 38108 6356 38164
rect 2380 34860 2436 34916
rect 4956 36594 5012 36596
rect 4956 36542 4958 36594
rect 4958 36542 5010 36594
rect 5010 36542 5012 36594
rect 4956 36540 5012 36542
rect 4060 35980 4116 36036
rect 3052 34860 3108 34916
rect 4172 36316 4228 36372
rect 8316 39116 8372 39172
rect 7532 38162 7588 38164
rect 7532 38110 7534 38162
rect 7534 38110 7586 38162
rect 7586 38110 7588 38162
rect 7532 38108 7588 38110
rect 8876 38108 8932 38164
rect 6636 37100 6692 37156
rect 12684 39788 12740 39844
rect 12796 39564 12852 39620
rect 13916 39618 13972 39620
rect 13916 39566 13918 39618
rect 13918 39566 13970 39618
rect 13970 39566 13972 39618
rect 13916 39564 13972 39566
rect 12236 38668 12292 38724
rect 13468 38722 13524 38724
rect 13468 38670 13470 38722
rect 13470 38670 13522 38722
rect 13522 38670 13524 38722
rect 13468 38668 13524 38670
rect 7644 36876 7700 36932
rect 8764 36930 8820 36932
rect 8764 36878 8766 36930
rect 8766 36878 8818 36930
rect 8818 36878 8820 36930
rect 8764 36876 8820 36878
rect 6188 36540 6244 36596
rect 8316 36594 8372 36596
rect 8316 36542 8318 36594
rect 8318 36542 8370 36594
rect 8370 36542 8372 36594
rect 8316 36540 8372 36542
rect 11004 36594 11060 36596
rect 11004 36542 11006 36594
rect 11006 36542 11058 36594
rect 11058 36542 11060 36594
rect 11004 36540 11060 36542
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4172 34972 4228 35028
rect 5628 34914 5684 34916
rect 5628 34862 5630 34914
rect 5630 34862 5682 34914
rect 5682 34862 5684 34914
rect 5628 34860 5684 34862
rect 4060 34636 4116 34692
rect 4620 34636 4676 34692
rect 5516 34636 5572 34692
rect 4956 34578 5012 34580
rect 4956 34526 4958 34578
rect 4958 34526 5010 34578
rect 5010 34526 5012 34578
rect 4956 34524 5012 34526
rect 9772 36428 9828 36484
rect 5852 34636 5908 34692
rect 8540 34690 8596 34692
rect 8540 34638 8542 34690
rect 8542 34638 8594 34690
rect 8594 34638 8596 34690
rect 8540 34636 8596 34638
rect 9324 34636 9380 34692
rect 5740 34578 5796 34580
rect 5740 34526 5742 34578
rect 5742 34526 5794 34578
rect 5794 34526 5796 34578
rect 5740 34524 5796 34526
rect 8988 34578 9044 34580
rect 8988 34526 8990 34578
rect 8990 34526 9042 34578
rect 9042 34526 9044 34578
rect 8988 34524 9044 34526
rect 9884 34690 9940 34692
rect 9884 34638 9886 34690
rect 9886 34638 9938 34690
rect 9938 34638 9940 34690
rect 9884 34636 9940 34638
rect 4284 33628 4340 33684
rect 2716 33068 2772 33124
rect 3276 33068 3332 33124
rect 2380 30828 2436 30884
rect 2716 30828 2772 30884
rect 1820 30044 1876 30100
rect 1932 29708 1988 29764
rect 4476 33290 4532 33292
rect 4476 33238 4478 33290
rect 4478 33238 4530 33290
rect 4530 33238 4532 33290
rect 4476 33236 4532 33238
rect 4580 33290 4636 33292
rect 4580 33238 4582 33290
rect 4582 33238 4634 33290
rect 4634 33238 4636 33290
rect 4580 33236 4636 33238
rect 4684 33290 4740 33292
rect 4684 33238 4686 33290
rect 4686 33238 4738 33290
rect 4738 33238 4740 33290
rect 4684 33236 4740 33238
rect 4844 33122 4900 33124
rect 4844 33070 4846 33122
rect 4846 33070 4898 33122
rect 4898 33070 4900 33122
rect 4844 33068 4900 33070
rect 3388 32732 3444 32788
rect 4396 32732 4452 32788
rect 5852 33682 5908 33684
rect 5852 33630 5854 33682
rect 5854 33630 5906 33682
rect 5906 33630 5908 33682
rect 5852 33628 5908 33630
rect 4956 31836 5012 31892
rect 4476 31274 4532 31276
rect 4476 31222 4478 31274
rect 4478 31222 4530 31274
rect 4530 31222 4532 31274
rect 4476 31220 4532 31222
rect 4580 31274 4636 31276
rect 4580 31222 4582 31274
rect 4582 31222 4634 31274
rect 4634 31222 4636 31274
rect 4580 31220 4636 31222
rect 4684 31274 4740 31276
rect 4684 31222 4686 31274
rect 4686 31222 4738 31274
rect 4738 31222 4740 31274
rect 4684 31220 4740 31222
rect 4732 30268 4788 30324
rect 4956 30546 5012 30548
rect 4956 30494 4958 30546
rect 4958 30494 5010 30546
rect 5010 30494 5012 30546
rect 4956 30492 5012 30494
rect 3836 30098 3892 30100
rect 3836 30046 3838 30098
rect 3838 30046 3890 30098
rect 3890 30046 3892 30098
rect 3836 30044 3892 30046
rect 1820 27858 1876 27860
rect 1820 27806 1822 27858
rect 1822 27806 1874 27858
rect 1874 27806 1876 27858
rect 1820 27804 1876 27806
rect 2380 27804 2436 27860
rect 3724 29762 3780 29764
rect 3724 29710 3726 29762
rect 3726 29710 3778 29762
rect 3778 29710 3780 29762
rect 3724 29708 3780 29710
rect 3388 29484 3444 29540
rect 3276 29426 3332 29428
rect 3276 29374 3278 29426
rect 3278 29374 3330 29426
rect 3330 29374 3332 29426
rect 3276 29372 3332 29374
rect 5852 31890 5908 31892
rect 5852 31838 5854 31890
rect 5854 31838 5906 31890
rect 5906 31838 5908 31890
rect 5852 31836 5908 31838
rect 5628 30882 5684 30884
rect 5628 30830 5630 30882
rect 5630 30830 5682 30882
rect 5682 30830 5684 30882
rect 5628 30828 5684 30830
rect 5740 30546 5796 30548
rect 5740 30494 5742 30546
rect 5742 30494 5794 30546
rect 5794 30494 5796 30546
rect 5740 30492 5796 30494
rect 10108 34578 10164 34580
rect 10108 34526 10110 34578
rect 10110 34526 10162 34578
rect 10162 34526 10164 34578
rect 10108 34524 10164 34526
rect 9436 34466 9492 34468
rect 9436 34414 9438 34466
rect 9438 34414 9490 34466
rect 9490 34414 9492 34466
rect 9436 34412 9492 34414
rect 10332 34412 10388 34468
rect 17948 40850 18004 40852
rect 17948 40798 17950 40850
rect 17950 40798 18002 40850
rect 18002 40798 18004 40850
rect 17948 40796 18004 40798
rect 16492 39730 16548 39732
rect 16492 39678 16494 39730
rect 16494 39678 16546 39730
rect 16546 39678 16548 39730
rect 16492 39676 16548 39678
rect 19852 42476 19908 42532
rect 21420 42642 21476 42644
rect 21420 42590 21422 42642
rect 21422 42590 21474 42642
rect 21474 42590 21476 42642
rect 21420 42588 21476 42590
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 23436 44882 23492 44884
rect 23436 44830 23438 44882
rect 23438 44830 23490 44882
rect 23490 44830 23492 44882
rect 23436 44828 23492 44830
rect 22540 43708 22596 43764
rect 22540 43484 22596 43540
rect 22316 42754 22372 42756
rect 22316 42702 22318 42754
rect 22318 42702 22370 42754
rect 22370 42702 22372 42754
rect 22316 42700 22372 42702
rect 23996 44044 24052 44100
rect 24668 44044 24724 44100
rect 23884 43708 23940 43764
rect 23100 43596 23156 43652
rect 22204 42588 22260 42644
rect 26572 47740 26628 47796
rect 26572 47068 26628 47124
rect 27580 46956 27636 47012
rect 26460 45778 26516 45780
rect 26460 45726 26462 45778
rect 26462 45726 26514 45778
rect 26514 45726 26516 45778
rect 26460 45724 26516 45726
rect 26348 44882 26404 44884
rect 26348 44830 26350 44882
rect 26350 44830 26402 44882
rect 26402 44830 26404 44882
rect 26348 44828 26404 44830
rect 27580 45948 27636 46004
rect 27804 46620 27860 46676
rect 27804 44828 27860 44884
rect 28140 44828 28196 44884
rect 27244 44098 27300 44100
rect 27244 44046 27246 44098
rect 27246 44046 27298 44098
rect 27298 44046 27300 44098
rect 27244 44044 27300 44046
rect 26684 43708 26740 43764
rect 27692 43986 27748 43988
rect 27692 43934 27694 43986
rect 27694 43934 27746 43986
rect 27746 43934 27748 43986
rect 27692 43932 27748 43934
rect 24668 43596 24724 43652
rect 23884 43484 23940 43540
rect 23100 42700 23156 42756
rect 23436 42754 23492 42756
rect 23436 42702 23438 42754
rect 23438 42702 23490 42754
rect 23490 42702 23492 42754
rect 23436 42700 23492 42702
rect 22764 42588 22820 42644
rect 21420 42028 21476 42084
rect 18508 41916 18564 41972
rect 20524 41970 20580 41972
rect 20524 41918 20526 41970
rect 20526 41918 20578 41970
rect 20578 41918 20580 41970
rect 20524 41916 20580 41918
rect 21980 41916 22036 41972
rect 21308 41074 21364 41076
rect 21308 41022 21310 41074
rect 21310 41022 21362 41074
rect 21362 41022 21364 41074
rect 21308 41020 21364 41022
rect 18172 40796 18228 40852
rect 18956 40796 19012 40852
rect 18396 39676 18452 39732
rect 17388 39004 17444 39060
rect 18732 39004 18788 39060
rect 16828 38556 16884 38612
rect 13580 36876 13636 36932
rect 17052 37996 17108 38052
rect 17836 38722 17892 38724
rect 17836 38670 17838 38722
rect 17838 38670 17890 38722
rect 17890 38670 17892 38722
rect 17836 38668 17892 38670
rect 18508 38722 18564 38724
rect 18508 38670 18510 38722
rect 18510 38670 18562 38722
rect 18562 38670 18564 38722
rect 18508 38668 18564 38670
rect 17948 38050 18004 38052
rect 17948 37998 17950 38050
rect 17950 37998 18002 38050
rect 18002 37998 18004 38050
rect 17948 37996 18004 37998
rect 17500 37884 17556 37940
rect 18396 37826 18452 37828
rect 18396 37774 18398 37826
rect 18398 37774 18450 37826
rect 18450 37774 18452 37826
rect 18396 37772 18452 37774
rect 16828 37714 16884 37716
rect 16828 37662 16830 37714
rect 16830 37662 16882 37714
rect 16882 37662 16884 37714
rect 16828 37660 16884 37662
rect 14700 36764 14756 36820
rect 14812 36876 14868 36932
rect 13468 36482 13524 36484
rect 13468 36430 13470 36482
rect 13470 36430 13522 36482
rect 13522 36430 13524 36482
rect 13468 36428 13524 36430
rect 12124 35922 12180 35924
rect 12124 35870 12126 35922
rect 12126 35870 12178 35922
rect 12178 35870 12180 35922
rect 12124 35868 12180 35870
rect 15036 36818 15092 36820
rect 15036 36766 15038 36818
rect 15038 36766 15090 36818
rect 15090 36766 15092 36818
rect 15036 36764 15092 36766
rect 15484 36764 15540 36820
rect 14476 35922 14532 35924
rect 14476 35870 14478 35922
rect 14478 35870 14530 35922
rect 14530 35870 14532 35922
rect 14476 35868 14532 35870
rect 14588 35810 14644 35812
rect 14588 35758 14590 35810
rect 14590 35758 14642 35810
rect 14642 35758 14644 35810
rect 14588 35756 14644 35758
rect 12124 34690 12180 34692
rect 12124 34638 12126 34690
rect 12126 34638 12178 34690
rect 12178 34638 12180 34690
rect 12124 34636 12180 34638
rect 13468 34636 13524 34692
rect 10892 34076 10948 34132
rect 11900 34412 11956 34468
rect 11004 33516 11060 33572
rect 12908 34466 12964 34468
rect 12908 34414 12910 34466
rect 12910 34414 12962 34466
rect 12962 34414 12964 34466
rect 12908 34412 12964 34414
rect 12572 34300 12628 34356
rect 12124 34130 12180 34132
rect 12124 34078 12126 34130
rect 12126 34078 12178 34130
rect 12178 34078 12180 34130
rect 12124 34076 12180 34078
rect 13020 34076 13076 34132
rect 13580 33906 13636 33908
rect 13580 33854 13582 33906
rect 13582 33854 13634 33906
rect 13634 33854 13636 33906
rect 13580 33852 13636 33854
rect 15036 34018 15092 34020
rect 15036 33966 15038 34018
rect 15038 33966 15090 34018
rect 15090 33966 15092 34018
rect 15036 33964 15092 33966
rect 12908 33628 12964 33684
rect 12460 33516 12516 33572
rect 14476 33794 14532 33796
rect 14476 33742 14478 33794
rect 14478 33742 14530 33794
rect 14530 33742 14532 33794
rect 14476 33740 14532 33742
rect 14364 33682 14420 33684
rect 14364 33630 14366 33682
rect 14366 33630 14418 33682
rect 14418 33630 14420 33682
rect 14364 33628 14420 33630
rect 14700 33010 14756 33012
rect 14700 32958 14702 33010
rect 14702 32958 14754 33010
rect 14754 32958 14756 33010
rect 14700 32956 14756 32958
rect 14588 32732 14644 32788
rect 12796 32508 12852 32564
rect 10780 32396 10836 32452
rect 11788 32450 11844 32452
rect 11788 32398 11790 32450
rect 11790 32398 11842 32450
rect 11842 32398 11844 32450
rect 11788 32396 11844 32398
rect 11340 31836 11396 31892
rect 9324 30546 9380 30548
rect 9324 30494 9326 30546
rect 9326 30494 9378 30546
rect 9378 30494 9380 30546
rect 9324 30492 9380 30494
rect 6076 30268 6132 30324
rect 3836 28924 3892 28980
rect 5068 29372 5124 29428
rect 4476 29258 4532 29260
rect 4476 29206 4478 29258
rect 4478 29206 4530 29258
rect 4530 29206 4532 29258
rect 4476 29204 4532 29206
rect 4580 29258 4636 29260
rect 4580 29206 4582 29258
rect 4582 29206 4634 29258
rect 4634 29206 4636 29258
rect 4580 29204 4636 29206
rect 4684 29258 4740 29260
rect 4684 29206 4686 29258
rect 4686 29206 4738 29258
rect 4738 29206 4740 29258
rect 4684 29204 4740 29206
rect 4284 29036 4340 29092
rect 4508 28924 4564 28980
rect 5068 28754 5124 28756
rect 5068 28702 5070 28754
rect 5070 28702 5122 28754
rect 5122 28702 5124 28754
rect 5068 28700 5124 28702
rect 2940 27804 2996 27860
rect 3388 27858 3444 27860
rect 3388 27806 3390 27858
rect 3390 27806 3442 27858
rect 3442 27806 3444 27858
rect 3388 27804 3444 27806
rect 4284 27804 4340 27860
rect 6188 29820 6244 29876
rect 6748 30380 6804 30436
rect 5516 29036 5572 29092
rect 8540 29986 8596 29988
rect 8540 29934 8542 29986
rect 8542 29934 8594 29986
rect 8594 29934 8596 29986
rect 8540 29932 8596 29934
rect 9660 30044 9716 30100
rect 9324 29932 9380 29988
rect 6748 28924 6804 28980
rect 6972 29820 7028 29876
rect 6188 28754 6244 28756
rect 6188 28702 6190 28754
rect 6190 28702 6242 28754
rect 6242 28702 6244 28754
rect 6188 28700 6244 28702
rect 5068 27804 5124 27860
rect 5740 27804 5796 27860
rect 4476 27242 4532 27244
rect 4476 27190 4478 27242
rect 4478 27190 4530 27242
rect 4530 27190 4532 27242
rect 4476 27188 4532 27190
rect 4580 27242 4636 27244
rect 4580 27190 4582 27242
rect 4582 27190 4634 27242
rect 4634 27190 4636 27242
rect 4580 27188 4636 27190
rect 4684 27242 4740 27244
rect 4684 27190 4686 27242
rect 4686 27190 4738 27242
rect 4738 27190 4740 27242
rect 4684 27188 4740 27190
rect 7308 29820 7364 29876
rect 7868 29372 7924 29428
rect 8764 29484 8820 29540
rect 8876 29426 8932 29428
rect 8876 29374 8878 29426
rect 8878 29374 8930 29426
rect 8930 29374 8932 29426
rect 8876 29372 8932 29374
rect 10444 30492 10500 30548
rect 10332 30098 10388 30100
rect 10332 30046 10334 30098
rect 10334 30046 10386 30098
rect 10386 30046 10388 30098
rect 10332 30044 10388 30046
rect 9996 29762 10052 29764
rect 9996 29710 9998 29762
rect 9998 29710 10050 29762
rect 10050 29710 10052 29762
rect 9996 29708 10052 29710
rect 8988 28588 9044 28644
rect 8428 28530 8484 28532
rect 8428 28478 8430 28530
rect 8430 28478 8482 28530
rect 8482 28478 8484 28530
rect 8428 28476 8484 28478
rect 9660 29036 9716 29092
rect 9100 28476 9156 28532
rect 10108 29372 10164 29428
rect 14364 31890 14420 31892
rect 14364 31838 14366 31890
rect 14366 31838 14418 31890
rect 14418 31838 14420 31890
rect 14364 31836 14420 31838
rect 13916 31778 13972 31780
rect 13916 31726 13918 31778
rect 13918 31726 13970 31778
rect 13970 31726 13972 31778
rect 13916 31724 13972 31726
rect 14476 31778 14532 31780
rect 14476 31726 14478 31778
rect 14478 31726 14530 31778
rect 14530 31726 14532 31778
rect 14476 31724 14532 31726
rect 13468 31276 13524 31332
rect 12460 30546 12516 30548
rect 12460 30494 12462 30546
rect 12462 30494 12514 30546
rect 12514 30494 12516 30546
rect 12460 30492 12516 30494
rect 11340 29036 11396 29092
rect 10444 28924 10500 28980
rect 17836 36652 17892 36708
rect 15820 36594 15876 36596
rect 15820 36542 15822 36594
rect 15822 36542 15874 36594
rect 15874 36542 15876 36594
rect 15820 36540 15876 36542
rect 16604 35420 16660 35476
rect 16156 34860 16212 34916
rect 18508 36706 18564 36708
rect 18508 36654 18510 36706
rect 18510 36654 18562 36706
rect 18562 36654 18564 36706
rect 18508 36652 18564 36654
rect 18060 36594 18116 36596
rect 18060 36542 18062 36594
rect 18062 36542 18114 36594
rect 18114 36542 18116 36594
rect 18060 36540 18116 36542
rect 20188 40796 20244 40852
rect 19836 40346 19892 40348
rect 19836 40294 19838 40346
rect 19838 40294 19890 40346
rect 19890 40294 19892 40346
rect 19836 40292 19892 40294
rect 19940 40346 19996 40348
rect 19940 40294 19942 40346
rect 19942 40294 19994 40346
rect 19994 40294 19996 40346
rect 19940 40292 19996 40294
rect 20044 40346 20100 40348
rect 20044 40294 20046 40346
rect 20046 40294 20098 40346
rect 20098 40294 20100 40346
rect 20044 40292 20100 40294
rect 19964 38834 20020 38836
rect 19964 38782 19966 38834
rect 19966 38782 20018 38834
rect 20018 38782 20020 38834
rect 19964 38780 20020 38782
rect 19836 38330 19892 38332
rect 19836 38278 19838 38330
rect 19838 38278 19890 38330
rect 19890 38278 19892 38330
rect 19836 38276 19892 38278
rect 19940 38330 19996 38332
rect 19940 38278 19942 38330
rect 19942 38278 19994 38330
rect 19994 38278 19996 38330
rect 19940 38276 19996 38278
rect 20044 38330 20100 38332
rect 20044 38278 20046 38330
rect 20046 38278 20098 38330
rect 20098 38278 20100 38330
rect 20044 38276 20100 38278
rect 19068 37996 19124 38052
rect 18844 36988 18900 37044
rect 19404 37826 19460 37828
rect 19404 37774 19406 37826
rect 19406 37774 19458 37826
rect 19458 37774 19460 37826
rect 19404 37772 19460 37774
rect 20748 40850 20804 40852
rect 20748 40798 20750 40850
rect 20750 40798 20802 40850
rect 20802 40798 20804 40850
rect 20748 40796 20804 40798
rect 21420 40460 21476 40516
rect 21644 39788 21700 39844
rect 19964 37826 20020 37828
rect 19964 37774 19966 37826
rect 19966 37774 20018 37826
rect 20018 37774 20020 37826
rect 19964 37772 20020 37774
rect 20412 39004 20468 39060
rect 21644 39058 21700 39060
rect 21644 39006 21646 39058
rect 21646 39006 21698 39058
rect 21698 39006 21700 39058
rect 21644 39004 21700 39006
rect 21868 38780 21924 38836
rect 20412 38556 20468 38612
rect 20412 37938 20468 37940
rect 20412 37886 20414 37938
rect 20414 37886 20466 37938
rect 20466 37886 20468 37938
rect 20412 37884 20468 37886
rect 20636 37772 20692 37828
rect 19964 36988 20020 37044
rect 19068 36764 19124 36820
rect 19180 36930 19236 36932
rect 19180 36878 19182 36930
rect 19182 36878 19234 36930
rect 19234 36878 19236 36930
rect 19180 36876 19236 36878
rect 17948 35474 18004 35476
rect 17948 35422 17950 35474
rect 17950 35422 18002 35474
rect 18002 35422 18004 35474
rect 17948 35420 18004 35422
rect 16156 33964 16212 34020
rect 15932 33794 15988 33796
rect 15932 33742 15934 33794
rect 15934 33742 15986 33794
rect 15986 33742 15988 33794
rect 15932 33740 15988 33742
rect 15708 32844 15764 32900
rect 15372 32786 15428 32788
rect 15372 32734 15374 32786
rect 15374 32734 15426 32786
rect 15426 32734 15428 32786
rect 15372 32732 15428 32734
rect 16044 32284 16100 32340
rect 15372 31778 15428 31780
rect 15372 31726 15374 31778
rect 15374 31726 15426 31778
rect 15426 31726 15428 31778
rect 15372 31724 15428 31726
rect 14924 31666 14980 31668
rect 14924 31614 14926 31666
rect 14926 31614 14978 31666
rect 14978 31614 14980 31666
rect 14924 31612 14980 31614
rect 15932 31052 15988 31108
rect 15036 30994 15092 30996
rect 15036 30942 15038 30994
rect 15038 30942 15090 30994
rect 15090 30942 15092 30994
rect 15036 30940 15092 30942
rect 20412 36988 20468 37044
rect 20076 36876 20132 36932
rect 19836 36314 19892 36316
rect 19836 36262 19838 36314
rect 19838 36262 19890 36314
rect 19890 36262 19892 36314
rect 19836 36260 19892 36262
rect 19940 36314 19996 36316
rect 19940 36262 19942 36314
rect 19942 36262 19994 36314
rect 19994 36262 19996 36314
rect 19940 36260 19996 36262
rect 20044 36314 20100 36316
rect 20044 36262 20046 36314
rect 20046 36262 20098 36314
rect 20098 36262 20100 36314
rect 20044 36260 20100 36262
rect 20076 36092 20132 36148
rect 19740 35922 19796 35924
rect 19740 35870 19742 35922
rect 19742 35870 19794 35922
rect 19794 35870 19796 35922
rect 19740 35868 19796 35870
rect 18956 35308 19012 35364
rect 19180 34972 19236 35028
rect 19628 35810 19684 35812
rect 19628 35758 19630 35810
rect 19630 35758 19682 35810
rect 19682 35758 19684 35810
rect 19628 35756 19684 35758
rect 19516 34860 19572 34916
rect 18396 33794 18452 33796
rect 18396 33742 18398 33794
rect 18398 33742 18450 33794
rect 18450 33742 18452 33794
rect 18396 33740 18452 33742
rect 18396 32732 18452 32788
rect 20524 35308 20580 35364
rect 20300 34972 20356 35028
rect 18956 32844 19012 32900
rect 19292 32956 19348 33012
rect 16380 31724 16436 31780
rect 16828 31276 16884 31332
rect 17948 32562 18004 32564
rect 17948 32510 17950 32562
rect 17950 32510 18002 32562
rect 18002 32510 18004 32562
rect 17948 32508 18004 32510
rect 17836 31500 17892 31556
rect 19180 30828 19236 30884
rect 13468 30492 13524 30548
rect 13916 30604 13972 30660
rect 13580 30434 13636 30436
rect 13580 30382 13582 30434
rect 13582 30382 13634 30434
rect 13634 30382 13636 30434
rect 13580 30380 13636 30382
rect 12908 29708 12964 29764
rect 12796 28978 12852 28980
rect 12796 28926 12798 28978
rect 12798 28926 12850 28978
rect 12850 28926 12852 28978
rect 12796 28924 12852 28926
rect 13468 29090 13524 29092
rect 13468 29038 13470 29090
rect 13470 29038 13522 29090
rect 13522 29038 13524 29090
rect 13468 29036 13524 29038
rect 12908 28700 12964 28756
rect 13916 29596 13972 29652
rect 14588 30492 14644 30548
rect 14252 30156 14308 30212
rect 14028 28924 14084 28980
rect 14476 28754 14532 28756
rect 14476 28702 14478 28754
rect 14478 28702 14530 28754
rect 14530 28702 14532 28754
rect 14476 28700 14532 28702
rect 12796 28588 12852 28644
rect 15484 30658 15540 30660
rect 15484 30606 15486 30658
rect 15486 30606 15538 30658
rect 15538 30606 15540 30658
rect 15484 30604 15540 30606
rect 16044 30380 16100 30436
rect 17724 30492 17780 30548
rect 18284 30380 18340 30436
rect 17724 30044 17780 30100
rect 15260 29874 15316 29876
rect 15260 29822 15262 29874
rect 15262 29822 15314 29874
rect 15314 29822 15316 29874
rect 15260 29820 15316 29822
rect 19836 34298 19892 34300
rect 19836 34246 19838 34298
rect 19838 34246 19890 34298
rect 19890 34246 19892 34298
rect 19836 34244 19892 34246
rect 19940 34298 19996 34300
rect 19940 34246 19942 34298
rect 19942 34246 19994 34298
rect 19994 34246 19996 34298
rect 19940 34244 19996 34246
rect 20044 34298 20100 34300
rect 20044 34246 20046 34298
rect 20046 34246 20098 34298
rect 20098 34246 20100 34298
rect 20044 34244 20100 34246
rect 20524 33628 20580 33684
rect 20412 33010 20468 33012
rect 20412 32958 20414 33010
rect 20414 32958 20466 33010
rect 20466 32958 20468 33010
rect 20412 32956 20468 32958
rect 19836 32282 19892 32284
rect 19836 32230 19838 32282
rect 19838 32230 19890 32282
rect 19890 32230 19892 32282
rect 19836 32228 19892 32230
rect 19940 32282 19996 32284
rect 19940 32230 19942 32282
rect 19942 32230 19994 32282
rect 19994 32230 19996 32282
rect 19940 32228 19996 32230
rect 20044 32282 20100 32284
rect 20044 32230 20046 32282
rect 20046 32230 20098 32282
rect 20098 32230 20100 32282
rect 20044 32228 20100 32230
rect 20188 31836 20244 31892
rect 20188 31276 20244 31332
rect 19180 29820 19236 29876
rect 19836 30266 19892 30268
rect 19836 30214 19838 30266
rect 19838 30214 19890 30266
rect 19890 30214 19892 30266
rect 19836 30212 19892 30214
rect 19940 30266 19996 30268
rect 19940 30214 19942 30266
rect 19942 30214 19994 30266
rect 19994 30214 19996 30266
rect 19940 30212 19996 30214
rect 20044 30266 20100 30268
rect 20044 30214 20046 30266
rect 20046 30214 20098 30266
rect 20098 30214 20100 30266
rect 20044 30212 20100 30214
rect 19628 29820 19684 29876
rect 19628 28812 19684 28868
rect 19516 28700 19572 28756
rect 14700 28588 14756 28644
rect 15036 28642 15092 28644
rect 15036 28590 15038 28642
rect 15038 28590 15090 28642
rect 15090 28590 15092 28642
rect 15036 28588 15092 28590
rect 17836 28588 17892 28644
rect 15932 26738 15988 26740
rect 15932 26686 15934 26738
rect 15934 26686 15986 26738
rect 15986 26686 15988 26738
rect 15932 26684 15988 26686
rect 14588 25788 14644 25844
rect 4476 25226 4532 25228
rect 4476 25174 4478 25226
rect 4478 25174 4530 25226
rect 4530 25174 4532 25226
rect 4476 25172 4532 25174
rect 4580 25226 4636 25228
rect 4580 25174 4582 25226
rect 4582 25174 4634 25226
rect 4634 25174 4636 25226
rect 4580 25172 4636 25174
rect 4684 25226 4740 25228
rect 4684 25174 4686 25226
rect 4686 25174 4738 25226
rect 4738 25174 4740 25226
rect 4684 25172 4740 25174
rect 11676 23714 11732 23716
rect 11676 23662 11678 23714
rect 11678 23662 11730 23714
rect 11730 23662 11732 23714
rect 11676 23660 11732 23662
rect 13468 23660 13524 23716
rect 15148 23660 15204 23716
rect 4476 23210 4532 23212
rect 4476 23158 4478 23210
rect 4478 23158 4530 23210
rect 4530 23158 4532 23210
rect 4476 23156 4532 23158
rect 4580 23210 4636 23212
rect 4580 23158 4582 23210
rect 4582 23158 4634 23210
rect 4634 23158 4636 23210
rect 4580 23156 4636 23158
rect 4684 23210 4740 23212
rect 4684 23158 4686 23210
rect 4686 23158 4738 23210
rect 4738 23158 4740 23210
rect 4684 23156 4740 23158
rect 16716 25954 16772 25956
rect 16716 25902 16718 25954
rect 16718 25902 16770 25954
rect 16770 25902 16772 25954
rect 16716 25900 16772 25902
rect 17052 26626 17108 26628
rect 17052 26574 17054 26626
rect 17054 26574 17106 26626
rect 17106 26574 17108 26626
rect 17052 26572 17108 26574
rect 20300 28754 20356 28756
rect 20300 28702 20302 28754
rect 20302 28702 20354 28754
rect 20354 28702 20356 28754
rect 20300 28700 20356 28702
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 17948 26572 18004 26628
rect 17724 26012 17780 26068
rect 17612 25842 17668 25844
rect 17612 25790 17614 25842
rect 17614 25790 17666 25842
rect 17666 25790 17668 25842
rect 17612 25788 17668 25790
rect 18956 26348 19012 26404
rect 18172 25900 18228 25956
rect 19852 26348 19908 26404
rect 19836 26234 19892 26236
rect 19836 26182 19838 26234
rect 19838 26182 19890 26234
rect 19890 26182 19892 26234
rect 19836 26180 19892 26182
rect 19940 26234 19996 26236
rect 19940 26182 19942 26234
rect 19942 26182 19994 26234
rect 19994 26182 19996 26234
rect 19940 26180 19996 26182
rect 20044 26234 20100 26236
rect 20044 26182 20046 26234
rect 20046 26182 20098 26234
rect 20098 26182 20100 26234
rect 20044 26180 20100 26182
rect 21532 38556 21588 38612
rect 21308 37884 21364 37940
rect 21084 37660 21140 37716
rect 21420 36876 21476 36932
rect 21756 36988 21812 37044
rect 21420 36652 21476 36708
rect 21644 36594 21700 36596
rect 21644 36542 21646 36594
rect 21646 36542 21698 36594
rect 21698 36542 21700 36594
rect 21644 36540 21700 36542
rect 21756 36034 21812 36036
rect 21756 35982 21758 36034
rect 21758 35982 21810 36034
rect 21810 35982 21812 36034
rect 21756 35980 21812 35982
rect 20748 35868 20804 35924
rect 23772 41916 23828 41972
rect 26124 41970 26180 41972
rect 26124 41918 26126 41970
rect 26126 41918 26178 41970
rect 26178 41918 26180 41970
rect 26124 41916 26180 41918
rect 26348 41916 26404 41972
rect 28140 43932 28196 43988
rect 28588 46002 28644 46004
rect 28588 45950 28590 46002
rect 28590 45950 28642 46002
rect 28642 45950 28644 46002
rect 28588 45948 28644 45950
rect 28588 43932 28644 43988
rect 27804 42812 27860 42868
rect 29260 45724 29316 45780
rect 29484 44882 29540 44884
rect 29484 44830 29486 44882
rect 29486 44830 29538 44882
rect 29538 44830 29540 44882
rect 29484 44828 29540 44830
rect 28812 43986 28868 43988
rect 28812 43934 28814 43986
rect 28814 43934 28866 43986
rect 28866 43934 28868 43986
rect 28812 43932 28868 43934
rect 26908 42028 26964 42084
rect 26796 41692 26852 41748
rect 26012 41580 26068 41636
rect 22540 40684 22596 40740
rect 23100 40684 23156 40740
rect 23884 40738 23940 40740
rect 23884 40686 23886 40738
rect 23886 40686 23938 40738
rect 23938 40686 23940 40738
rect 23884 40684 23940 40686
rect 22652 39842 22708 39844
rect 22652 39790 22654 39842
rect 22654 39790 22706 39842
rect 22706 39790 22708 39842
rect 22652 39788 22708 39790
rect 22092 37938 22148 37940
rect 22092 37886 22094 37938
rect 22094 37886 22146 37938
rect 22146 37886 22148 37938
rect 22092 37884 22148 37886
rect 22204 37660 22260 37716
rect 24668 40066 24724 40068
rect 24668 40014 24670 40066
rect 24670 40014 24722 40066
rect 24722 40014 24724 40066
rect 24668 40012 24724 40014
rect 25116 40572 25172 40628
rect 24220 39900 24276 39956
rect 25116 39954 25172 39956
rect 25116 39902 25118 39954
rect 25118 39902 25170 39954
rect 25170 39902 25172 39954
rect 25116 39900 25172 39902
rect 25452 40012 25508 40068
rect 26572 40348 26628 40404
rect 22988 38668 23044 38724
rect 26460 39788 26516 39844
rect 22652 37660 22708 37716
rect 21980 36876 22036 36932
rect 21980 36706 22036 36708
rect 21980 36654 21982 36706
rect 21982 36654 22034 36706
rect 22034 36654 22036 36706
rect 21980 36652 22036 36654
rect 22204 36706 22260 36708
rect 22204 36654 22206 36706
rect 22206 36654 22258 36706
rect 22258 36654 22260 36706
rect 22204 36652 22260 36654
rect 21980 36034 22036 36036
rect 21980 35982 21982 36034
rect 21982 35982 22034 36034
rect 22034 35982 22036 36034
rect 21980 35980 22036 35982
rect 23548 37938 23604 37940
rect 23548 37886 23550 37938
rect 23550 37886 23602 37938
rect 23602 37886 23604 37938
rect 23548 37884 23604 37886
rect 22540 36652 22596 36708
rect 22540 35698 22596 35700
rect 22540 35646 22542 35698
rect 22542 35646 22594 35698
rect 22594 35646 22596 35698
rect 22540 35644 22596 35646
rect 22876 36092 22932 36148
rect 25116 38780 25172 38836
rect 26012 38220 26068 38276
rect 24892 37660 24948 37716
rect 23548 36540 23604 36596
rect 23100 35644 23156 35700
rect 23212 35756 23268 35812
rect 22540 34972 22596 35028
rect 22540 34802 22596 34804
rect 22540 34750 22542 34802
rect 22542 34750 22594 34802
rect 22594 34750 22596 34802
rect 22540 34748 22596 34750
rect 22428 34636 22484 34692
rect 21532 33682 21588 33684
rect 21532 33630 21534 33682
rect 21534 33630 21586 33682
rect 21586 33630 21588 33682
rect 21532 33628 21588 33630
rect 21980 33628 22036 33684
rect 21084 32956 21140 33012
rect 20972 31890 21028 31892
rect 20972 31838 20974 31890
rect 20974 31838 21026 31890
rect 21026 31838 21028 31890
rect 20972 31836 21028 31838
rect 21868 31890 21924 31892
rect 21868 31838 21870 31890
rect 21870 31838 21922 31890
rect 21922 31838 21924 31890
rect 21868 31836 21924 31838
rect 20748 31500 20804 31556
rect 20860 31778 20916 31780
rect 20860 31726 20862 31778
rect 20862 31726 20914 31778
rect 20914 31726 20916 31778
rect 20860 31724 20916 31726
rect 21420 31724 21476 31780
rect 21756 31500 21812 31556
rect 20860 31388 20916 31444
rect 21308 28754 21364 28756
rect 21308 28702 21310 28754
rect 21310 28702 21362 28754
rect 21362 28702 21364 28754
rect 21308 28700 21364 28702
rect 20748 28642 20804 28644
rect 20748 28590 20750 28642
rect 20750 28590 20802 28642
rect 20802 28590 20804 28642
rect 20748 28588 20804 28590
rect 21756 28588 21812 28644
rect 20860 27746 20916 27748
rect 20860 27694 20862 27746
rect 20862 27694 20914 27746
rect 20914 27694 20916 27746
rect 20860 27692 20916 27694
rect 21644 27356 21700 27412
rect 21868 26572 21924 26628
rect 20748 26514 20804 26516
rect 20748 26462 20750 26514
rect 20750 26462 20802 26514
rect 20802 26462 20804 26514
rect 20748 26460 20804 26462
rect 18620 25394 18676 25396
rect 18620 25342 18622 25394
rect 18622 25342 18674 25394
rect 18674 25342 18676 25394
rect 18620 25340 18676 25342
rect 20972 26348 21028 26404
rect 17500 23714 17556 23716
rect 17500 23662 17502 23714
rect 17502 23662 17554 23714
rect 17554 23662 17556 23714
rect 17500 23660 17556 23662
rect 19404 24780 19460 24836
rect 19180 23826 19236 23828
rect 19180 23774 19182 23826
rect 19182 23774 19234 23826
rect 19234 23774 19236 23826
rect 19180 23772 19236 23774
rect 18844 23714 18900 23716
rect 18844 23662 18846 23714
rect 18846 23662 18898 23714
rect 18898 23662 18900 23714
rect 18844 23660 18900 23662
rect 20188 24556 20244 24612
rect 19836 24218 19892 24220
rect 19836 24166 19838 24218
rect 19838 24166 19890 24218
rect 19890 24166 19892 24218
rect 19836 24164 19892 24166
rect 19940 24218 19996 24220
rect 19940 24166 19942 24218
rect 19942 24166 19994 24218
rect 19994 24166 19996 24218
rect 19940 24164 19996 24166
rect 20044 24218 20100 24220
rect 20044 24166 20046 24218
rect 20046 24166 20098 24218
rect 20098 24166 20100 24218
rect 20044 24164 20100 24166
rect 21420 26012 21476 26068
rect 21868 26012 21924 26068
rect 21420 25676 21476 25732
rect 24220 36540 24276 36596
rect 24108 35810 24164 35812
rect 24108 35758 24110 35810
rect 24110 35758 24162 35810
rect 24162 35758 24164 35810
rect 24108 35756 24164 35758
rect 24780 36034 24836 36036
rect 24780 35982 24782 36034
rect 24782 35982 24834 36034
rect 24834 35982 24836 36034
rect 24780 35980 24836 35982
rect 23772 35644 23828 35700
rect 23548 34802 23604 34804
rect 23548 34750 23550 34802
rect 23550 34750 23602 34802
rect 23602 34750 23604 34802
rect 23548 34748 23604 34750
rect 23772 34690 23828 34692
rect 23772 34638 23774 34690
rect 23774 34638 23826 34690
rect 23826 34638 23828 34690
rect 23772 34636 23828 34638
rect 22428 33628 22484 33684
rect 22764 33628 22820 33684
rect 23212 34524 23268 34580
rect 23212 33740 23268 33796
rect 22764 31612 22820 31668
rect 22876 31500 22932 31556
rect 23884 32284 23940 32340
rect 23212 31778 23268 31780
rect 23212 31726 23214 31778
rect 23214 31726 23266 31778
rect 23266 31726 23268 31778
rect 23212 31724 23268 31726
rect 24444 35756 24500 35812
rect 24668 33682 24724 33684
rect 24668 33630 24670 33682
rect 24670 33630 24722 33682
rect 24722 33630 24724 33682
rect 24668 33628 24724 33630
rect 24220 31948 24276 32004
rect 24108 31890 24164 31892
rect 24108 31838 24110 31890
rect 24110 31838 24162 31890
rect 24162 31838 24164 31890
rect 24108 31836 24164 31838
rect 24108 31500 24164 31556
rect 23772 31388 23828 31444
rect 22652 30492 22708 30548
rect 22316 28754 22372 28756
rect 22316 28702 22318 28754
rect 22318 28702 22370 28754
rect 22370 28702 22372 28754
rect 22316 28700 22372 28702
rect 23100 29932 23156 29988
rect 22988 28700 23044 28756
rect 22204 27746 22260 27748
rect 22204 27694 22206 27746
rect 22206 27694 22258 27746
rect 22258 27694 22260 27746
rect 22204 27692 22260 27694
rect 22092 26460 22148 26516
rect 21644 24834 21700 24836
rect 21644 24782 21646 24834
rect 21646 24782 21698 24834
rect 21698 24782 21700 24834
rect 21644 24780 21700 24782
rect 22092 24834 22148 24836
rect 22092 24782 22094 24834
rect 22094 24782 22146 24834
rect 22146 24782 22148 24834
rect 22092 24780 22148 24782
rect 21084 24668 21140 24724
rect 20300 24332 20356 24388
rect 20748 23884 20804 23940
rect 22540 26850 22596 26852
rect 22540 26798 22542 26850
rect 22542 26798 22594 26850
rect 22594 26798 22596 26850
rect 22540 26796 22596 26798
rect 23660 27692 23716 27748
rect 22876 27410 22932 27412
rect 22876 27358 22878 27410
rect 22878 27358 22930 27410
rect 22930 27358 22932 27410
rect 22876 27356 22932 27358
rect 23996 30770 24052 30772
rect 23996 30718 23998 30770
rect 23998 30718 24050 30770
rect 24050 30718 24052 30770
rect 23996 30716 24052 30718
rect 24332 29986 24388 29988
rect 24332 29934 24334 29986
rect 24334 29934 24386 29986
rect 24386 29934 24388 29986
rect 24332 29932 24388 29934
rect 23884 29484 23940 29540
rect 24556 29932 24612 29988
rect 24780 32284 24836 32340
rect 25788 37938 25844 37940
rect 25788 37886 25790 37938
rect 25790 37886 25842 37938
rect 25842 37886 25844 37938
rect 25788 37884 25844 37886
rect 25340 36652 25396 36708
rect 25116 36540 25172 36596
rect 25228 33628 25284 33684
rect 25340 31948 25396 32004
rect 25228 31612 25284 31668
rect 25004 31500 25060 31556
rect 24444 29820 24500 29876
rect 24332 29708 24388 29764
rect 24220 29148 24276 29204
rect 24220 28924 24276 28980
rect 25116 31106 25172 31108
rect 25116 31054 25118 31106
rect 25118 31054 25170 31106
rect 25170 31054 25172 31106
rect 25116 31052 25172 31054
rect 25004 30658 25060 30660
rect 25004 30606 25006 30658
rect 25006 30606 25058 30658
rect 25058 30606 25060 30658
rect 25004 30604 25060 30606
rect 25004 29708 25060 29764
rect 25228 29484 25284 29540
rect 25004 28924 25060 28980
rect 25116 28754 25172 28756
rect 25116 28702 25118 28754
rect 25118 28702 25170 28754
rect 25170 28702 25172 28754
rect 25116 28700 25172 28702
rect 24444 27746 24500 27748
rect 24444 27694 24446 27746
rect 24446 27694 24498 27746
rect 24498 27694 24500 27746
rect 24444 27692 24500 27694
rect 22204 24668 22260 24724
rect 21756 24444 21812 24500
rect 21532 23884 21588 23940
rect 19836 22202 19892 22204
rect 19836 22150 19838 22202
rect 19838 22150 19890 22202
rect 19890 22150 19892 22202
rect 19836 22148 19892 22150
rect 19940 22202 19996 22204
rect 19940 22150 19942 22202
rect 19942 22150 19994 22202
rect 19994 22150 19996 22202
rect 19940 22148 19996 22150
rect 20044 22202 20100 22204
rect 20044 22150 20046 22202
rect 20046 22150 20098 22202
rect 20098 22150 20100 22202
rect 20044 22148 20100 22150
rect 19852 21698 19908 21700
rect 19852 21646 19854 21698
rect 19854 21646 19906 21698
rect 19906 21646 19908 21698
rect 19852 21644 19908 21646
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 18508 20690 18564 20692
rect 18508 20638 18510 20690
rect 18510 20638 18562 20690
rect 18562 20638 18564 20690
rect 18508 20636 18564 20638
rect 4476 19178 4532 19180
rect 4476 19126 4478 19178
rect 4478 19126 4530 19178
rect 4530 19126 4532 19178
rect 4476 19124 4532 19126
rect 4580 19178 4636 19180
rect 4580 19126 4582 19178
rect 4582 19126 4634 19178
rect 4634 19126 4636 19178
rect 4580 19124 4636 19126
rect 4684 19178 4740 19180
rect 4684 19126 4686 19178
rect 4686 19126 4738 19178
rect 4738 19126 4740 19178
rect 4684 19124 4740 19126
rect 17500 18674 17556 18676
rect 17500 18622 17502 18674
rect 17502 18622 17554 18674
rect 17554 18622 17556 18674
rect 17500 18620 17556 18622
rect 16604 18562 16660 18564
rect 16604 18510 16606 18562
rect 16606 18510 16658 18562
rect 16658 18510 16660 18562
rect 16604 18508 16660 18510
rect 18396 19068 18452 19124
rect 18284 18674 18340 18676
rect 18284 18622 18286 18674
rect 18286 18622 18338 18674
rect 18338 18622 18340 18674
rect 18284 18620 18340 18622
rect 17724 18562 17780 18564
rect 17724 18510 17726 18562
rect 17726 18510 17778 18562
rect 17778 18510 17780 18562
rect 17724 18508 17780 18510
rect 16828 17554 16884 17556
rect 16828 17502 16830 17554
rect 16830 17502 16882 17554
rect 16882 17502 16884 17554
rect 16828 17500 16884 17502
rect 19292 20524 19348 20580
rect 19740 20466 19796 20468
rect 19740 20414 19742 20466
rect 19742 20414 19794 20466
rect 19794 20414 19796 20466
rect 19740 20412 19796 20414
rect 19852 20300 19908 20356
rect 20300 21868 20356 21924
rect 21868 23772 21924 23828
rect 22428 25730 22484 25732
rect 22428 25678 22430 25730
rect 22430 25678 22482 25730
rect 22482 25678 22484 25730
rect 22428 25676 22484 25678
rect 22540 26236 22596 26292
rect 22764 26066 22820 26068
rect 22764 26014 22766 26066
rect 22766 26014 22818 26066
rect 22818 26014 22820 26066
rect 22764 26012 22820 26014
rect 23548 26626 23604 26628
rect 23548 26574 23550 26626
rect 23550 26574 23602 26626
rect 23602 26574 23604 26626
rect 23548 26572 23604 26574
rect 23324 26514 23380 26516
rect 23324 26462 23326 26514
rect 23326 26462 23378 26514
rect 23378 26462 23380 26514
rect 23324 26460 23380 26462
rect 23772 26460 23828 26516
rect 23212 26348 23268 26404
rect 22316 24556 22372 24612
rect 22316 23772 22372 23828
rect 19836 20186 19892 20188
rect 19836 20134 19838 20186
rect 19838 20134 19890 20186
rect 19890 20134 19892 20186
rect 19836 20132 19892 20134
rect 19940 20186 19996 20188
rect 19940 20134 19942 20186
rect 19942 20134 19994 20186
rect 19994 20134 19996 20186
rect 19940 20132 19996 20134
rect 20044 20186 20100 20188
rect 20044 20134 20046 20186
rect 20046 20134 20098 20186
rect 20098 20134 20100 20186
rect 20044 20132 20100 20134
rect 20300 20636 20356 20692
rect 20748 20188 20804 20244
rect 20636 20076 20692 20132
rect 20188 19740 20244 19796
rect 21084 19794 21140 19796
rect 21084 19742 21086 19794
rect 21086 19742 21138 19794
rect 21138 19742 21140 19794
rect 21084 19740 21140 19742
rect 19516 19068 19572 19124
rect 18508 18508 18564 18564
rect 18956 18508 19012 18564
rect 18284 18396 18340 18452
rect 19180 18450 19236 18452
rect 19180 18398 19182 18450
rect 19182 18398 19234 18450
rect 19234 18398 19236 18450
rect 19180 18396 19236 18398
rect 20188 19068 20244 19124
rect 20300 18956 20356 19012
rect 19740 18674 19796 18676
rect 19740 18622 19742 18674
rect 19742 18622 19794 18674
rect 19794 18622 19796 18674
rect 19740 18620 19796 18622
rect 19836 18170 19892 18172
rect 19836 18118 19838 18170
rect 19838 18118 19890 18170
rect 19890 18118 19892 18170
rect 19836 18116 19892 18118
rect 19940 18170 19996 18172
rect 19940 18118 19942 18170
rect 19942 18118 19994 18170
rect 19994 18118 19996 18170
rect 19940 18116 19996 18118
rect 20044 18170 20100 18172
rect 20044 18118 20046 18170
rect 20046 18118 20098 18170
rect 20098 18118 20100 18170
rect 20044 18116 20100 18118
rect 4476 17162 4532 17164
rect 4476 17110 4478 17162
rect 4478 17110 4530 17162
rect 4530 17110 4532 17162
rect 4476 17108 4532 17110
rect 4580 17162 4636 17164
rect 4580 17110 4582 17162
rect 4582 17110 4634 17162
rect 4634 17110 4636 17162
rect 4580 17108 4636 17110
rect 4684 17162 4740 17164
rect 4684 17110 4686 17162
rect 4686 17110 4738 17162
rect 4738 17110 4740 17162
rect 4684 17108 4740 17110
rect 15036 16658 15092 16660
rect 15036 16606 15038 16658
rect 15038 16606 15090 16658
rect 15090 16606 15092 16658
rect 15036 16604 15092 16606
rect 17612 16604 17668 16660
rect 18284 17500 18340 17556
rect 4476 15146 4532 15148
rect 4476 15094 4478 15146
rect 4478 15094 4530 15146
rect 4530 15094 4532 15146
rect 4476 15092 4532 15094
rect 4580 15146 4636 15148
rect 4580 15094 4582 15146
rect 4582 15094 4634 15146
rect 4634 15094 4636 15146
rect 4580 15092 4636 15094
rect 4684 15146 4740 15148
rect 4684 15094 4686 15146
rect 4686 15094 4738 15146
rect 4738 15094 4740 15146
rect 4684 15092 4740 15094
rect 17612 13468 17668 13524
rect 4476 13130 4532 13132
rect 4476 13078 4478 13130
rect 4478 13078 4530 13130
rect 4530 13078 4532 13130
rect 4476 13076 4532 13078
rect 4580 13130 4636 13132
rect 4580 13078 4582 13130
rect 4582 13078 4634 13130
rect 4634 13078 4636 13130
rect 4580 13076 4636 13078
rect 4684 13130 4740 13132
rect 4684 13078 4686 13130
rect 4686 13078 4738 13130
rect 4738 13078 4740 13130
rect 4684 13076 4740 13078
rect 18732 17554 18788 17556
rect 18732 17502 18734 17554
rect 18734 17502 18786 17554
rect 18786 17502 18788 17554
rect 18732 17500 18788 17502
rect 21532 20578 21588 20580
rect 21532 20526 21534 20578
rect 21534 20526 21586 20578
rect 21586 20526 21588 20578
rect 21532 20524 21588 20526
rect 21420 18956 21476 19012
rect 22092 20578 22148 20580
rect 22092 20526 22094 20578
rect 22094 20526 22146 20578
rect 22146 20526 22148 20578
rect 22092 20524 22148 20526
rect 22876 24498 22932 24500
rect 22876 24446 22878 24498
rect 22878 24446 22930 24498
rect 22930 24446 22932 24498
rect 22876 24444 22932 24446
rect 22652 24332 22708 24388
rect 22540 23884 22596 23940
rect 23436 25842 23492 25844
rect 23436 25790 23438 25842
rect 23438 25790 23490 25842
rect 23490 25790 23492 25842
rect 23436 25788 23492 25790
rect 23324 24722 23380 24724
rect 23324 24670 23326 24722
rect 23326 24670 23378 24722
rect 23378 24670 23380 24722
rect 23324 24668 23380 24670
rect 23548 24332 23604 24388
rect 23100 23826 23156 23828
rect 23100 23774 23102 23826
rect 23102 23774 23154 23826
rect 23154 23774 23156 23826
rect 23100 23772 23156 23774
rect 23548 23884 23604 23940
rect 23660 23660 23716 23716
rect 23212 23548 23268 23604
rect 23884 24610 23940 24612
rect 23884 24558 23886 24610
rect 23886 24558 23938 24610
rect 23938 24558 23940 24610
rect 23884 24556 23940 24558
rect 25004 28530 25060 28532
rect 25004 28478 25006 28530
rect 25006 28478 25058 28530
rect 25058 28478 25060 28530
rect 25004 28476 25060 28478
rect 25564 35922 25620 35924
rect 25564 35870 25566 35922
rect 25566 35870 25618 35922
rect 25618 35870 25620 35922
rect 25564 35868 25620 35870
rect 26348 37714 26404 37716
rect 26348 37662 26350 37714
rect 26350 37662 26402 37714
rect 26402 37662 26404 37714
rect 26348 37660 26404 37662
rect 25900 35810 25956 35812
rect 25900 35758 25902 35810
rect 25902 35758 25954 35810
rect 25954 35758 25956 35810
rect 25900 35756 25956 35758
rect 25900 34578 25956 34580
rect 25900 34526 25902 34578
rect 25902 34526 25954 34578
rect 25954 34526 25956 34578
rect 25900 34524 25956 34526
rect 26796 34018 26852 34020
rect 26796 33966 26798 34018
rect 26798 33966 26850 34018
rect 26850 33966 26852 34018
rect 26796 33964 26852 33966
rect 25788 33292 25844 33348
rect 26460 33852 26516 33908
rect 26124 32844 26180 32900
rect 25788 30828 25844 30884
rect 26012 31724 26068 31780
rect 26460 31836 26516 31892
rect 26348 31500 26404 31556
rect 26236 30828 26292 30884
rect 25900 30716 25956 30772
rect 25564 30658 25620 30660
rect 25564 30606 25566 30658
rect 25566 30606 25618 30658
rect 25618 30606 25620 30658
rect 25564 30604 25620 30606
rect 26348 30658 26404 30660
rect 26348 30606 26350 30658
rect 26350 30606 26402 30658
rect 26402 30606 26404 30658
rect 26348 30604 26404 30606
rect 26012 30268 26068 30324
rect 26460 30380 26516 30436
rect 25788 30156 25844 30212
rect 25564 30098 25620 30100
rect 25564 30046 25566 30098
rect 25566 30046 25618 30098
rect 25618 30046 25620 30098
rect 25564 30044 25620 30046
rect 27132 41970 27188 41972
rect 27132 41918 27134 41970
rect 27134 41918 27186 41970
rect 27186 41918 27188 41970
rect 27132 41916 27188 41918
rect 28028 42588 28084 42644
rect 28028 42028 28084 42084
rect 27020 41580 27076 41636
rect 27020 40348 27076 40404
rect 27132 40012 27188 40068
rect 27692 39900 27748 39956
rect 27580 39788 27636 39844
rect 27132 39228 27188 39284
rect 27580 38834 27636 38836
rect 27580 38782 27582 38834
rect 27582 38782 27634 38834
rect 27634 38782 27636 38834
rect 27580 38780 27636 38782
rect 27244 37660 27300 37716
rect 27356 36652 27412 36708
rect 27356 36092 27412 36148
rect 27020 35922 27076 35924
rect 27020 35870 27022 35922
rect 27022 35870 27074 35922
rect 27074 35870 27076 35922
rect 27020 35868 27076 35870
rect 27132 35308 27188 35364
rect 27580 33964 27636 34020
rect 27132 33906 27188 33908
rect 27132 33854 27134 33906
rect 27134 33854 27186 33906
rect 27186 33854 27188 33906
rect 27132 33852 27188 33854
rect 27692 33794 27748 33796
rect 27692 33742 27694 33794
rect 27694 33742 27746 33794
rect 27746 33742 27748 33794
rect 27692 33740 27748 33742
rect 28588 42812 28644 42868
rect 29484 40796 29540 40852
rect 29372 40626 29428 40628
rect 29372 40574 29374 40626
rect 29374 40574 29426 40626
rect 29426 40574 29428 40626
rect 29372 40572 29428 40574
rect 29260 40460 29316 40516
rect 28476 40012 28532 40068
rect 29260 39954 29316 39956
rect 29260 39902 29262 39954
rect 29262 39902 29314 39954
rect 29314 39902 29316 39954
rect 29260 39900 29316 39902
rect 28364 39228 28420 39284
rect 28364 38892 28420 38948
rect 28252 38332 28308 38388
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 35196 55466 35252 55468
rect 35196 55414 35198 55466
rect 35198 55414 35250 55466
rect 35250 55414 35252 55466
rect 35196 55412 35252 55414
rect 35300 55466 35356 55468
rect 35300 55414 35302 55466
rect 35302 55414 35354 55466
rect 35354 55414 35356 55466
rect 35300 55412 35356 55414
rect 35404 55466 35460 55468
rect 35404 55414 35406 55466
rect 35406 55414 35458 55466
rect 35458 55414 35460 55466
rect 35404 55412 35460 55414
rect 50556 54458 50612 54460
rect 50556 54406 50558 54458
rect 50558 54406 50610 54458
rect 50610 54406 50612 54458
rect 50556 54404 50612 54406
rect 50660 54458 50716 54460
rect 50660 54406 50662 54458
rect 50662 54406 50714 54458
rect 50714 54406 50716 54458
rect 50660 54404 50716 54406
rect 50764 54458 50820 54460
rect 50764 54406 50766 54458
rect 50766 54406 50818 54458
rect 50818 54406 50820 54458
rect 50764 54404 50820 54406
rect 55244 53788 55300 53844
rect 35196 53450 35252 53452
rect 35196 53398 35198 53450
rect 35198 53398 35250 53450
rect 35250 53398 35252 53450
rect 35196 53396 35252 53398
rect 35300 53450 35356 53452
rect 35300 53398 35302 53450
rect 35302 53398 35354 53450
rect 35354 53398 35356 53450
rect 35300 53396 35356 53398
rect 35404 53450 35460 53452
rect 35404 53398 35406 53450
rect 35406 53398 35458 53450
rect 35458 53398 35460 53450
rect 35404 53396 35460 53398
rect 50556 52442 50612 52444
rect 50556 52390 50558 52442
rect 50558 52390 50610 52442
rect 50610 52390 50612 52442
rect 50556 52388 50612 52390
rect 50660 52442 50716 52444
rect 50660 52390 50662 52442
rect 50662 52390 50714 52442
rect 50714 52390 50716 52442
rect 50660 52388 50716 52390
rect 50764 52442 50820 52444
rect 50764 52390 50766 52442
rect 50766 52390 50818 52442
rect 50818 52390 50820 52442
rect 50764 52388 50820 52390
rect 35196 51434 35252 51436
rect 35196 51382 35198 51434
rect 35198 51382 35250 51434
rect 35250 51382 35252 51434
rect 35196 51380 35252 51382
rect 35300 51434 35356 51436
rect 35300 51382 35302 51434
rect 35302 51382 35354 51434
rect 35354 51382 35356 51434
rect 35300 51380 35356 51382
rect 35404 51434 35460 51436
rect 35404 51382 35406 51434
rect 35406 51382 35458 51434
rect 35458 51382 35460 51434
rect 35404 51380 35460 51382
rect 50556 50426 50612 50428
rect 50556 50374 50558 50426
rect 50558 50374 50610 50426
rect 50610 50374 50612 50426
rect 50556 50372 50612 50374
rect 50660 50426 50716 50428
rect 50660 50374 50662 50426
rect 50662 50374 50714 50426
rect 50714 50374 50716 50426
rect 50660 50372 50716 50374
rect 50764 50426 50820 50428
rect 50764 50374 50766 50426
rect 50766 50374 50818 50426
rect 50818 50374 50820 50426
rect 50764 50372 50820 50374
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 36988 48972 37044 49028
rect 31276 48914 31332 48916
rect 31276 48862 31278 48914
rect 31278 48862 31330 48914
rect 31330 48862 31332 48914
rect 31276 48860 31332 48862
rect 30828 48802 30884 48804
rect 30828 48750 30830 48802
rect 30830 48750 30882 48802
rect 30882 48750 30884 48802
rect 30828 48748 30884 48750
rect 29708 46674 29764 46676
rect 29708 46622 29710 46674
rect 29710 46622 29762 46674
rect 29762 46622 29764 46674
rect 29708 46620 29764 46622
rect 30940 45388 30996 45444
rect 30268 45276 30324 45332
rect 29932 44882 29988 44884
rect 29932 44830 29934 44882
rect 29934 44830 29986 44882
rect 29986 44830 29988 44882
rect 29932 44828 29988 44830
rect 29932 43932 29988 43988
rect 32732 48914 32788 48916
rect 32732 48862 32734 48914
rect 32734 48862 32786 48914
rect 32786 48862 32788 48914
rect 32732 48860 32788 48862
rect 31948 48802 32004 48804
rect 31948 48750 31950 48802
rect 31950 48750 32002 48802
rect 32002 48750 32004 48802
rect 31948 48748 32004 48750
rect 31500 46620 31556 46676
rect 37436 48972 37492 49028
rect 40348 48972 40404 49028
rect 35196 47402 35252 47404
rect 35196 47350 35198 47402
rect 35198 47350 35250 47402
rect 35250 47350 35252 47402
rect 35196 47348 35252 47350
rect 35300 47402 35356 47404
rect 35300 47350 35302 47402
rect 35302 47350 35354 47402
rect 35354 47350 35356 47402
rect 35300 47348 35356 47350
rect 35404 47402 35460 47404
rect 35404 47350 35406 47402
rect 35406 47350 35458 47402
rect 35458 47350 35460 47402
rect 35404 47348 35460 47350
rect 31948 45724 32004 45780
rect 31276 45276 31332 45332
rect 31948 44828 32004 44884
rect 32620 46620 32676 46676
rect 33292 45724 33348 45780
rect 33180 45276 33236 45332
rect 33180 44044 33236 44100
rect 31276 43708 31332 43764
rect 32284 43762 32340 43764
rect 32284 43710 32286 43762
rect 32286 43710 32338 43762
rect 32338 43710 32340 43762
rect 32284 43708 32340 43710
rect 29820 42642 29876 42644
rect 29820 42590 29822 42642
rect 29822 42590 29874 42642
rect 29874 42590 29876 42642
rect 29820 42588 29876 42590
rect 34636 45778 34692 45780
rect 34636 45726 34638 45778
rect 34638 45726 34690 45778
rect 34690 45726 34692 45778
rect 34636 45724 34692 45726
rect 35084 45890 35140 45892
rect 35084 45838 35086 45890
rect 35086 45838 35138 45890
rect 35138 45838 35140 45890
rect 35084 45836 35140 45838
rect 35196 45386 35252 45388
rect 35196 45334 35198 45386
rect 35198 45334 35250 45386
rect 35250 45334 35252 45386
rect 35196 45332 35252 45334
rect 35300 45386 35356 45388
rect 35300 45334 35302 45386
rect 35302 45334 35354 45386
rect 35354 45334 35356 45386
rect 35300 45332 35356 45334
rect 35404 45386 35460 45388
rect 35404 45334 35406 45386
rect 35406 45334 35458 45386
rect 35458 45334 35460 45386
rect 35404 45332 35460 45334
rect 33516 43874 33572 43876
rect 33516 43822 33518 43874
rect 33518 43822 33570 43874
rect 33570 43822 33572 43874
rect 33516 43820 33572 43822
rect 33180 43708 33236 43764
rect 34412 44044 34468 44100
rect 33292 42754 33348 42756
rect 33292 42702 33294 42754
rect 33294 42702 33346 42754
rect 33346 42702 33348 42754
rect 33292 42700 33348 42702
rect 32060 41916 32116 41972
rect 30044 41858 30100 41860
rect 30044 41806 30046 41858
rect 30046 41806 30098 41858
rect 30098 41806 30100 41858
rect 30044 41804 30100 41806
rect 30492 41746 30548 41748
rect 30492 41694 30494 41746
rect 30494 41694 30546 41746
rect 30546 41694 30548 41746
rect 30492 41692 30548 41694
rect 30380 40908 30436 40964
rect 29820 40738 29876 40740
rect 29820 40686 29822 40738
rect 29822 40686 29874 40738
rect 29874 40686 29876 40738
rect 29820 40684 29876 40686
rect 29820 40348 29876 40404
rect 30268 40236 30324 40292
rect 29372 36764 29428 36820
rect 29260 36706 29316 36708
rect 29260 36654 29262 36706
rect 29262 36654 29314 36706
rect 29314 36654 29316 36706
rect 29260 36652 29316 36654
rect 28028 35308 28084 35364
rect 28028 34466 28084 34468
rect 28028 34414 28030 34466
rect 28030 34414 28082 34466
rect 28082 34414 28084 34466
rect 28028 34412 28084 34414
rect 28588 34578 28644 34580
rect 28588 34526 28590 34578
rect 28590 34526 28642 34578
rect 28642 34526 28644 34578
rect 28588 34524 28644 34526
rect 28700 33794 28756 33796
rect 28700 33742 28702 33794
rect 28702 33742 28754 33794
rect 28754 33742 28756 33794
rect 28700 33740 28756 33742
rect 29260 34524 29316 34580
rect 29484 34412 29540 34468
rect 29036 33628 29092 33684
rect 27020 32786 27076 32788
rect 27020 32734 27022 32786
rect 27022 32734 27074 32786
rect 27074 32734 27076 32786
rect 27020 32732 27076 32734
rect 27916 33068 27972 33124
rect 28364 33068 28420 33124
rect 28588 32732 28644 32788
rect 26684 31052 26740 31108
rect 27020 32172 27076 32228
rect 26684 30546 26740 30548
rect 26684 30494 26686 30546
rect 26686 30494 26738 30546
rect 26738 30494 26740 30546
rect 26684 30492 26740 30494
rect 27692 32450 27748 32452
rect 27692 32398 27694 32450
rect 27694 32398 27746 32450
rect 27746 32398 27748 32450
rect 27692 32396 27748 32398
rect 27580 32172 27636 32228
rect 27356 31948 27412 32004
rect 27468 31724 27524 31780
rect 27020 31612 27076 31668
rect 26908 31442 26964 31444
rect 26908 31390 26910 31442
rect 26910 31390 26962 31442
rect 26962 31390 26964 31442
rect 26908 31388 26964 31390
rect 26908 30658 26964 30660
rect 26908 30606 26910 30658
rect 26910 30606 26962 30658
rect 26962 30606 26964 30658
rect 26908 30604 26964 30606
rect 25788 29932 25844 29988
rect 25564 29874 25620 29876
rect 25564 29822 25566 29874
rect 25566 29822 25618 29874
rect 25618 29822 25620 29874
rect 25564 29820 25620 29822
rect 25676 29708 25732 29764
rect 24892 27916 24948 27972
rect 24668 27746 24724 27748
rect 24668 27694 24670 27746
rect 24670 27694 24722 27746
rect 24722 27694 24724 27746
rect 24668 27692 24724 27694
rect 24556 26796 24612 26852
rect 26572 29708 26628 29764
rect 26348 28812 26404 28868
rect 25900 28530 25956 28532
rect 25900 28478 25902 28530
rect 25902 28478 25954 28530
rect 25954 28478 25956 28530
rect 25900 28476 25956 28478
rect 26124 28364 26180 28420
rect 25228 27970 25284 27972
rect 25228 27918 25230 27970
rect 25230 27918 25282 27970
rect 25282 27918 25284 27970
rect 25228 27916 25284 27918
rect 25228 27020 25284 27076
rect 24332 26402 24388 26404
rect 24332 26350 24334 26402
rect 24334 26350 24386 26402
rect 24386 26350 24388 26402
rect 24332 26348 24388 26350
rect 24220 26236 24276 26292
rect 24668 26738 24724 26740
rect 24668 26686 24670 26738
rect 24670 26686 24722 26738
rect 24722 26686 24724 26738
rect 24668 26684 24724 26686
rect 25004 26684 25060 26740
rect 24444 26012 24500 26068
rect 24556 26572 24612 26628
rect 23212 21644 23268 21700
rect 23772 20802 23828 20804
rect 23772 20750 23774 20802
rect 23774 20750 23826 20802
rect 23826 20750 23828 20802
rect 23772 20748 23828 20750
rect 22764 20188 22820 20244
rect 22204 19852 22260 19908
rect 22316 20076 22372 20132
rect 21756 19740 21812 19796
rect 21420 18732 21476 18788
rect 22876 20076 22932 20132
rect 20748 18508 20804 18564
rect 19964 17612 20020 17668
rect 19292 16716 19348 16772
rect 18620 16604 18676 16660
rect 19180 16322 19236 16324
rect 19180 16270 19182 16322
rect 19182 16270 19234 16322
rect 19234 16270 19236 16322
rect 19180 16268 19236 16270
rect 20412 17666 20468 17668
rect 20412 17614 20414 17666
rect 20414 17614 20466 17666
rect 20466 17614 20468 17666
rect 20412 17612 20468 17614
rect 20076 16716 20132 16772
rect 20524 16604 20580 16660
rect 20188 16434 20244 16436
rect 20188 16382 20190 16434
rect 20190 16382 20242 16434
rect 20242 16382 20244 16434
rect 20188 16380 20244 16382
rect 19836 16154 19892 16156
rect 19836 16102 19838 16154
rect 19838 16102 19890 16154
rect 19890 16102 19892 16154
rect 19836 16100 19892 16102
rect 19940 16154 19996 16156
rect 19940 16102 19942 16154
rect 19942 16102 19994 16154
rect 19994 16102 19996 16154
rect 19940 16100 19996 16102
rect 20044 16154 20100 16156
rect 20044 16102 20046 16154
rect 20046 16102 20098 16154
rect 20098 16102 20100 16154
rect 20044 16100 20100 16102
rect 20748 15820 20804 15876
rect 21084 16268 21140 16324
rect 20860 15596 20916 15652
rect 21308 16604 21364 16660
rect 21308 15596 21364 15652
rect 20300 14754 20356 14756
rect 20300 14702 20302 14754
rect 20302 14702 20354 14754
rect 20354 14702 20356 14754
rect 20300 14700 20356 14702
rect 19852 14418 19908 14420
rect 19852 14366 19854 14418
rect 19854 14366 19906 14418
rect 19906 14366 19908 14418
rect 19852 14364 19908 14366
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 18620 13468 18676 13524
rect 19404 13522 19460 13524
rect 19404 13470 19406 13522
rect 19406 13470 19458 13522
rect 19458 13470 19460 13522
rect 19404 13468 19460 13470
rect 18284 12236 18340 12292
rect 19836 12122 19892 12124
rect 19836 12070 19838 12122
rect 19838 12070 19890 12122
rect 19890 12070 19892 12122
rect 19836 12068 19892 12070
rect 19940 12122 19996 12124
rect 19940 12070 19942 12122
rect 19942 12070 19994 12122
rect 19994 12070 19996 12122
rect 19940 12068 19996 12070
rect 20044 12122 20100 12124
rect 20044 12070 20046 12122
rect 20046 12070 20098 12122
rect 20098 12070 20100 12122
rect 20044 12068 20100 12070
rect 4476 11114 4532 11116
rect 4476 11062 4478 11114
rect 4478 11062 4530 11114
rect 4530 11062 4532 11114
rect 4476 11060 4532 11062
rect 4580 11114 4636 11116
rect 4580 11062 4582 11114
rect 4582 11062 4634 11114
rect 4634 11062 4636 11114
rect 4580 11060 4636 11062
rect 4684 11114 4740 11116
rect 4684 11062 4686 11114
rect 4686 11062 4738 11114
rect 4738 11062 4740 11114
rect 4684 11060 4740 11062
rect 16380 10108 16436 10164
rect 17500 10108 17556 10164
rect 16940 9996 16996 10052
rect 19068 10610 19124 10612
rect 19068 10558 19070 10610
rect 19070 10558 19122 10610
rect 19122 10558 19124 10610
rect 19068 10556 19124 10558
rect 19852 10556 19908 10612
rect 19740 10386 19796 10388
rect 19740 10334 19742 10386
rect 19742 10334 19794 10386
rect 19794 10334 19796 10386
rect 19740 10332 19796 10334
rect 18396 10108 18452 10164
rect 18284 9996 18340 10052
rect 18284 9436 18340 9492
rect 19836 10106 19892 10108
rect 19836 10054 19838 10106
rect 19838 10054 19890 10106
rect 19890 10054 19892 10106
rect 19836 10052 19892 10054
rect 19940 10106 19996 10108
rect 19940 10054 19942 10106
rect 19942 10054 19994 10106
rect 19994 10054 19996 10106
rect 19940 10052 19996 10054
rect 20044 10106 20100 10108
rect 20044 10054 20046 10106
rect 20046 10054 20098 10106
rect 20098 10054 20100 10106
rect 20044 10052 20100 10054
rect 19628 9602 19684 9604
rect 19628 9550 19630 9602
rect 19630 9550 19682 9602
rect 19682 9550 19684 9602
rect 19628 9548 19684 9550
rect 4476 9098 4532 9100
rect 4476 9046 4478 9098
rect 4478 9046 4530 9098
rect 4530 9046 4532 9098
rect 4476 9044 4532 9046
rect 4580 9098 4636 9100
rect 4580 9046 4582 9098
rect 4582 9046 4634 9098
rect 4634 9046 4636 9098
rect 4580 9044 4636 9046
rect 4684 9098 4740 9100
rect 4684 9046 4686 9098
rect 4686 9046 4738 9098
rect 4738 9046 4740 9098
rect 4684 9044 4740 9046
rect 18956 9490 19012 9492
rect 18956 9438 18958 9490
rect 18958 9438 19010 9490
rect 19010 9438 19012 9490
rect 18956 9436 19012 9438
rect 18956 8482 19012 8484
rect 18956 8430 18958 8482
rect 18958 8430 19010 8482
rect 19010 8430 19012 8482
rect 18956 8428 19012 8430
rect 19516 8764 19572 8820
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4620 6748 4676 6804
rect 4172 6354 4228 6356
rect 4172 6302 4174 6354
rect 4174 6302 4226 6354
rect 4226 6302 4228 6354
rect 4172 6300 4228 6302
rect 20188 9436 20244 9492
rect 19852 8706 19908 8708
rect 19852 8654 19854 8706
rect 19854 8654 19906 8706
rect 19906 8654 19908 8706
rect 19852 8652 19908 8654
rect 20300 9548 20356 9604
rect 20636 11452 20692 11508
rect 20636 10780 20692 10836
rect 20636 9548 20692 9604
rect 20524 8764 20580 8820
rect 20972 14700 21028 14756
rect 21980 16716 22036 16772
rect 21868 16380 21924 16436
rect 21644 15820 21700 15876
rect 21420 14252 21476 14308
rect 23212 18844 23268 18900
rect 23996 23884 24052 23940
rect 24332 23772 24388 23828
rect 23996 23660 24052 23716
rect 22876 18562 22932 18564
rect 22876 18510 22878 18562
rect 22878 18510 22930 18562
rect 22930 18510 22932 18562
rect 22876 18508 22932 18510
rect 25116 26012 25172 26068
rect 24556 25618 24612 25620
rect 24556 25566 24558 25618
rect 24558 25566 24610 25618
rect 24610 25566 24612 25618
rect 24556 25564 24612 25566
rect 24668 24722 24724 24724
rect 24668 24670 24670 24722
rect 24670 24670 24722 24722
rect 24722 24670 24724 24722
rect 24668 24668 24724 24670
rect 24556 24610 24612 24612
rect 24556 24558 24558 24610
rect 24558 24558 24610 24610
rect 24610 24558 24612 24610
rect 24556 24556 24612 24558
rect 24444 23660 24500 23716
rect 24668 23490 24724 23492
rect 24668 23438 24670 23490
rect 24670 23438 24722 23490
rect 24722 23438 24724 23490
rect 24668 23436 24724 23438
rect 24668 22540 24724 22596
rect 24668 21586 24724 21588
rect 24668 21534 24670 21586
rect 24670 21534 24722 21586
rect 24722 21534 24724 21586
rect 24668 21532 24724 21534
rect 24220 21196 24276 21252
rect 24668 20802 24724 20804
rect 24668 20750 24670 20802
rect 24670 20750 24722 20802
rect 24722 20750 24724 20802
rect 24668 20748 24724 20750
rect 24108 20188 24164 20244
rect 24892 25676 24948 25732
rect 25676 26738 25732 26740
rect 25676 26686 25678 26738
rect 25678 26686 25730 26738
rect 25730 26686 25732 26738
rect 25676 26684 25732 26686
rect 26012 26908 26068 26964
rect 26572 28476 26628 28532
rect 26796 30268 26852 30324
rect 27020 30044 27076 30100
rect 27132 31388 27188 31444
rect 27356 30268 27412 30324
rect 27132 29820 27188 29876
rect 27580 31106 27636 31108
rect 27580 31054 27582 31106
rect 27582 31054 27634 31106
rect 27634 31054 27636 31106
rect 27580 31052 27636 31054
rect 27916 30770 27972 30772
rect 27916 30718 27918 30770
rect 27918 30718 27970 30770
rect 27970 30718 27972 30770
rect 27916 30716 27972 30718
rect 28364 32002 28420 32004
rect 28364 31950 28366 32002
rect 28366 31950 28418 32002
rect 28418 31950 28420 32002
rect 28364 31948 28420 31950
rect 30044 38946 30100 38948
rect 30044 38894 30046 38946
rect 30046 38894 30098 38946
rect 30098 38894 30100 38946
rect 30044 38892 30100 38894
rect 30716 40460 30772 40516
rect 31164 40738 31220 40740
rect 31164 40686 31166 40738
rect 31166 40686 31218 40738
rect 31218 40686 31220 40738
rect 31164 40684 31220 40686
rect 30604 38892 30660 38948
rect 30716 36818 30772 36820
rect 30716 36766 30718 36818
rect 30718 36766 30770 36818
rect 30770 36766 30772 36818
rect 30716 36764 30772 36766
rect 30156 36034 30212 36036
rect 30156 35982 30158 36034
rect 30158 35982 30210 36034
rect 30210 35982 30212 36034
rect 30156 35980 30212 35982
rect 29932 32844 29988 32900
rect 30716 33628 30772 33684
rect 29820 31724 29876 31780
rect 28252 30882 28308 30884
rect 28252 30830 28254 30882
rect 28254 30830 28306 30882
rect 28306 30830 28308 30882
rect 28252 30828 28308 30830
rect 30940 31836 30996 31892
rect 35868 45724 35924 45780
rect 35980 45836 36036 45892
rect 36316 47794 36372 47796
rect 36316 47742 36318 47794
rect 36318 47742 36370 47794
rect 36370 47742 36372 47794
rect 36316 47740 36372 47742
rect 37100 47740 37156 47796
rect 40012 48636 40068 48692
rect 38108 47740 38164 47796
rect 35980 44940 36036 44996
rect 35644 44658 35700 44660
rect 35644 44606 35646 44658
rect 35646 44606 35698 44658
rect 35698 44606 35700 44658
rect 35644 44604 35700 44606
rect 36092 45724 36148 45780
rect 35644 44098 35700 44100
rect 35644 44046 35646 44098
rect 35646 44046 35698 44098
rect 35698 44046 35700 44098
rect 35644 44044 35700 44046
rect 35532 43820 35588 43876
rect 39004 46898 39060 46900
rect 39004 46846 39006 46898
rect 39006 46846 39058 46898
rect 39058 46846 39060 46898
rect 39004 46844 39060 46846
rect 38332 45276 38388 45332
rect 37660 44994 37716 44996
rect 37660 44942 37662 44994
rect 37662 44942 37714 44994
rect 37714 44942 37716 44994
rect 37660 44940 37716 44942
rect 36428 44658 36484 44660
rect 36428 44606 36430 44658
rect 36430 44606 36482 44658
rect 36482 44606 36484 44658
rect 36428 44604 36484 44606
rect 36764 43874 36820 43876
rect 36764 43822 36766 43874
rect 36766 43822 36818 43874
rect 36818 43822 36820 43874
rect 36764 43820 36820 43822
rect 37212 44658 37268 44660
rect 37212 44606 37214 44658
rect 37214 44606 37266 44658
rect 37266 44606 37268 44658
rect 37212 44604 37268 44606
rect 36092 43708 36148 43764
rect 37100 43708 37156 43764
rect 33404 41970 33460 41972
rect 33404 41918 33406 41970
rect 33406 41918 33458 41970
rect 33458 41918 33460 41970
rect 33404 41916 33460 41918
rect 34636 41970 34692 41972
rect 34636 41918 34638 41970
rect 34638 41918 34690 41970
rect 34690 41918 34692 41970
rect 34636 41916 34692 41918
rect 32732 41132 32788 41188
rect 32508 40684 32564 40740
rect 31612 40236 31668 40292
rect 32508 40236 32564 40292
rect 33068 40236 33124 40292
rect 35196 43370 35252 43372
rect 35196 43318 35198 43370
rect 35198 43318 35250 43370
rect 35250 43318 35252 43370
rect 35196 43316 35252 43318
rect 35300 43370 35356 43372
rect 35300 43318 35302 43370
rect 35302 43318 35354 43370
rect 35354 43318 35356 43370
rect 35300 43316 35356 43318
rect 35404 43370 35460 43372
rect 35404 43318 35406 43370
rect 35406 43318 35458 43370
rect 35458 43318 35460 43370
rect 35404 43316 35460 43318
rect 35308 42754 35364 42756
rect 35308 42702 35310 42754
rect 35310 42702 35362 42754
rect 35362 42702 35364 42754
rect 35308 42700 35364 42702
rect 35196 41354 35252 41356
rect 35196 41302 35198 41354
rect 35198 41302 35250 41354
rect 35250 41302 35252 41354
rect 35196 41300 35252 41302
rect 35300 41354 35356 41356
rect 35300 41302 35302 41354
rect 35302 41302 35354 41354
rect 35354 41302 35356 41354
rect 35300 41300 35356 41302
rect 35404 41354 35460 41356
rect 35404 41302 35406 41354
rect 35406 41302 35458 41354
rect 35458 41302 35460 41354
rect 35404 41300 35460 41302
rect 34972 41132 35028 41188
rect 34412 40684 34468 40740
rect 34076 40348 34132 40404
rect 38780 44940 38836 44996
rect 39900 46674 39956 46676
rect 39900 46622 39902 46674
rect 39902 46622 39954 46674
rect 39954 46622 39956 46674
rect 39900 46620 39956 46622
rect 41244 48860 41300 48916
rect 40796 48802 40852 48804
rect 40796 48750 40798 48802
rect 40798 48750 40850 48802
rect 40850 48750 40852 48802
rect 40796 48748 40852 48750
rect 40236 46898 40292 46900
rect 40236 46846 40238 46898
rect 40238 46846 40290 46898
rect 40290 46846 40292 46898
rect 40236 46844 40292 46846
rect 40684 46620 40740 46676
rect 41132 46844 41188 46900
rect 40124 46172 40180 46228
rect 40908 46172 40964 46228
rect 39004 45388 39060 45444
rect 37996 43820 38052 43876
rect 37436 41804 37492 41860
rect 37324 40908 37380 40964
rect 36764 40684 36820 40740
rect 37100 40460 37156 40516
rect 35532 39788 35588 39844
rect 36428 39676 36484 39732
rect 35644 39564 35700 39620
rect 33628 38892 33684 38948
rect 34412 38946 34468 38948
rect 34412 38894 34414 38946
rect 34414 38894 34466 38946
rect 34466 38894 34468 38946
rect 34412 38892 34468 38894
rect 32508 37714 32564 37716
rect 32508 37662 32510 37714
rect 32510 37662 32562 37714
rect 32562 37662 32564 37714
rect 32508 37660 32564 37662
rect 32172 35810 32228 35812
rect 32172 35758 32174 35810
rect 32174 35758 32226 35810
rect 32226 35758 32228 35810
rect 32172 35756 32228 35758
rect 32060 34802 32116 34804
rect 32060 34750 32062 34802
rect 32062 34750 32114 34802
rect 32114 34750 32116 34802
rect 32060 34748 32116 34750
rect 32060 33740 32116 33796
rect 31612 32844 31668 32900
rect 29708 30716 29764 30772
rect 28588 30380 28644 30436
rect 29148 30604 29204 30660
rect 29036 30268 29092 30324
rect 28140 30098 28196 30100
rect 28140 30046 28142 30098
rect 28142 30046 28194 30098
rect 28194 30046 28196 30098
rect 28140 30044 28196 30046
rect 27692 29708 27748 29764
rect 27020 29484 27076 29540
rect 27468 29596 27524 29652
rect 26908 28924 26964 28980
rect 27020 28364 27076 28420
rect 26348 27746 26404 27748
rect 26348 27694 26350 27746
rect 26350 27694 26402 27746
rect 26402 27694 26404 27746
rect 26348 27692 26404 27694
rect 25564 26460 25620 26516
rect 25340 25452 25396 25508
rect 25564 25564 25620 25620
rect 25228 25340 25284 25396
rect 25452 24668 25508 24724
rect 25340 24610 25396 24612
rect 25340 24558 25342 24610
rect 25342 24558 25394 24610
rect 25394 24558 25396 24610
rect 25340 24556 25396 24558
rect 26348 27020 26404 27076
rect 28476 29596 28532 29652
rect 28924 29650 28980 29652
rect 28924 29598 28926 29650
rect 28926 29598 28978 29650
rect 28978 29598 28980 29650
rect 28924 29596 28980 29598
rect 29036 29372 29092 29428
rect 27580 28866 27636 28868
rect 27580 28814 27582 28866
rect 27582 28814 27634 28866
rect 27634 28814 27636 28866
rect 27580 28812 27636 28814
rect 29260 30380 29316 30436
rect 29596 30156 29652 30212
rect 29260 29762 29316 29764
rect 29260 29710 29262 29762
rect 29262 29710 29314 29762
rect 29314 29710 29316 29762
rect 29260 29708 29316 29710
rect 29148 28700 29204 28756
rect 29484 28812 29540 28868
rect 29932 29762 29988 29764
rect 29932 29710 29934 29762
rect 29934 29710 29986 29762
rect 29986 29710 29988 29762
rect 29932 29708 29988 29710
rect 29820 29148 29876 29204
rect 29820 27916 29876 27972
rect 29596 26908 29652 26964
rect 29708 27580 29764 27636
rect 26908 26012 26964 26068
rect 26124 25900 26180 25956
rect 25900 25730 25956 25732
rect 25900 25678 25902 25730
rect 25902 25678 25954 25730
rect 25954 25678 25956 25730
rect 25900 25676 25956 25678
rect 25788 25228 25844 25284
rect 26124 24668 26180 24724
rect 25676 24444 25732 24500
rect 25228 23660 25284 23716
rect 25116 22540 25172 22596
rect 25116 21196 25172 21252
rect 24556 19570 24612 19572
rect 24556 19518 24558 19570
rect 24558 19518 24610 19570
rect 24610 19518 24612 19570
rect 24556 19516 24612 19518
rect 23548 17836 23604 17892
rect 24444 17836 24500 17892
rect 23772 16716 23828 16772
rect 22988 16434 23044 16436
rect 22988 16382 22990 16434
rect 22990 16382 23042 16434
rect 23042 16382 23044 16434
rect 22988 16380 23044 16382
rect 22988 15820 23044 15876
rect 22988 15650 23044 15652
rect 22988 15598 22990 15650
rect 22990 15598 23042 15650
rect 23042 15598 23044 15650
rect 22988 15596 23044 15598
rect 24220 15820 24276 15876
rect 23884 15708 23940 15764
rect 22428 14700 22484 14756
rect 21420 13858 21476 13860
rect 21420 13806 21422 13858
rect 21422 13806 21474 13858
rect 21474 13806 21476 13858
rect 21420 13804 21476 13806
rect 21644 13692 21700 13748
rect 21308 12236 21364 12292
rect 21084 10556 21140 10612
rect 22316 14252 22372 14308
rect 22316 13746 22372 13748
rect 22316 13694 22318 13746
rect 22318 13694 22370 13746
rect 22370 13694 22372 13746
rect 22316 13692 22372 13694
rect 25004 16716 25060 16772
rect 24668 15708 24724 15764
rect 24332 15650 24388 15652
rect 24332 15598 24334 15650
rect 24334 15598 24386 15650
rect 24386 15598 24388 15650
rect 24332 15596 24388 15598
rect 23212 13858 23268 13860
rect 23212 13806 23214 13858
rect 23214 13806 23266 13858
rect 23266 13806 23268 13858
rect 23212 13804 23268 13806
rect 24220 13858 24276 13860
rect 24220 13806 24222 13858
rect 24222 13806 24274 13858
rect 24274 13806 24276 13858
rect 24220 13804 24276 13806
rect 22876 11954 22932 11956
rect 22876 11902 22878 11954
rect 22878 11902 22930 11954
rect 22930 11902 22932 11954
rect 22876 11900 22932 11902
rect 22316 11564 22372 11620
rect 21980 11340 22036 11396
rect 21980 10780 22036 10836
rect 21308 10498 21364 10500
rect 21308 10446 21310 10498
rect 21310 10446 21362 10498
rect 21362 10446 21364 10498
rect 21308 10444 21364 10446
rect 20860 8652 20916 8708
rect 20188 8540 20244 8596
rect 19852 8428 19908 8484
rect 19836 8090 19892 8092
rect 19836 8038 19838 8090
rect 19838 8038 19890 8090
rect 19890 8038 19892 8090
rect 19836 8036 19892 8038
rect 19940 8090 19996 8092
rect 19940 8038 19942 8090
rect 19942 8038 19994 8090
rect 19994 8038 19996 8090
rect 19940 8036 19996 8038
rect 20044 8090 20100 8092
rect 20044 8038 20046 8090
rect 20046 8038 20098 8090
rect 20098 8038 20100 8090
rect 20044 8036 20100 8038
rect 20748 8540 20804 8596
rect 20636 8428 20692 8484
rect 21532 8652 21588 8708
rect 20412 6636 20468 6692
rect 19404 6524 19460 6580
rect 20076 6524 20132 6580
rect 18172 6354 18228 6356
rect 18172 6302 18174 6354
rect 18174 6302 18226 6354
rect 18226 6302 18228 6354
rect 18172 6300 18228 6302
rect 19836 6074 19892 6076
rect 19836 6022 19838 6074
rect 19838 6022 19890 6074
rect 19890 6022 19892 6074
rect 19836 6020 19892 6022
rect 19940 6074 19996 6076
rect 19940 6022 19942 6074
rect 19942 6022 19994 6074
rect 19994 6022 19996 6074
rect 19940 6020 19996 6022
rect 20044 6074 20100 6076
rect 20044 6022 20046 6074
rect 20046 6022 20098 6074
rect 20098 6022 20100 6074
rect 20044 6020 20100 6022
rect 21196 6578 21252 6580
rect 21196 6526 21198 6578
rect 21198 6526 21250 6578
rect 21250 6526 21252 6578
rect 21196 6524 21252 6526
rect 20636 6412 20692 6468
rect 20524 6354 20580 6356
rect 20524 6302 20526 6354
rect 20526 6302 20578 6354
rect 20578 6302 20580 6354
rect 20524 6300 20580 6302
rect 21980 10610 22036 10612
rect 21980 10558 21982 10610
rect 21982 10558 22034 10610
rect 22034 10558 22036 10610
rect 21980 10556 22036 10558
rect 22428 10332 22484 10388
rect 23100 11730 23156 11732
rect 23100 11678 23102 11730
rect 23102 11678 23154 11730
rect 23154 11678 23156 11730
rect 23100 11676 23156 11678
rect 24668 14588 24724 14644
rect 24444 14530 24500 14532
rect 24444 14478 24446 14530
rect 24446 14478 24498 14530
rect 24498 14478 24500 14530
rect 24444 14476 24500 14478
rect 24444 13804 24500 13860
rect 23548 11618 23604 11620
rect 23548 11566 23550 11618
rect 23550 11566 23602 11618
rect 23602 11566 23604 11618
rect 23548 11564 23604 11566
rect 23324 11340 23380 11396
rect 22204 8482 22260 8484
rect 22204 8430 22206 8482
rect 22206 8430 22258 8482
rect 22258 8430 22260 8482
rect 22204 8428 22260 8430
rect 22876 10108 22932 10164
rect 21532 7532 21588 7588
rect 22540 7644 22596 7700
rect 21980 6636 22036 6692
rect 22204 6300 22260 6356
rect 23436 11452 23492 11508
rect 24332 11900 24388 11956
rect 25004 11900 25060 11956
rect 23884 8764 23940 8820
rect 23660 8594 23716 8596
rect 23660 8542 23662 8594
rect 23662 8542 23714 8594
rect 23714 8542 23716 8594
rect 23660 8540 23716 8542
rect 24220 11618 24276 11620
rect 24220 11566 24222 11618
rect 24222 11566 24274 11618
rect 24274 11566 24276 11618
rect 24220 11564 24276 11566
rect 25788 23996 25844 24052
rect 25788 23826 25844 23828
rect 25788 23774 25790 23826
rect 25790 23774 25842 23826
rect 25842 23774 25844 23826
rect 25788 23772 25844 23774
rect 25788 23548 25844 23604
rect 25564 22594 25620 22596
rect 25564 22542 25566 22594
rect 25566 22542 25618 22594
rect 25618 22542 25620 22594
rect 25564 22540 25620 22542
rect 25676 21810 25732 21812
rect 25676 21758 25678 21810
rect 25678 21758 25730 21810
rect 25730 21758 25732 21810
rect 25676 21756 25732 21758
rect 25452 21586 25508 21588
rect 25452 21534 25454 21586
rect 25454 21534 25506 21586
rect 25506 21534 25508 21586
rect 25452 21532 25508 21534
rect 26572 25900 26628 25956
rect 26348 25340 26404 25396
rect 26684 25788 26740 25844
rect 27020 25842 27076 25844
rect 27020 25790 27022 25842
rect 27022 25790 27074 25842
rect 27074 25790 27076 25842
rect 27020 25788 27076 25790
rect 27356 26514 27412 26516
rect 27356 26462 27358 26514
rect 27358 26462 27410 26514
rect 27410 26462 27412 26514
rect 27356 26460 27412 26462
rect 26572 25564 26628 25620
rect 26460 24722 26516 24724
rect 26460 24670 26462 24722
rect 26462 24670 26514 24722
rect 26514 24670 26516 24722
rect 26460 24668 26516 24670
rect 26908 25340 26964 25396
rect 26796 25058 26852 25060
rect 26796 25006 26798 25058
rect 26798 25006 26850 25058
rect 26850 25006 26852 25058
rect 26796 25004 26852 25006
rect 26460 24444 26516 24500
rect 26348 24050 26404 24052
rect 26348 23998 26350 24050
rect 26350 23998 26402 24050
rect 26402 23998 26404 24050
rect 26348 23996 26404 23998
rect 26684 23884 26740 23940
rect 26684 23548 26740 23604
rect 26348 23436 26404 23492
rect 27244 25340 27300 25396
rect 27244 23938 27300 23940
rect 27244 23886 27246 23938
rect 27246 23886 27298 23938
rect 27298 23886 27300 23938
rect 27244 23884 27300 23886
rect 26796 22876 26852 22932
rect 26908 22594 26964 22596
rect 26908 22542 26910 22594
rect 26910 22542 26962 22594
rect 26962 22542 26964 22594
rect 26908 22540 26964 22542
rect 27692 25564 27748 25620
rect 27468 24610 27524 24612
rect 27468 24558 27470 24610
rect 27470 24558 27522 24610
rect 27522 24558 27524 24610
rect 27468 24556 27524 24558
rect 27916 25900 27972 25956
rect 29484 26236 29540 26292
rect 28588 25900 28644 25956
rect 29372 25954 29428 25956
rect 29372 25902 29374 25954
rect 29374 25902 29426 25954
rect 29426 25902 29428 25954
rect 29372 25900 29428 25902
rect 28028 25618 28084 25620
rect 28028 25566 28030 25618
rect 28030 25566 28082 25618
rect 28082 25566 28084 25618
rect 28028 25564 28084 25566
rect 28588 25564 28644 25620
rect 27580 24444 27636 24500
rect 27692 24332 27748 24388
rect 27468 23884 27524 23940
rect 27580 23826 27636 23828
rect 27580 23774 27582 23826
rect 27582 23774 27634 23826
rect 27634 23774 27636 23826
rect 27580 23772 27636 23774
rect 27468 22876 27524 22932
rect 26236 20972 26292 21028
rect 26348 21756 26404 21812
rect 27356 21810 27412 21812
rect 27356 21758 27358 21810
rect 27358 21758 27410 21810
rect 27410 21758 27412 21810
rect 27356 21756 27412 21758
rect 26460 21698 26516 21700
rect 26460 21646 26462 21698
rect 26462 21646 26514 21698
rect 26514 21646 26516 21698
rect 26460 21644 26516 21646
rect 26796 21196 26852 21252
rect 25340 20188 25396 20244
rect 27244 20466 27300 20468
rect 27244 20414 27246 20466
rect 27246 20414 27298 20466
rect 27298 20414 27300 20466
rect 27244 20412 27300 20414
rect 26012 19906 26068 19908
rect 26012 19854 26014 19906
rect 26014 19854 26066 19906
rect 26066 19854 26068 19906
rect 26012 19852 26068 19854
rect 25228 18844 25284 18900
rect 25676 18450 25732 18452
rect 25676 18398 25678 18450
rect 25678 18398 25730 18450
rect 25730 18398 25732 18450
rect 25676 18396 25732 18398
rect 27356 19740 27412 19796
rect 25340 17554 25396 17556
rect 25340 17502 25342 17554
rect 25342 17502 25394 17554
rect 25394 17502 25396 17554
rect 25340 17500 25396 17502
rect 25340 15820 25396 15876
rect 25788 15762 25844 15764
rect 25788 15710 25790 15762
rect 25790 15710 25842 15762
rect 25842 15710 25844 15762
rect 25788 15708 25844 15710
rect 25452 14476 25508 14532
rect 25788 14364 25844 14420
rect 25452 13858 25508 13860
rect 25452 13806 25454 13858
rect 25454 13806 25506 13858
rect 25506 13806 25508 13858
rect 25452 13804 25508 13806
rect 26012 15650 26068 15652
rect 26012 15598 26014 15650
rect 26014 15598 26066 15650
rect 26066 15598 26068 15650
rect 26012 15596 26068 15598
rect 26348 17890 26404 17892
rect 26348 17838 26350 17890
rect 26350 17838 26402 17890
rect 26402 17838 26404 17890
rect 26348 17836 26404 17838
rect 26908 19570 26964 19572
rect 26908 19518 26910 19570
rect 26910 19518 26962 19570
rect 26962 19518 26964 19570
rect 26908 19516 26964 19518
rect 26684 18898 26740 18900
rect 26684 18846 26686 18898
rect 26686 18846 26738 18898
rect 26738 18846 26740 18898
rect 26684 18844 26740 18846
rect 26572 17724 26628 17780
rect 27356 17500 27412 17556
rect 27244 16770 27300 16772
rect 27244 16718 27246 16770
rect 27246 16718 27298 16770
rect 27298 16718 27300 16770
rect 27244 16716 27300 16718
rect 26012 14642 26068 14644
rect 26012 14590 26014 14642
rect 26014 14590 26066 14642
rect 26066 14590 26068 14642
rect 26012 14588 26068 14590
rect 26236 14530 26292 14532
rect 26236 14478 26238 14530
rect 26238 14478 26290 14530
rect 26290 14478 26292 14530
rect 26236 14476 26292 14478
rect 26348 14364 26404 14420
rect 26236 14252 26292 14308
rect 25116 11676 25172 11732
rect 25340 11730 25396 11732
rect 25340 11678 25342 11730
rect 25342 11678 25394 11730
rect 25394 11678 25396 11730
rect 25340 11676 25396 11678
rect 25004 11452 25060 11508
rect 24108 10386 24164 10388
rect 24108 10334 24110 10386
rect 24110 10334 24162 10386
rect 24162 10334 24164 10386
rect 24108 10332 24164 10334
rect 24220 9996 24276 10052
rect 24668 8764 24724 8820
rect 23996 7644 24052 7700
rect 22988 7586 23044 7588
rect 22988 7534 22990 7586
rect 22990 7534 23042 7586
rect 23042 7534 23044 7586
rect 22988 7532 23044 7534
rect 25340 9996 25396 10052
rect 24892 7868 24948 7924
rect 25004 7532 25060 7588
rect 25116 8540 25172 8596
rect 26572 14306 26628 14308
rect 26572 14254 26574 14306
rect 26574 14254 26626 14306
rect 26626 14254 26628 14306
rect 26572 14252 26628 14254
rect 27020 15260 27076 15316
rect 26684 13804 26740 13860
rect 26796 14700 26852 14756
rect 26908 14642 26964 14644
rect 26908 14590 26910 14642
rect 26910 14590 26962 14642
rect 26962 14590 26964 14642
rect 26908 14588 26964 14590
rect 27132 11788 27188 11844
rect 26348 11506 26404 11508
rect 26348 11454 26350 11506
rect 26350 11454 26402 11506
rect 26402 11454 26404 11506
rect 26348 11452 26404 11454
rect 27804 21532 27860 21588
rect 27804 20188 27860 20244
rect 27692 17500 27748 17556
rect 27468 15372 27524 15428
rect 27580 16268 27636 16324
rect 27468 15148 27524 15204
rect 27468 14588 27524 14644
rect 27356 13356 27412 13412
rect 27804 15036 27860 15092
rect 27692 14418 27748 14420
rect 27692 14366 27694 14418
rect 27694 14366 27746 14418
rect 27746 14366 27748 14418
rect 27692 14364 27748 14366
rect 27020 9996 27076 10052
rect 27244 8540 27300 8596
rect 25116 6636 25172 6692
rect 24332 6524 24388 6580
rect 24668 6524 24724 6580
rect 24332 6300 24388 6356
rect 4476 5066 4532 5068
rect 4476 5014 4478 5066
rect 4478 5014 4530 5066
rect 4530 5014 4532 5066
rect 4476 5012 4532 5014
rect 4580 5066 4636 5068
rect 4580 5014 4582 5066
rect 4582 5014 4634 5066
rect 4634 5014 4636 5066
rect 4580 5012 4636 5014
rect 4684 5066 4740 5068
rect 4684 5014 4686 5066
rect 4686 5014 4738 5066
rect 4738 5014 4740 5066
rect 4684 5012 4740 5014
rect 23996 4674 24052 4676
rect 23996 4622 23998 4674
rect 23998 4622 24050 4674
rect 24050 4622 24052 4674
rect 23996 4620 24052 4622
rect 25228 6524 25284 6580
rect 25900 6524 25956 6580
rect 26124 7586 26180 7588
rect 26124 7534 26126 7586
rect 26126 7534 26178 7586
rect 26178 7534 26180 7586
rect 26124 7532 26180 7534
rect 25340 6354 25396 6356
rect 25340 6302 25342 6354
rect 25342 6302 25394 6354
rect 25394 6302 25396 6354
rect 25340 6300 25396 6302
rect 25452 4674 25508 4676
rect 25452 4622 25454 4674
rect 25454 4622 25506 4674
rect 25506 4622 25508 4674
rect 25452 4620 25508 4622
rect 26348 5458 26404 5460
rect 26348 5406 26350 5458
rect 26350 5406 26402 5458
rect 26402 5406 26404 5458
rect 26348 5404 26404 5406
rect 25900 4620 25956 4676
rect 27804 11788 27860 11844
rect 28924 24556 28980 24612
rect 29260 24556 29316 24612
rect 28028 23772 28084 23828
rect 29596 25564 29652 25620
rect 30828 30658 30884 30660
rect 30828 30606 30830 30658
rect 30830 30606 30882 30658
rect 30882 30606 30884 30658
rect 30828 30604 30884 30606
rect 30044 29036 30100 29092
rect 31388 30156 31444 30212
rect 30156 28754 30212 28756
rect 30156 28702 30158 28754
rect 30158 28702 30210 28754
rect 30210 28702 30212 28754
rect 30156 28700 30212 28702
rect 30716 28924 30772 28980
rect 30380 28812 30436 28868
rect 29932 26012 29988 26068
rect 32172 33516 32228 33572
rect 31948 32898 32004 32900
rect 31948 32846 31950 32898
rect 31950 32846 32002 32898
rect 32002 32846 32004 32898
rect 31948 32844 32004 32846
rect 31836 32060 31892 32116
rect 31836 31890 31892 31892
rect 31836 31838 31838 31890
rect 31838 31838 31890 31890
rect 31890 31838 31892 31890
rect 31836 31836 31892 31838
rect 31276 29484 31332 29540
rect 31612 29596 31668 29652
rect 31276 29036 31332 29092
rect 31052 28588 31108 28644
rect 30828 27970 30884 27972
rect 30828 27918 30830 27970
rect 30830 27918 30882 27970
rect 30882 27918 30884 27970
rect 30828 27916 30884 27918
rect 30604 26738 30660 26740
rect 30604 26686 30606 26738
rect 30606 26686 30658 26738
rect 30658 26686 30660 26738
rect 30604 26684 30660 26686
rect 30156 26124 30212 26180
rect 30604 26236 30660 26292
rect 30156 25506 30212 25508
rect 30156 25454 30158 25506
rect 30158 25454 30210 25506
rect 30210 25454 30212 25506
rect 30156 25452 30212 25454
rect 30828 25842 30884 25844
rect 30828 25790 30830 25842
rect 30830 25790 30882 25842
rect 30882 25790 30884 25842
rect 30828 25788 30884 25790
rect 30716 25004 30772 25060
rect 30044 24892 30100 24948
rect 30828 24946 30884 24948
rect 30828 24894 30830 24946
rect 30830 24894 30882 24946
rect 30882 24894 30884 24946
rect 30828 24892 30884 24894
rect 31836 29596 31892 29652
rect 31724 29036 31780 29092
rect 31500 28866 31556 28868
rect 31500 28814 31502 28866
rect 31502 28814 31554 28866
rect 31554 28814 31556 28866
rect 31500 28812 31556 28814
rect 31836 28364 31892 28420
rect 31500 27580 31556 27636
rect 31612 26796 31668 26852
rect 31388 26460 31444 26516
rect 31388 25900 31444 25956
rect 31724 26572 31780 26628
rect 32508 34524 32564 34580
rect 32396 33794 32452 33796
rect 32396 33742 32398 33794
rect 32398 33742 32450 33794
rect 32450 33742 32452 33794
rect 32396 33740 32452 33742
rect 32508 33458 32564 33460
rect 32508 33406 32510 33458
rect 32510 33406 32562 33458
rect 32562 33406 32564 33458
rect 32508 33404 32564 33406
rect 35196 39338 35252 39340
rect 35196 39286 35198 39338
rect 35198 39286 35250 39338
rect 35250 39286 35252 39338
rect 35196 39284 35252 39286
rect 35300 39338 35356 39340
rect 35300 39286 35302 39338
rect 35302 39286 35354 39338
rect 35354 39286 35356 39338
rect 35300 39284 35356 39286
rect 35404 39338 35460 39340
rect 35404 39286 35406 39338
rect 35406 39286 35458 39338
rect 35458 39286 35460 39338
rect 35404 39284 35460 39286
rect 34524 38444 34580 38500
rect 34748 38892 34804 38948
rect 34636 35586 34692 35588
rect 34636 35534 34638 35586
rect 34638 35534 34690 35586
rect 34690 35534 34692 35586
rect 34636 35532 34692 35534
rect 32732 34748 32788 34804
rect 32732 34578 32788 34580
rect 32732 34526 32734 34578
rect 32734 34526 32786 34578
rect 32786 34526 32788 34578
rect 32732 34524 32788 34526
rect 33404 34524 33460 34580
rect 33180 33852 33236 33908
rect 32732 33740 32788 33796
rect 33516 33794 33572 33796
rect 33516 33742 33518 33794
rect 33518 33742 33570 33794
rect 33570 33742 33572 33794
rect 33516 33740 33572 33742
rect 34076 33628 34132 33684
rect 32620 32172 32676 32228
rect 32060 30658 32116 30660
rect 32060 30606 32062 30658
rect 32062 30606 32114 30658
rect 32114 30606 32116 30658
rect 32060 30604 32116 30606
rect 32732 31612 32788 31668
rect 33068 32172 33124 32228
rect 32620 30044 32676 30100
rect 32172 29596 32228 29652
rect 32172 29260 32228 29316
rect 32620 28812 32676 28868
rect 33292 33404 33348 33460
rect 34188 33404 34244 33460
rect 33628 31724 33684 31780
rect 32956 30492 33012 30548
rect 33628 30492 33684 30548
rect 33516 29820 33572 29876
rect 33180 29762 33236 29764
rect 33180 29710 33182 29762
rect 33182 29710 33234 29762
rect 33234 29710 33236 29762
rect 33180 29708 33236 29710
rect 33292 28924 33348 28980
rect 32956 28754 33012 28756
rect 32956 28702 32958 28754
rect 32958 28702 33010 28754
rect 33010 28702 33012 28754
rect 32956 28700 33012 28702
rect 32620 28476 32676 28532
rect 32172 27692 32228 27748
rect 32620 27804 32676 27860
rect 31948 26684 32004 26740
rect 32284 26796 32340 26852
rect 32508 26738 32564 26740
rect 32508 26686 32510 26738
rect 32510 26686 32562 26738
rect 32562 26686 32564 26738
rect 32508 26684 32564 26686
rect 32060 26514 32116 26516
rect 32060 26462 32062 26514
rect 32062 26462 32114 26514
rect 32114 26462 32116 26514
rect 32060 26460 32116 26462
rect 31724 26236 31780 26292
rect 32508 26236 32564 26292
rect 33180 27468 33236 27524
rect 31164 25618 31220 25620
rect 31164 25566 31166 25618
rect 31166 25566 31218 25618
rect 31218 25566 31220 25618
rect 31164 25564 31220 25566
rect 29596 24444 29652 24500
rect 29820 24332 29876 24388
rect 29372 23996 29428 24052
rect 28140 21756 28196 21812
rect 28700 21810 28756 21812
rect 28700 21758 28702 21810
rect 28702 21758 28754 21810
rect 28754 21758 28756 21810
rect 28700 21756 28756 21758
rect 28588 21644 28644 21700
rect 28588 21196 28644 21252
rect 28476 20412 28532 20468
rect 30268 24610 30324 24612
rect 30268 24558 30270 24610
rect 30270 24558 30322 24610
rect 30322 24558 30324 24610
rect 30268 24556 30324 24558
rect 30604 24498 30660 24500
rect 30604 24446 30606 24498
rect 30606 24446 30658 24498
rect 30658 24446 30660 24498
rect 30604 24444 30660 24446
rect 30044 22540 30100 22596
rect 29820 20860 29876 20916
rect 30604 24050 30660 24052
rect 30604 23998 30606 24050
rect 30606 23998 30658 24050
rect 30658 23998 30660 24050
rect 30604 23996 30660 23998
rect 30716 23436 30772 23492
rect 30156 22482 30212 22484
rect 30156 22430 30158 22482
rect 30158 22430 30210 22482
rect 30210 22430 30212 22482
rect 30156 22428 30212 22430
rect 30716 22316 30772 22372
rect 31164 23884 31220 23940
rect 31164 22764 31220 22820
rect 29148 20300 29204 20356
rect 29484 20466 29540 20468
rect 29484 20414 29486 20466
rect 29486 20414 29538 20466
rect 29538 20414 29540 20466
rect 29484 20412 29540 20414
rect 28028 18732 28084 18788
rect 28588 18786 28644 18788
rect 28588 18734 28590 18786
rect 28590 18734 28642 18786
rect 28642 18734 28644 18786
rect 28588 18732 28644 18734
rect 29260 19852 29316 19908
rect 31500 24498 31556 24500
rect 31500 24446 31502 24498
rect 31502 24446 31554 24498
rect 31554 24446 31556 24498
rect 31500 24444 31556 24446
rect 31388 23938 31444 23940
rect 31388 23886 31390 23938
rect 31390 23886 31442 23938
rect 31442 23886 31444 23938
rect 31388 23884 31444 23886
rect 31724 25730 31780 25732
rect 31724 25678 31726 25730
rect 31726 25678 31778 25730
rect 31778 25678 31780 25730
rect 31724 25676 31780 25678
rect 32172 25730 32228 25732
rect 32172 25678 32174 25730
rect 32174 25678 32226 25730
rect 32226 25678 32228 25730
rect 32172 25676 32228 25678
rect 32620 25676 32676 25732
rect 32060 25452 32116 25508
rect 31724 23772 31780 23828
rect 31500 23548 31556 23604
rect 31164 22594 31220 22596
rect 31164 22542 31166 22594
rect 31166 22542 31218 22594
rect 31218 22542 31220 22594
rect 31164 22540 31220 22542
rect 31948 24610 32004 24612
rect 31948 24558 31950 24610
rect 31950 24558 32002 24610
rect 32002 24558 32004 24610
rect 31948 24556 32004 24558
rect 32060 23660 32116 23716
rect 31948 23548 32004 23604
rect 32508 23436 32564 23492
rect 31612 22540 31668 22596
rect 32284 22482 32340 22484
rect 32284 22430 32286 22482
rect 32286 22430 32338 22482
rect 32338 22430 32340 22482
rect 32284 22428 32340 22430
rect 31836 22316 31892 22372
rect 31052 21756 31108 21812
rect 30268 21698 30324 21700
rect 30268 21646 30270 21698
rect 30270 21646 30322 21698
rect 30322 21646 30324 21698
rect 30268 21644 30324 21646
rect 30268 20914 30324 20916
rect 30268 20862 30270 20914
rect 30270 20862 30322 20914
rect 30322 20862 30324 20914
rect 30268 20860 30324 20862
rect 29820 20300 29876 20356
rect 29596 19794 29652 19796
rect 29596 19742 29598 19794
rect 29598 19742 29650 19794
rect 29650 19742 29652 19794
rect 29596 19740 29652 19742
rect 30380 20412 30436 20468
rect 30492 20636 30548 20692
rect 30380 19852 30436 19908
rect 30268 19628 30324 19684
rect 29596 19180 29652 19236
rect 29484 18732 29540 18788
rect 29932 19180 29988 19236
rect 28812 18284 28868 18340
rect 28028 16604 28084 16660
rect 28028 16268 28084 16324
rect 28812 16828 28868 16884
rect 29820 18396 29876 18452
rect 29260 16716 29316 16772
rect 29372 16828 29428 16884
rect 28364 15372 28420 15428
rect 28140 14418 28196 14420
rect 28140 14366 28142 14418
rect 28142 14366 28194 14418
rect 28194 14366 28196 14418
rect 28140 14364 28196 14366
rect 28140 13634 28196 13636
rect 28140 13582 28142 13634
rect 28142 13582 28194 13634
rect 28194 13582 28196 13634
rect 28140 13580 28196 13582
rect 28028 13356 28084 13412
rect 28028 11788 28084 11844
rect 28476 15260 28532 15316
rect 28812 14812 28868 14868
rect 30828 20690 30884 20692
rect 30828 20638 30830 20690
rect 30830 20638 30882 20690
rect 30882 20638 30884 20690
rect 30828 20636 30884 20638
rect 30828 20412 30884 20468
rect 31276 20412 31332 20468
rect 31052 19682 31108 19684
rect 31052 19630 31054 19682
rect 31054 19630 31106 19682
rect 31106 19630 31108 19682
rect 31052 19628 31108 19630
rect 33516 28924 33572 28980
rect 33516 28140 33572 28196
rect 33516 27858 33572 27860
rect 33516 27806 33518 27858
rect 33518 27806 33570 27858
rect 33570 27806 33572 27858
rect 33516 27804 33572 27806
rect 33740 29762 33796 29764
rect 33740 29710 33742 29762
rect 33742 29710 33794 29762
rect 33794 29710 33796 29762
rect 33740 29708 33796 29710
rect 34188 29820 34244 29876
rect 34076 28642 34132 28644
rect 34076 28590 34078 28642
rect 34078 28590 34130 28642
rect 34130 28590 34132 28642
rect 34076 28588 34132 28590
rect 36092 38892 36148 38948
rect 36988 39564 37044 39620
rect 37548 41580 37604 41636
rect 38668 41692 38724 41748
rect 39004 43820 39060 43876
rect 40012 43820 40068 43876
rect 41692 49026 41748 49028
rect 41692 48974 41694 49026
rect 41694 48974 41746 49026
rect 41746 48974 41748 49026
rect 41692 48972 41748 48974
rect 42364 48972 42420 49028
rect 41804 48860 41860 48916
rect 42140 48860 42196 48916
rect 41356 48748 41412 48804
rect 43484 48860 43540 48916
rect 42812 48748 42868 48804
rect 41244 46620 41300 46676
rect 41580 46620 41636 46676
rect 43708 48860 43764 48916
rect 41468 45276 41524 45332
rect 41132 44658 41188 44660
rect 41132 44606 41134 44658
rect 41134 44606 41186 44658
rect 41186 44606 41188 44658
rect 41132 44604 41188 44606
rect 41244 43874 41300 43876
rect 41244 43822 41246 43874
rect 41246 43822 41298 43874
rect 41298 43822 41300 43874
rect 41244 43820 41300 43822
rect 40012 41804 40068 41860
rect 37884 40908 37940 40964
rect 37660 40460 37716 40516
rect 37884 39676 37940 39732
rect 35308 37660 35364 37716
rect 35196 37322 35252 37324
rect 35196 37270 35198 37322
rect 35198 37270 35250 37322
rect 35250 37270 35252 37322
rect 35196 37268 35252 37270
rect 35300 37322 35356 37324
rect 35300 37270 35302 37322
rect 35302 37270 35354 37322
rect 35354 37270 35356 37322
rect 35300 37268 35356 37270
rect 35404 37322 35460 37324
rect 35404 37270 35406 37322
rect 35406 37270 35458 37322
rect 35458 37270 35460 37322
rect 35404 37268 35460 37270
rect 37548 38892 37604 38948
rect 36428 36594 36484 36596
rect 36428 36542 36430 36594
rect 36430 36542 36482 36594
rect 36482 36542 36484 36594
rect 36428 36540 36484 36542
rect 34972 35810 35028 35812
rect 34972 35758 34974 35810
rect 34974 35758 35026 35810
rect 35026 35758 35028 35810
rect 34972 35756 35028 35758
rect 36428 36092 36484 36148
rect 36876 36092 36932 36148
rect 35980 35532 36036 35588
rect 36204 35756 36260 35812
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34412 34524 34468 34580
rect 35644 34914 35700 34916
rect 35644 34862 35646 34914
rect 35646 34862 35698 34914
rect 35698 34862 35700 34914
rect 35644 34860 35700 34862
rect 36092 34802 36148 34804
rect 36092 34750 36094 34802
rect 36094 34750 36146 34802
rect 36146 34750 36148 34802
rect 36092 34748 36148 34750
rect 35196 34690 35252 34692
rect 35196 34638 35198 34690
rect 35198 34638 35250 34690
rect 35250 34638 35252 34690
rect 35196 34636 35252 34638
rect 35196 33964 35252 34020
rect 34972 33852 35028 33908
rect 34860 33794 34916 33796
rect 34860 33742 34862 33794
rect 34862 33742 34914 33794
rect 34914 33742 34916 33794
rect 34860 33740 34916 33742
rect 34748 33404 34804 33460
rect 34748 31778 34804 31780
rect 34748 31726 34750 31778
rect 34750 31726 34802 31778
rect 34802 31726 34804 31778
rect 34748 31724 34804 31726
rect 34412 30658 34468 30660
rect 34412 30606 34414 30658
rect 34414 30606 34466 30658
rect 34466 30606 34468 30658
rect 34412 30604 34468 30606
rect 34860 30156 34916 30212
rect 34524 29596 34580 29652
rect 34636 29260 34692 29316
rect 34860 29484 34916 29540
rect 34524 28924 34580 28980
rect 33852 27858 33908 27860
rect 33852 27806 33854 27858
rect 33854 27806 33906 27858
rect 33906 27806 33908 27858
rect 33852 27804 33908 27806
rect 33628 27132 33684 27188
rect 34188 27692 34244 27748
rect 33292 26684 33348 26740
rect 32956 26460 33012 26516
rect 33852 26514 33908 26516
rect 33852 26462 33854 26514
rect 33854 26462 33906 26514
rect 33906 26462 33908 26514
rect 33852 26460 33908 26462
rect 33516 26236 33572 26292
rect 32844 25564 32900 25620
rect 33180 23772 33236 23828
rect 33404 25564 33460 25620
rect 33068 23714 33124 23716
rect 33068 23662 33070 23714
rect 33070 23662 33122 23714
rect 33122 23662 33124 23714
rect 33068 23660 33124 23662
rect 33852 25676 33908 25732
rect 32844 23436 32900 23492
rect 33628 24332 33684 24388
rect 33516 23548 33572 23604
rect 32620 22316 32676 22372
rect 32284 20636 32340 20692
rect 31836 20300 31892 20356
rect 33068 20690 33124 20692
rect 33068 20638 33070 20690
rect 33070 20638 33122 20690
rect 33122 20638 33124 20690
rect 33068 20636 33124 20638
rect 33516 20466 33572 20468
rect 33516 20414 33518 20466
rect 33518 20414 33570 20466
rect 33570 20414 33572 20466
rect 33516 20412 33572 20414
rect 32060 19740 32116 19796
rect 32844 19740 32900 19796
rect 31724 19628 31780 19684
rect 30828 17836 30884 17892
rect 30492 16604 30548 16660
rect 29484 15148 29540 15204
rect 29708 14812 29764 14868
rect 29260 14364 29316 14420
rect 29260 13858 29316 13860
rect 29260 13806 29262 13858
rect 29262 13806 29314 13858
rect 29314 13806 29316 13858
rect 29260 13804 29316 13806
rect 32284 19682 32340 19684
rect 32284 19630 32286 19682
rect 32286 19630 32338 19682
rect 32338 19630 32340 19682
rect 32284 19628 32340 19630
rect 30604 15036 30660 15092
rect 30604 14812 30660 14868
rect 28588 13468 28644 13524
rect 28812 13580 28868 13636
rect 31276 15148 31332 15204
rect 31836 15036 31892 15092
rect 30380 13804 30436 13860
rect 30044 13580 30100 13636
rect 28364 12908 28420 12964
rect 28140 10722 28196 10724
rect 28140 10670 28142 10722
rect 28142 10670 28194 10722
rect 28194 10670 28196 10722
rect 28140 10668 28196 10670
rect 30156 13522 30212 13524
rect 30156 13470 30158 13522
rect 30158 13470 30210 13522
rect 30210 13470 30212 13522
rect 30156 13468 30212 13470
rect 31836 14476 31892 14532
rect 32284 15148 32340 15204
rect 33404 20076 33460 20132
rect 33964 22818 34020 22820
rect 33964 22766 33966 22818
rect 33966 22766 34018 22818
rect 34018 22766 34020 22818
rect 33964 22764 34020 22766
rect 34188 26626 34244 26628
rect 34188 26574 34190 26626
rect 34190 26574 34242 26626
rect 34242 26574 34244 26626
rect 34188 26572 34244 26574
rect 34636 28028 34692 28084
rect 34524 27804 34580 27860
rect 35868 33964 35924 34020
rect 36764 35810 36820 35812
rect 36764 35758 36766 35810
rect 36766 35758 36818 35810
rect 36818 35758 36820 35810
rect 36764 35756 36820 35758
rect 37324 35810 37380 35812
rect 37324 35758 37326 35810
rect 37326 35758 37378 35810
rect 37378 35758 37380 35810
rect 37324 35756 37380 35758
rect 35644 33740 35700 33796
rect 35532 33682 35588 33684
rect 35532 33630 35534 33682
rect 35534 33630 35586 33682
rect 35586 33630 35588 33682
rect 35532 33628 35588 33630
rect 35196 33290 35252 33292
rect 35196 33238 35198 33290
rect 35198 33238 35250 33290
rect 35250 33238 35252 33290
rect 35196 33236 35252 33238
rect 35300 33290 35356 33292
rect 35300 33238 35302 33290
rect 35302 33238 35354 33290
rect 35354 33238 35356 33290
rect 35300 33236 35356 33238
rect 35404 33290 35460 33292
rect 35404 33238 35406 33290
rect 35406 33238 35458 33290
rect 35458 33238 35460 33290
rect 35404 33236 35460 33238
rect 35756 33404 35812 33460
rect 35644 31836 35700 31892
rect 35532 31724 35588 31780
rect 35196 31274 35252 31276
rect 35196 31222 35198 31274
rect 35198 31222 35250 31274
rect 35250 31222 35252 31274
rect 35196 31220 35252 31222
rect 35300 31274 35356 31276
rect 35300 31222 35302 31274
rect 35302 31222 35354 31274
rect 35354 31222 35356 31274
rect 35300 31220 35356 31222
rect 35404 31274 35460 31276
rect 35404 31222 35406 31274
rect 35406 31222 35458 31274
rect 35458 31222 35460 31274
rect 35404 31220 35460 31222
rect 35756 31724 35812 31780
rect 38892 41580 38948 41636
rect 38556 40684 38612 40740
rect 38108 38946 38164 38948
rect 38108 38894 38110 38946
rect 38110 38894 38162 38946
rect 38162 38894 38164 38946
rect 38108 38892 38164 38894
rect 38220 39676 38276 39732
rect 37884 38668 37940 38724
rect 37772 38220 37828 38276
rect 37884 37996 37940 38052
rect 37660 36540 37716 36596
rect 37548 34860 37604 34916
rect 37660 34748 37716 34804
rect 38556 38220 38612 38276
rect 37884 34636 37940 34692
rect 36988 34018 37044 34020
rect 36988 33966 36990 34018
rect 36990 33966 37042 34018
rect 37042 33966 37044 34018
rect 36988 33964 37044 33966
rect 37324 32956 37380 33012
rect 37996 33404 38052 33460
rect 38108 32956 38164 33012
rect 37772 31890 37828 31892
rect 37772 31838 37774 31890
rect 37774 31838 37826 31890
rect 37826 31838 37828 31890
rect 37772 31836 37828 31838
rect 36540 31388 36596 31444
rect 35532 30492 35588 30548
rect 35532 30044 35588 30100
rect 35420 29762 35476 29764
rect 35420 29710 35422 29762
rect 35422 29710 35474 29762
rect 35474 29710 35476 29762
rect 35420 29708 35476 29710
rect 35196 29538 35252 29540
rect 35196 29486 35198 29538
rect 35198 29486 35250 29538
rect 35250 29486 35252 29538
rect 35196 29484 35252 29486
rect 35196 29258 35252 29260
rect 35196 29206 35198 29258
rect 35198 29206 35250 29258
rect 35250 29206 35252 29258
rect 35196 29204 35252 29206
rect 35300 29258 35356 29260
rect 35300 29206 35302 29258
rect 35302 29206 35354 29258
rect 35354 29206 35356 29258
rect 35300 29204 35356 29206
rect 35404 29258 35460 29260
rect 35404 29206 35406 29258
rect 35406 29206 35458 29258
rect 35458 29206 35460 29258
rect 35404 29204 35460 29206
rect 35756 30716 35812 30772
rect 35980 30268 36036 30324
rect 35196 28140 35252 28196
rect 35532 28082 35588 28084
rect 35532 28030 35534 28082
rect 35534 28030 35586 28082
rect 35586 28030 35588 28082
rect 35532 28028 35588 28030
rect 34188 23826 34244 23828
rect 34188 23774 34190 23826
rect 34190 23774 34242 23826
rect 34242 23774 34244 23826
rect 34188 23772 34244 23774
rect 34412 25954 34468 25956
rect 34412 25902 34414 25954
rect 34414 25902 34466 25954
rect 34466 25902 34468 25954
rect 34412 25900 34468 25902
rect 35084 27746 35140 27748
rect 35084 27694 35086 27746
rect 35086 27694 35138 27746
rect 35138 27694 35140 27746
rect 35084 27692 35140 27694
rect 35084 27468 35140 27524
rect 35196 27242 35252 27244
rect 35196 27190 35198 27242
rect 35198 27190 35250 27242
rect 35250 27190 35252 27242
rect 35196 27188 35252 27190
rect 35300 27242 35356 27244
rect 35300 27190 35302 27242
rect 35302 27190 35354 27242
rect 35354 27190 35356 27242
rect 35300 27188 35356 27190
rect 35404 27242 35460 27244
rect 35404 27190 35406 27242
rect 35406 27190 35458 27242
rect 35458 27190 35460 27242
rect 35404 27188 35460 27190
rect 35644 27746 35700 27748
rect 35644 27694 35646 27746
rect 35646 27694 35698 27746
rect 35698 27694 35700 27746
rect 35644 27692 35700 27694
rect 35532 26796 35588 26852
rect 35868 26684 35924 26740
rect 35196 26514 35252 26516
rect 35196 26462 35198 26514
rect 35198 26462 35250 26514
rect 35250 26462 35252 26514
rect 35196 26460 35252 26462
rect 35868 26514 35924 26516
rect 35868 26462 35870 26514
rect 35870 26462 35922 26514
rect 35922 26462 35924 26514
rect 35868 26460 35924 26462
rect 36988 31778 37044 31780
rect 36988 31726 36990 31778
rect 36990 31726 37042 31778
rect 37042 31726 37044 31778
rect 36988 31724 37044 31726
rect 37324 30716 37380 30772
rect 36652 30268 36708 30324
rect 36540 30156 36596 30212
rect 36204 29874 36260 29876
rect 36204 29822 36206 29874
rect 36206 29822 36258 29874
rect 36258 29822 36260 29874
rect 36204 29820 36260 29822
rect 36988 29820 37044 29876
rect 36092 28924 36148 28980
rect 35532 25900 35588 25956
rect 34972 25618 35028 25620
rect 34972 25566 34974 25618
rect 34974 25566 35026 25618
rect 35026 25566 35028 25618
rect 34972 25564 35028 25566
rect 34972 25340 35028 25396
rect 35644 25618 35700 25620
rect 35644 25566 35646 25618
rect 35646 25566 35698 25618
rect 35698 25566 35700 25618
rect 35644 25564 35700 25566
rect 35196 25226 35252 25228
rect 35196 25174 35198 25226
rect 35198 25174 35250 25226
rect 35250 25174 35252 25226
rect 35196 25172 35252 25174
rect 35300 25226 35356 25228
rect 35300 25174 35302 25226
rect 35302 25174 35354 25226
rect 35354 25174 35356 25226
rect 35300 25172 35356 25174
rect 35404 25226 35460 25228
rect 35404 25174 35406 25226
rect 35406 25174 35458 25226
rect 35458 25174 35460 25226
rect 35404 25172 35460 25174
rect 34748 24556 34804 24612
rect 35532 24498 35588 24500
rect 35532 24446 35534 24498
rect 35534 24446 35586 24498
rect 35586 24446 35588 24498
rect 35532 24444 35588 24446
rect 34636 23602 34692 23604
rect 34636 23550 34638 23602
rect 34638 23550 34690 23602
rect 34690 23550 34692 23602
rect 34636 23548 34692 23550
rect 34412 21810 34468 21812
rect 34412 21758 34414 21810
rect 34414 21758 34466 21810
rect 34466 21758 34468 21810
rect 34412 21756 34468 21758
rect 34076 21586 34132 21588
rect 34076 21534 34078 21586
rect 34078 21534 34130 21586
rect 34130 21534 34132 21586
rect 34076 21532 34132 21534
rect 35868 25452 35924 25508
rect 37100 29650 37156 29652
rect 37100 29598 37102 29650
rect 37102 29598 37154 29650
rect 37154 29598 37156 29650
rect 37100 29596 37156 29598
rect 37660 31388 37716 31444
rect 38444 30492 38500 30548
rect 37996 30268 38052 30324
rect 37212 29484 37268 29540
rect 37548 29484 37604 29540
rect 38332 28588 38388 28644
rect 36092 25452 36148 25508
rect 36540 26572 36596 26628
rect 37660 26572 37716 26628
rect 36428 25676 36484 25732
rect 36876 25676 36932 25732
rect 36204 25340 36260 25396
rect 36652 24780 36708 24836
rect 35980 24498 36036 24500
rect 35980 24446 35982 24498
rect 35982 24446 36034 24498
rect 36034 24446 36036 24498
rect 35980 24444 36036 24446
rect 35532 23548 35588 23604
rect 35196 23210 35252 23212
rect 35196 23158 35198 23210
rect 35198 23158 35250 23210
rect 35250 23158 35252 23210
rect 35196 23156 35252 23158
rect 35300 23210 35356 23212
rect 35300 23158 35302 23210
rect 35302 23158 35354 23210
rect 35354 23158 35356 23210
rect 35300 23156 35356 23158
rect 35404 23210 35460 23212
rect 35404 23158 35406 23210
rect 35406 23158 35458 23210
rect 35458 23158 35460 23210
rect 35404 23156 35460 23158
rect 35532 22764 35588 22820
rect 34972 21810 35028 21812
rect 34972 21758 34974 21810
rect 34974 21758 35026 21810
rect 35026 21758 35028 21810
rect 34972 21756 35028 21758
rect 33852 20300 33908 20356
rect 35084 21420 35140 21476
rect 33964 20076 34020 20132
rect 34300 20636 34356 20692
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 21026 35252 21028
rect 35196 20974 35198 21026
rect 35198 20974 35250 21026
rect 35250 20974 35252 21026
rect 35196 20972 35252 20974
rect 35196 20300 35252 20356
rect 35196 19178 35252 19180
rect 35196 19126 35198 19178
rect 35198 19126 35250 19178
rect 35250 19126 35252 19178
rect 35196 19124 35252 19126
rect 35300 19178 35356 19180
rect 35300 19126 35302 19178
rect 35302 19126 35354 19178
rect 35354 19126 35356 19178
rect 35300 19124 35356 19126
rect 35404 19178 35460 19180
rect 35404 19126 35406 19178
rect 35406 19126 35458 19178
rect 35458 19126 35460 19178
rect 35404 19124 35460 19126
rect 37548 25730 37604 25732
rect 37548 25678 37550 25730
rect 37550 25678 37602 25730
rect 37602 25678 37604 25730
rect 37548 25676 37604 25678
rect 37436 25564 37492 25620
rect 37772 25564 37828 25620
rect 38220 26684 38276 26740
rect 37548 25452 37604 25508
rect 36876 24444 36932 24500
rect 36204 22818 36260 22820
rect 36204 22766 36206 22818
rect 36206 22766 36258 22818
rect 36258 22766 36260 22818
rect 36204 22764 36260 22766
rect 36428 23602 36484 23604
rect 36428 23550 36430 23602
rect 36430 23550 36482 23602
rect 36482 23550 36484 23602
rect 36428 23548 36484 23550
rect 37996 26236 38052 26292
rect 37996 25676 38052 25732
rect 37884 24780 37940 24836
rect 35980 21868 36036 21924
rect 35644 21810 35700 21812
rect 35644 21758 35646 21810
rect 35646 21758 35698 21810
rect 35698 21758 35700 21810
rect 35644 21756 35700 21758
rect 36204 21474 36260 21476
rect 36204 21422 36206 21474
rect 36206 21422 36258 21474
rect 36258 21422 36260 21474
rect 36204 21420 36260 21422
rect 37996 22540 38052 22596
rect 37100 21756 37156 21812
rect 36316 20802 36372 20804
rect 36316 20750 36318 20802
rect 36318 20750 36370 20802
rect 36370 20750 36372 20802
rect 36316 20748 36372 20750
rect 35644 19292 35700 19348
rect 35980 18674 36036 18676
rect 35980 18622 35982 18674
rect 35982 18622 36034 18674
rect 36034 18622 36036 18674
rect 35980 18620 36036 18622
rect 37212 20802 37268 20804
rect 37212 20750 37214 20802
rect 37214 20750 37266 20802
rect 37266 20750 37268 20802
rect 37212 20748 37268 20750
rect 39900 41746 39956 41748
rect 39900 41694 39902 41746
rect 39902 41694 39954 41746
rect 39954 41694 39956 41746
rect 39900 41692 39956 41694
rect 39228 39058 39284 39060
rect 39228 39006 39230 39058
rect 39230 39006 39282 39058
rect 39282 39006 39284 39058
rect 39228 39004 39284 39006
rect 38892 38722 38948 38724
rect 38892 38670 38894 38722
rect 38894 38670 38946 38722
rect 38946 38670 38948 38722
rect 38892 38668 38948 38670
rect 40348 40908 40404 40964
rect 39900 40066 39956 40068
rect 39900 40014 39902 40066
rect 39902 40014 39954 40066
rect 39954 40014 39956 40066
rect 39900 40012 39956 40014
rect 40460 39004 40516 39060
rect 38892 35980 38948 36036
rect 40348 37996 40404 38052
rect 39228 35810 39284 35812
rect 39228 35758 39230 35810
rect 39230 35758 39282 35810
rect 39282 35758 39284 35810
rect 39228 35756 39284 35758
rect 38780 34076 38836 34132
rect 39228 34018 39284 34020
rect 39228 33966 39230 34018
rect 39230 33966 39282 34018
rect 39282 33966 39284 34018
rect 39228 33964 39284 33966
rect 38668 33628 38724 33684
rect 39116 33404 39172 33460
rect 39788 37772 39844 37828
rect 40348 37548 40404 37604
rect 41132 41916 41188 41972
rect 40908 41858 40964 41860
rect 40908 41806 40910 41858
rect 40910 41806 40962 41858
rect 40962 41806 40964 41858
rect 40908 41804 40964 41806
rect 41580 41580 41636 41636
rect 41244 40738 41300 40740
rect 41244 40686 41246 40738
rect 41246 40686 41298 40738
rect 41298 40686 41300 40738
rect 41244 40684 41300 40686
rect 40908 40012 40964 40068
rect 42924 45276 42980 45332
rect 43036 46508 43092 46564
rect 50556 48410 50612 48412
rect 50556 48358 50558 48410
rect 50558 48358 50610 48410
rect 50610 48358 50612 48410
rect 50556 48356 50612 48358
rect 50660 48410 50716 48412
rect 50660 48358 50662 48410
rect 50662 48358 50714 48410
rect 50714 48358 50716 48410
rect 50660 48356 50716 48358
rect 50764 48410 50820 48412
rect 50764 48358 50766 48410
rect 50766 48358 50818 48410
rect 50818 48358 50820 48410
rect 50764 48356 50820 48358
rect 44044 46562 44100 46564
rect 44044 46510 44046 46562
rect 44046 46510 44098 46562
rect 44098 46510 44100 46562
rect 44044 46508 44100 46510
rect 50556 46394 50612 46396
rect 50556 46342 50558 46394
rect 50558 46342 50610 46394
rect 50610 46342 50612 46394
rect 50556 46340 50612 46342
rect 50660 46394 50716 46396
rect 50660 46342 50662 46394
rect 50662 46342 50714 46394
rect 50714 46342 50716 46394
rect 50660 46340 50716 46342
rect 50764 46394 50820 46396
rect 50764 46342 50766 46394
rect 50766 46342 50818 46394
rect 50818 46342 50820 46394
rect 50764 46340 50820 46342
rect 45164 44658 45220 44660
rect 45164 44606 45166 44658
rect 45166 44606 45218 44658
rect 45218 44606 45220 44658
rect 45164 44604 45220 44606
rect 43148 43708 43204 43764
rect 42588 41916 42644 41972
rect 42364 40012 42420 40068
rect 41356 39004 41412 39060
rect 41132 38892 41188 38948
rect 41244 38668 41300 38724
rect 40908 37826 40964 37828
rect 40908 37774 40910 37826
rect 40910 37774 40962 37826
rect 40962 37774 40964 37826
rect 40908 37772 40964 37774
rect 39676 35980 39732 36036
rect 39340 33516 39396 33572
rect 39452 34860 39508 34916
rect 39228 32956 39284 33012
rect 39116 32898 39172 32900
rect 39116 32846 39118 32898
rect 39118 32846 39170 32898
rect 39170 32846 39172 32898
rect 39116 32844 39172 32846
rect 39228 32620 39284 32676
rect 39228 30716 39284 30772
rect 39676 32620 39732 32676
rect 40348 36092 40404 36148
rect 40348 35698 40404 35700
rect 40348 35646 40350 35698
rect 40350 35646 40402 35698
rect 40402 35646 40404 35698
rect 40348 35644 40404 35646
rect 40796 34636 40852 34692
rect 40348 34188 40404 34244
rect 40572 34188 40628 34244
rect 40348 34018 40404 34020
rect 40348 33966 40350 34018
rect 40350 33966 40402 34018
rect 40402 33966 40404 34018
rect 40348 33964 40404 33966
rect 40124 32674 40180 32676
rect 40124 32622 40126 32674
rect 40126 32622 40178 32674
rect 40178 32622 40180 32674
rect 40124 32620 40180 32622
rect 39900 31836 39956 31892
rect 40236 31836 40292 31892
rect 40348 31666 40404 31668
rect 40348 31614 40350 31666
rect 40350 31614 40402 31666
rect 40402 31614 40404 31666
rect 40348 31612 40404 31614
rect 40348 31276 40404 31332
rect 39676 30492 39732 30548
rect 39900 30716 39956 30772
rect 39452 30044 39508 30100
rect 40348 30492 40404 30548
rect 40124 30268 40180 30324
rect 39900 28866 39956 28868
rect 39900 28814 39902 28866
rect 39902 28814 39954 28866
rect 39954 28814 39956 28866
rect 39900 28812 39956 28814
rect 38556 28588 38612 28644
rect 41020 34748 41076 34804
rect 41020 34018 41076 34020
rect 41020 33966 41022 34018
rect 41022 33966 41074 34018
rect 41074 33966 41076 34018
rect 41020 33964 41076 33966
rect 41244 35980 41300 36036
rect 41244 33628 41300 33684
rect 43036 40908 43092 40964
rect 42700 40684 42756 40740
rect 41916 39842 41972 39844
rect 41916 39790 41918 39842
rect 41918 39790 41970 39842
rect 41970 39790 41972 39842
rect 41916 39788 41972 39790
rect 42028 38668 42084 38724
rect 43932 41970 43988 41972
rect 43932 41918 43934 41970
rect 43934 41918 43986 41970
rect 43986 41918 43988 41970
rect 43932 41916 43988 41918
rect 43484 41580 43540 41636
rect 44380 41916 44436 41972
rect 44268 41858 44324 41860
rect 44268 41806 44270 41858
rect 44270 41806 44322 41858
rect 44322 41806 44324 41858
rect 44268 41804 44324 41806
rect 44716 41916 44772 41972
rect 44940 41804 44996 41860
rect 45500 44604 45556 44660
rect 45724 43762 45780 43764
rect 45724 43710 45726 43762
rect 45726 43710 45778 43762
rect 45778 43710 45780 43762
rect 45724 43708 45780 43710
rect 45500 43596 45556 43652
rect 46508 43708 46564 43764
rect 45388 42140 45444 42196
rect 45388 41916 45444 41972
rect 44492 41692 44548 41748
rect 43932 40908 43988 40964
rect 43484 40796 43540 40852
rect 44044 40850 44100 40852
rect 44044 40798 44046 40850
rect 44046 40798 44098 40850
rect 44098 40798 44100 40850
rect 44044 40796 44100 40798
rect 42476 37826 42532 37828
rect 42476 37774 42478 37826
rect 42478 37774 42530 37826
rect 42530 37774 42532 37826
rect 42476 37772 42532 37774
rect 42252 37548 42308 37604
rect 42588 37660 42644 37716
rect 41916 35980 41972 36036
rect 42252 35980 42308 36036
rect 41580 34802 41636 34804
rect 41580 34750 41582 34802
rect 41582 34750 41634 34802
rect 41634 34750 41636 34802
rect 41580 34748 41636 34750
rect 41468 34188 41524 34244
rect 41692 34636 41748 34692
rect 43708 40066 43764 40068
rect 43708 40014 43710 40066
rect 43710 40014 43762 40066
rect 43762 40014 43764 40066
rect 43708 40012 43764 40014
rect 44940 39900 44996 39956
rect 46060 43484 46116 43540
rect 46732 43596 46788 43652
rect 50556 44378 50612 44380
rect 50556 44326 50558 44378
rect 50558 44326 50610 44378
rect 50610 44326 50612 44378
rect 50556 44324 50612 44326
rect 50660 44378 50716 44380
rect 50660 44326 50662 44378
rect 50662 44326 50714 44378
rect 50714 44326 50716 44378
rect 50660 44324 50716 44326
rect 50764 44378 50820 44380
rect 50764 44326 50766 44378
rect 50766 44326 50818 44378
rect 50818 44326 50820 44378
rect 50764 44324 50820 44326
rect 47292 43596 47348 43652
rect 47404 43484 47460 43540
rect 47964 43484 48020 43540
rect 47964 42866 48020 42868
rect 47964 42814 47966 42866
rect 47966 42814 48018 42866
rect 48018 42814 48020 42866
rect 47964 42812 48020 42814
rect 47516 42754 47572 42756
rect 47516 42702 47518 42754
rect 47518 42702 47570 42754
rect 47570 42702 47572 42754
rect 47516 42700 47572 42702
rect 46732 42140 46788 42196
rect 45612 41692 45668 41748
rect 45388 40850 45444 40852
rect 45388 40798 45390 40850
rect 45390 40798 45442 40850
rect 45442 40798 45444 40850
rect 45388 40796 45444 40798
rect 46732 40850 46788 40852
rect 46732 40798 46734 40850
rect 46734 40798 46786 40850
rect 46786 40798 46788 40850
rect 46732 40796 46788 40798
rect 46732 40124 46788 40180
rect 45724 39954 45780 39956
rect 45724 39902 45726 39954
rect 45726 39902 45778 39954
rect 45778 39902 45780 39954
rect 45724 39900 45780 39902
rect 44492 39842 44548 39844
rect 44492 39790 44494 39842
rect 44494 39790 44546 39842
rect 44546 39790 44548 39842
rect 44492 39788 44548 39790
rect 45388 39842 45444 39844
rect 45388 39790 45390 39842
rect 45390 39790 45442 39842
rect 45442 39790 45444 39842
rect 45388 39788 45444 39790
rect 44940 38780 44996 38836
rect 43036 37548 43092 37604
rect 43484 37772 43540 37828
rect 46508 38780 46564 38836
rect 47740 42140 47796 42196
rect 47516 41804 47572 41860
rect 47516 40850 47572 40852
rect 47516 40798 47518 40850
rect 47518 40798 47570 40850
rect 47570 40798 47572 40850
rect 47516 40796 47572 40798
rect 49420 42812 49476 42868
rect 48860 42700 48916 42756
rect 49084 42140 49140 42196
rect 48860 42028 48916 42084
rect 49308 42028 49364 42084
rect 48636 41804 48692 41860
rect 49196 41858 49252 41860
rect 49196 41806 49198 41858
rect 49198 41806 49250 41858
rect 49250 41806 49252 41858
rect 49196 41804 49252 41806
rect 48748 39900 48804 39956
rect 46844 39788 46900 39844
rect 45948 37884 46004 37940
rect 44492 37772 44548 37828
rect 43148 36540 43204 36596
rect 43484 36652 43540 36708
rect 44044 36652 44100 36708
rect 43820 35980 43876 36036
rect 43932 36540 43988 36596
rect 43148 35644 43204 35700
rect 42588 34860 42644 34916
rect 43596 34860 43652 34916
rect 42252 34690 42308 34692
rect 42252 34638 42254 34690
rect 42254 34638 42306 34690
rect 42306 34638 42308 34690
rect 42252 34636 42308 34638
rect 42364 34748 42420 34804
rect 41804 34076 41860 34132
rect 42812 34636 42868 34692
rect 43260 34524 43316 34580
rect 40908 31612 40964 31668
rect 40572 31052 40628 31108
rect 41132 31052 41188 31108
rect 41356 30770 41412 30772
rect 41356 30718 41358 30770
rect 41358 30718 41410 30770
rect 41410 30718 41412 30770
rect 41356 30716 41412 30718
rect 40796 29426 40852 29428
rect 40796 29374 40798 29426
rect 40798 29374 40850 29426
rect 40850 29374 40852 29426
rect 40796 29372 40852 29374
rect 41244 28866 41300 28868
rect 41244 28814 41246 28866
rect 41246 28814 41298 28866
rect 41298 28814 41300 28866
rect 41244 28812 41300 28814
rect 39116 28588 39172 28644
rect 38780 28476 38836 28532
rect 38780 26626 38836 26628
rect 38780 26574 38782 26626
rect 38782 26574 38834 26626
rect 38834 26574 38836 26626
rect 38780 26572 38836 26574
rect 39340 27020 39396 27076
rect 38668 26236 38724 26292
rect 38668 25676 38724 25732
rect 40348 26908 40404 26964
rect 39452 26796 39508 26852
rect 39676 25730 39732 25732
rect 39676 25678 39678 25730
rect 39678 25678 39730 25730
rect 39730 25678 39732 25730
rect 39676 25676 39732 25678
rect 38892 24668 38948 24724
rect 39788 24722 39844 24724
rect 39788 24670 39790 24722
rect 39790 24670 39842 24722
rect 39842 24670 39844 24722
rect 39788 24668 39844 24670
rect 38780 23826 38836 23828
rect 38780 23774 38782 23826
rect 38782 23774 38834 23826
rect 38834 23774 38836 23826
rect 38780 23772 38836 23774
rect 40348 25676 40404 25732
rect 39900 23772 39956 23828
rect 40012 23436 40068 23492
rect 39340 22988 39396 23044
rect 40124 23042 40180 23044
rect 40124 22990 40126 23042
rect 40126 22990 40178 23042
rect 40178 22990 40180 23042
rect 40124 22988 40180 22990
rect 40572 24332 40628 24388
rect 40572 23884 40628 23940
rect 40796 23490 40852 23492
rect 40796 23438 40798 23490
rect 40798 23438 40850 23490
rect 40850 23438 40852 23490
rect 40796 23436 40852 23438
rect 41020 27020 41076 27076
rect 41244 25676 41300 25732
rect 41468 24386 41524 24388
rect 41468 24334 41470 24386
rect 41470 24334 41522 24386
rect 41522 24334 41524 24386
rect 41468 24332 41524 24334
rect 41020 23884 41076 23940
rect 41356 23884 41412 23940
rect 41244 23548 41300 23604
rect 40572 22540 40628 22596
rect 38332 20748 38388 20804
rect 37100 20412 37156 20468
rect 38332 20466 38388 20468
rect 38332 20414 38334 20466
rect 38334 20414 38386 20466
rect 38386 20414 38388 20466
rect 38332 20412 38388 20414
rect 36316 18620 36372 18676
rect 36204 18508 36260 18564
rect 34748 18396 34804 18452
rect 34972 16770 35028 16772
rect 34972 16718 34974 16770
rect 34974 16718 35026 16770
rect 35026 16718 35028 16770
rect 34972 16716 35028 16718
rect 32732 14812 32788 14868
rect 32060 13858 32116 13860
rect 32060 13806 32062 13858
rect 32062 13806 32114 13858
rect 32114 13806 32116 13858
rect 32060 13804 32116 13806
rect 32508 13634 32564 13636
rect 32508 13582 32510 13634
rect 32510 13582 32562 13634
rect 32562 13582 32564 13634
rect 32508 13580 32564 13582
rect 30828 13468 30884 13524
rect 35308 18396 35364 18452
rect 37660 18620 37716 18676
rect 36428 18284 36484 18340
rect 37548 18508 37604 18564
rect 35196 17162 35252 17164
rect 35196 17110 35198 17162
rect 35198 17110 35250 17162
rect 35250 17110 35252 17162
rect 35196 17108 35252 17110
rect 35300 17162 35356 17164
rect 35300 17110 35302 17162
rect 35302 17110 35354 17162
rect 35354 17110 35356 17162
rect 35300 17108 35356 17110
rect 35404 17162 35460 17164
rect 35404 17110 35406 17162
rect 35406 17110 35458 17162
rect 35458 17110 35460 17162
rect 35404 17108 35460 17110
rect 36764 16716 36820 16772
rect 36204 15762 36260 15764
rect 36204 15710 36206 15762
rect 36206 15710 36258 15762
rect 36258 15710 36260 15762
rect 36204 15708 36260 15710
rect 37436 16716 37492 16772
rect 35084 15596 35140 15652
rect 33068 14812 33124 14868
rect 35196 15146 35252 15148
rect 35196 15094 35198 15146
rect 35198 15094 35250 15146
rect 35250 15094 35252 15146
rect 35196 15092 35252 15094
rect 35300 15146 35356 15148
rect 35300 15094 35302 15146
rect 35302 15094 35354 15146
rect 35354 15094 35356 15146
rect 35300 15092 35356 15094
rect 35404 15146 35460 15148
rect 35404 15094 35406 15146
rect 35406 15094 35458 15146
rect 35458 15094 35460 15146
rect 35404 15092 35460 15094
rect 33180 14642 33236 14644
rect 33180 14590 33182 14642
rect 33182 14590 33234 14642
rect 33234 14590 33236 14642
rect 33180 14588 33236 14590
rect 34076 14530 34132 14532
rect 34076 14478 34078 14530
rect 34078 14478 34130 14530
rect 34130 14478 34132 14530
rect 34076 14476 34132 14478
rect 33516 14306 33572 14308
rect 33516 14254 33518 14306
rect 33518 14254 33570 14306
rect 33570 14254 33572 14306
rect 33516 14252 33572 14254
rect 32844 13356 32900 13412
rect 31948 12962 32004 12964
rect 31948 12910 31950 12962
rect 31950 12910 32002 12962
rect 32002 12910 32004 12962
rect 31948 12908 32004 12910
rect 32844 12684 32900 12740
rect 33180 13692 33236 13748
rect 28252 10444 28308 10500
rect 27468 10108 27524 10164
rect 28588 9660 28644 9716
rect 27356 7756 27412 7812
rect 30044 10668 30100 10724
rect 29148 8540 29204 8596
rect 29260 9660 29316 9716
rect 29708 10498 29764 10500
rect 29708 10446 29710 10498
rect 29710 10446 29762 10498
rect 29762 10446 29764 10498
rect 29708 10444 29764 10446
rect 29596 9714 29652 9716
rect 29596 9662 29598 9714
rect 29598 9662 29650 9714
rect 29650 9662 29652 9714
rect 29596 9660 29652 9662
rect 30604 9660 30660 9716
rect 29372 8652 29428 8708
rect 30268 8706 30324 8708
rect 30268 8654 30270 8706
rect 30270 8654 30322 8706
rect 30322 8654 30324 8706
rect 30268 8652 30324 8654
rect 29820 8594 29876 8596
rect 29820 8542 29822 8594
rect 29822 8542 29874 8594
rect 29874 8542 29876 8594
rect 29820 8540 29876 8542
rect 27468 6636 27524 6692
rect 27020 6524 27076 6580
rect 28924 6636 28980 6692
rect 28812 6524 28868 6580
rect 27916 5794 27972 5796
rect 27916 5742 27918 5794
rect 27918 5742 27970 5794
rect 27970 5742 27972 5794
rect 27916 5740 27972 5742
rect 28476 5404 28532 5460
rect 26684 4620 26740 4676
rect 27692 4674 27748 4676
rect 27692 4622 27694 4674
rect 27694 4622 27746 4674
rect 27746 4622 27748 4674
rect 27692 4620 27748 4622
rect 30268 7922 30324 7924
rect 30268 7870 30270 7922
rect 30270 7870 30322 7922
rect 30322 7870 30324 7922
rect 30268 7868 30324 7870
rect 30716 10668 30772 10724
rect 30716 8706 30772 8708
rect 30716 8654 30718 8706
rect 30718 8654 30770 8706
rect 30770 8654 30772 8706
rect 30716 8652 30772 8654
rect 31276 10444 31332 10500
rect 32844 11788 32900 11844
rect 32172 9772 32228 9828
rect 32396 10444 32452 10500
rect 31164 8482 31220 8484
rect 31164 8430 31166 8482
rect 31166 8430 31218 8482
rect 31218 8430 31220 8482
rect 31164 8428 31220 8430
rect 31388 8594 31444 8596
rect 31388 8542 31390 8594
rect 31390 8542 31442 8594
rect 31442 8542 31444 8594
rect 31388 8540 31444 8542
rect 30380 6636 30436 6692
rect 29260 6578 29316 6580
rect 29260 6526 29262 6578
rect 29262 6526 29314 6578
rect 29314 6526 29316 6578
rect 29260 6524 29316 6526
rect 32060 8652 32116 8708
rect 33068 10498 33124 10500
rect 33068 10446 33070 10498
rect 33070 10446 33122 10498
rect 33122 10446 33124 10498
rect 33068 10444 33124 10446
rect 33740 13692 33796 13748
rect 33964 13634 34020 13636
rect 33964 13582 33966 13634
rect 33966 13582 34018 13634
rect 34018 13582 34020 13634
rect 33964 13580 34020 13582
rect 33628 13468 33684 13524
rect 34076 13468 34132 13524
rect 34524 12738 34580 12740
rect 34524 12686 34526 12738
rect 34526 12686 34578 12738
rect 34578 12686 34580 12738
rect 34524 12684 34580 12686
rect 32508 10332 32564 10388
rect 32732 9548 32788 9604
rect 32732 8428 32788 8484
rect 31836 6578 31892 6580
rect 31836 6526 31838 6578
rect 31838 6526 31890 6578
rect 31890 6526 31892 6578
rect 31836 6524 31892 6526
rect 31612 6412 31668 6468
rect 29148 5740 29204 5796
rect 29820 5740 29876 5796
rect 32396 6412 32452 6468
rect 32508 7532 32564 7588
rect 33292 8652 33348 8708
rect 32732 6636 32788 6692
rect 33068 6636 33124 6692
rect 34860 14812 34916 14868
rect 34748 13580 34804 13636
rect 36428 14754 36484 14756
rect 36428 14702 36430 14754
rect 36430 14702 36482 14754
rect 36482 14702 36484 14754
rect 36428 14700 36484 14702
rect 37100 14642 37156 14644
rect 37100 14590 37102 14642
rect 37102 14590 37154 14642
rect 37154 14590 37156 14642
rect 37100 14588 37156 14590
rect 35644 14530 35700 14532
rect 35644 14478 35646 14530
rect 35646 14478 35698 14530
rect 35698 14478 35700 14530
rect 35644 14476 35700 14478
rect 34860 13468 34916 13524
rect 37212 14252 37268 14308
rect 35196 13130 35252 13132
rect 35196 13078 35198 13130
rect 35198 13078 35250 13130
rect 35250 13078 35252 13130
rect 35196 13076 35252 13078
rect 35300 13130 35356 13132
rect 35300 13078 35302 13130
rect 35302 13078 35354 13130
rect 35354 13078 35356 13130
rect 35300 13076 35356 13078
rect 35404 13130 35460 13132
rect 35404 13078 35406 13130
rect 35406 13078 35458 13130
rect 35458 13078 35460 13130
rect 35404 13076 35460 13078
rect 36428 12796 36484 12852
rect 37100 12626 37156 12628
rect 37100 12574 37102 12626
rect 37102 12574 37154 12626
rect 37154 12574 37156 12626
rect 37100 12572 37156 12574
rect 34076 11676 34132 11732
rect 33740 10332 33796 10388
rect 33516 8092 33572 8148
rect 34076 7810 34132 7812
rect 34076 7758 34078 7810
rect 34078 7758 34130 7810
rect 34130 7758 34132 7810
rect 34076 7756 34132 7758
rect 35196 11114 35252 11116
rect 35196 11062 35198 11114
rect 35198 11062 35250 11114
rect 35250 11062 35252 11114
rect 35196 11060 35252 11062
rect 35300 11114 35356 11116
rect 35300 11062 35302 11114
rect 35302 11062 35354 11114
rect 35354 11062 35356 11114
rect 35300 11060 35356 11062
rect 35404 11114 35460 11116
rect 35404 11062 35406 11114
rect 35406 11062 35458 11114
rect 35458 11062 35460 11114
rect 35404 11060 35460 11062
rect 34748 9602 34804 9604
rect 34748 9550 34750 9602
rect 34750 9550 34802 9602
rect 34802 9550 34804 9602
rect 34748 9548 34804 9550
rect 35196 9098 35252 9100
rect 35196 9046 35198 9098
rect 35198 9046 35250 9098
rect 35250 9046 35252 9098
rect 35196 9044 35252 9046
rect 35300 9098 35356 9100
rect 35300 9046 35302 9098
rect 35302 9046 35354 9098
rect 35354 9046 35356 9098
rect 35300 9044 35356 9046
rect 35404 9098 35460 9100
rect 35404 9046 35406 9098
rect 35406 9046 35458 9098
rect 35458 9046 35460 9098
rect 35404 9044 35460 9046
rect 36092 9602 36148 9604
rect 36092 9550 36094 9602
rect 36094 9550 36146 9602
rect 36146 9550 36148 9602
rect 36092 9548 36148 9550
rect 35644 9490 35700 9492
rect 35644 9438 35646 9490
rect 35646 9438 35698 9490
rect 35698 9438 35700 9490
rect 35644 9436 35700 9438
rect 36540 9436 36596 9492
rect 38668 20300 38724 20356
rect 40012 20300 40068 20356
rect 38332 18620 38388 18676
rect 38556 18562 38612 18564
rect 38556 18510 38558 18562
rect 38558 18510 38610 18562
rect 38610 18510 38612 18562
rect 38556 18508 38612 18510
rect 38108 18284 38164 18340
rect 39340 18674 39396 18676
rect 39340 18622 39342 18674
rect 39342 18622 39394 18674
rect 39394 18622 39396 18674
rect 39340 18620 39396 18622
rect 40236 19458 40292 19460
rect 40236 19406 40238 19458
rect 40238 19406 40290 19458
rect 40290 19406 40292 19458
rect 40236 19404 40292 19406
rect 41020 22540 41076 22596
rect 41020 21644 41076 21700
rect 40796 20300 40852 20356
rect 40908 20188 40964 20244
rect 38220 16658 38276 16660
rect 38220 16606 38222 16658
rect 38222 16606 38274 16658
rect 38274 16606 38276 16658
rect 38220 16604 38276 16606
rect 37772 16546 37828 16548
rect 37772 16494 37774 16546
rect 37774 16494 37826 16546
rect 37826 16494 37828 16546
rect 37772 16492 37828 16494
rect 37436 15762 37492 15764
rect 37436 15710 37438 15762
rect 37438 15710 37490 15762
rect 37490 15710 37492 15762
rect 37436 15708 37492 15710
rect 37324 14588 37380 14644
rect 37996 15708 38052 15764
rect 37772 14476 37828 14532
rect 37884 14924 37940 14980
rect 37324 13804 37380 13860
rect 38332 15650 38388 15652
rect 38332 15598 38334 15650
rect 38334 15598 38386 15650
rect 38386 15598 38388 15650
rect 38332 15596 38388 15598
rect 38668 14924 38724 14980
rect 38220 14754 38276 14756
rect 38220 14702 38222 14754
rect 38222 14702 38274 14754
rect 38274 14702 38276 14754
rect 38220 14700 38276 14702
rect 39676 16716 39732 16772
rect 41468 23714 41524 23716
rect 41468 23662 41470 23714
rect 41470 23662 41522 23714
rect 41522 23662 41524 23714
rect 41468 23660 41524 23662
rect 41244 22540 41300 22596
rect 41356 21868 41412 21924
rect 41468 21756 41524 21812
rect 42700 33628 42756 33684
rect 41804 32508 41860 32564
rect 41916 32844 41972 32900
rect 41692 31052 41748 31108
rect 41804 31836 41860 31892
rect 41916 30828 41972 30884
rect 41580 21644 41636 21700
rect 41468 20524 41524 20580
rect 41580 20690 41636 20692
rect 41580 20638 41582 20690
rect 41582 20638 41634 20690
rect 41634 20638 41636 20690
rect 41580 20636 41636 20638
rect 41580 20188 41636 20244
rect 41356 19794 41412 19796
rect 41356 19742 41358 19794
rect 41358 19742 41410 19794
rect 41410 19742 41412 19794
rect 41356 19740 41412 19742
rect 41244 19404 41300 19460
rect 41356 18620 41412 18676
rect 40908 18562 40964 18564
rect 40908 18510 40910 18562
rect 40910 18510 40962 18562
rect 40962 18510 40964 18562
rect 40908 18508 40964 18510
rect 40796 18396 40852 18452
rect 39452 16546 39508 16548
rect 39452 16494 39454 16546
rect 39454 16494 39506 16546
rect 39506 16494 39508 16546
rect 39452 16492 39508 16494
rect 39564 15762 39620 15764
rect 39564 15710 39566 15762
rect 39566 15710 39618 15762
rect 39618 15710 39620 15762
rect 39564 15708 39620 15710
rect 37884 12850 37940 12852
rect 37884 12798 37886 12850
rect 37886 12798 37938 12850
rect 37938 12798 37940 12850
rect 37884 12796 37940 12798
rect 38108 13580 38164 13636
rect 38556 13522 38612 13524
rect 38556 13470 38558 13522
rect 38558 13470 38610 13522
rect 38610 13470 38612 13522
rect 38556 13468 38612 13470
rect 39228 14700 39284 14756
rect 39676 14700 39732 14756
rect 39004 13468 39060 13524
rect 41244 18396 41300 18452
rect 41356 17778 41412 17780
rect 41356 17726 41358 17778
rect 41358 17726 41410 17778
rect 41410 17726 41412 17778
rect 41356 17724 41412 17726
rect 41020 15708 41076 15764
rect 41580 19292 41636 19348
rect 43148 33628 43204 33684
rect 42812 32508 42868 32564
rect 43260 31948 43316 32004
rect 42812 31890 42868 31892
rect 42812 31838 42814 31890
rect 42814 31838 42866 31890
rect 42866 31838 42868 31890
rect 42812 31836 42868 31838
rect 42140 26908 42196 26964
rect 42028 26460 42084 26516
rect 42252 25900 42308 25956
rect 42812 23826 42868 23828
rect 42812 23774 42814 23826
rect 42814 23774 42866 23826
rect 42866 23774 42868 23826
rect 42812 23772 42868 23774
rect 42140 23660 42196 23716
rect 41916 21922 41972 21924
rect 41916 21870 41918 21922
rect 41918 21870 41970 21922
rect 41970 21870 41972 21922
rect 41916 21868 41972 21870
rect 41804 21756 41860 21812
rect 42364 21810 42420 21812
rect 42364 21758 42366 21810
rect 42366 21758 42418 21810
rect 42418 21758 42420 21810
rect 42364 21756 42420 21758
rect 43484 32508 43540 32564
rect 44380 36034 44436 36036
rect 44380 35982 44382 36034
rect 44382 35982 44434 36034
rect 44434 35982 44436 36034
rect 44380 35980 44436 35982
rect 44268 34748 44324 34804
rect 43820 33794 43876 33796
rect 43820 33742 43822 33794
rect 43822 33742 43874 33794
rect 43874 33742 43876 33794
rect 43820 33740 43876 33742
rect 44156 32562 44212 32564
rect 44156 32510 44158 32562
rect 44158 32510 44210 32562
rect 44210 32510 44212 32562
rect 44156 32508 44212 32510
rect 44044 31890 44100 31892
rect 44044 31838 44046 31890
rect 44046 31838 44098 31890
rect 44098 31838 44100 31890
rect 44044 31836 44100 31838
rect 43820 31612 43876 31668
rect 43708 30716 43764 30772
rect 43484 30044 43540 30100
rect 43372 29986 43428 29988
rect 43372 29934 43374 29986
rect 43374 29934 43426 29986
rect 43426 29934 43428 29986
rect 43372 29932 43428 29934
rect 44828 37772 44884 37828
rect 45276 37826 45332 37828
rect 45276 37774 45278 37826
rect 45278 37774 45330 37826
rect 45330 37774 45332 37826
rect 45276 37772 45332 37774
rect 44940 36764 44996 36820
rect 47180 38722 47236 38724
rect 47180 38670 47182 38722
rect 47182 38670 47234 38722
rect 47234 38670 47236 38722
rect 47180 38668 47236 38670
rect 48300 38668 48356 38724
rect 47292 37938 47348 37940
rect 47292 37886 47294 37938
rect 47294 37886 47346 37938
rect 47346 37886 47348 37938
rect 47292 37884 47348 37886
rect 46172 36818 46228 36820
rect 46172 36766 46174 36818
rect 46174 36766 46226 36818
rect 46226 36766 46228 36818
rect 46172 36764 46228 36766
rect 47180 36764 47236 36820
rect 46732 36706 46788 36708
rect 46732 36654 46734 36706
rect 46734 36654 46786 36706
rect 46786 36654 46788 36706
rect 46732 36652 46788 36654
rect 44828 36034 44884 36036
rect 44828 35982 44830 36034
rect 44830 35982 44882 36034
rect 44882 35982 44884 36034
rect 44828 35980 44884 35982
rect 45052 34690 45108 34692
rect 45052 34638 45054 34690
rect 45054 34638 45106 34690
rect 45106 34638 45108 34690
rect 45052 34636 45108 34638
rect 44380 32002 44436 32004
rect 44380 31950 44382 32002
rect 44382 31950 44434 32002
rect 44434 31950 44436 32002
rect 44380 31948 44436 31950
rect 44828 33852 44884 33908
rect 44268 31724 44324 31780
rect 44044 30882 44100 30884
rect 44044 30830 44046 30882
rect 44046 30830 44098 30882
rect 44098 30830 44100 30882
rect 44044 30828 44100 30830
rect 43932 30156 43988 30212
rect 44492 29762 44548 29764
rect 44492 29710 44494 29762
rect 44494 29710 44546 29762
rect 44546 29710 44548 29762
rect 44492 29708 44548 29710
rect 45612 36034 45668 36036
rect 45612 35982 45614 36034
rect 45614 35982 45666 36034
rect 45666 35982 45668 36034
rect 45612 35980 45668 35982
rect 46732 36034 46788 36036
rect 46732 35982 46734 36034
rect 46734 35982 46786 36034
rect 46786 35982 46788 36034
rect 46732 35980 46788 35982
rect 46396 35756 46452 35812
rect 45164 33068 45220 33124
rect 45500 34748 45556 34804
rect 44940 32956 44996 33012
rect 46620 34748 46676 34804
rect 45164 32562 45220 32564
rect 45164 32510 45166 32562
rect 45166 32510 45218 32562
rect 45218 32510 45220 32562
rect 45164 32508 45220 32510
rect 45164 31724 45220 31780
rect 44940 31612 44996 31668
rect 45388 31666 45444 31668
rect 45388 31614 45390 31666
rect 45390 31614 45442 31666
rect 45442 31614 45444 31666
rect 45388 31612 45444 31614
rect 46284 33906 46340 33908
rect 46284 33854 46286 33906
rect 46286 33854 46338 33906
rect 46338 33854 46340 33906
rect 46284 33852 46340 33854
rect 46060 33010 46116 33012
rect 46060 32958 46062 33010
rect 46062 32958 46114 33010
rect 46114 32958 46116 33010
rect 46060 32956 46116 32958
rect 47068 33906 47124 33908
rect 47068 33854 47070 33906
rect 47070 33854 47122 33906
rect 47122 33854 47124 33906
rect 47068 33852 47124 33854
rect 48188 36764 48244 36820
rect 47516 34748 47572 34804
rect 47740 36706 47796 36708
rect 47740 36654 47742 36706
rect 47742 36654 47794 36706
rect 47794 36654 47796 36706
rect 47740 36652 47796 36654
rect 47740 35980 47796 36036
rect 49196 39954 49252 39956
rect 49196 39902 49198 39954
rect 49198 39902 49250 39954
rect 49250 39902 49252 39954
rect 49196 39900 49252 39902
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 49420 41580 49476 41636
rect 49756 42140 49812 42196
rect 49868 42028 49924 42084
rect 50876 41916 50932 41972
rect 50876 41746 50932 41748
rect 50876 41694 50878 41746
rect 50878 41694 50930 41746
rect 50930 41694 50932 41746
rect 50876 41692 50932 41694
rect 49868 39954 49924 39956
rect 49868 39902 49870 39954
rect 49870 39902 49922 39954
rect 49922 39902 49924 39954
rect 49868 39900 49924 39902
rect 50556 40346 50612 40348
rect 50556 40294 50558 40346
rect 50558 40294 50610 40346
rect 50610 40294 50612 40346
rect 50556 40292 50612 40294
rect 50660 40346 50716 40348
rect 50660 40294 50662 40346
rect 50662 40294 50714 40346
rect 50714 40294 50716 40346
rect 50660 40292 50716 40294
rect 50764 40346 50820 40348
rect 50764 40294 50766 40346
rect 50766 40294 50818 40346
rect 50818 40294 50820 40346
rect 50764 40292 50820 40294
rect 50540 39842 50596 39844
rect 50540 39790 50542 39842
rect 50542 39790 50594 39842
rect 50594 39790 50596 39842
rect 50540 39788 50596 39790
rect 50988 39900 51044 39956
rect 51100 41804 51156 41860
rect 51660 42642 51716 42644
rect 51660 42590 51662 42642
rect 51662 42590 51714 42642
rect 51714 42590 51716 42642
rect 51660 42588 51716 42590
rect 51660 42028 51716 42084
rect 51212 41692 51268 41748
rect 52108 42140 52164 42196
rect 48860 37714 48916 37716
rect 48860 37662 48862 37714
rect 48862 37662 48914 37714
rect 48914 37662 48916 37714
rect 48860 37660 48916 37662
rect 50540 38668 50596 38724
rect 50092 37660 50148 37716
rect 50556 38330 50612 38332
rect 50556 38278 50558 38330
rect 50558 38278 50610 38330
rect 50610 38278 50612 38330
rect 50556 38276 50612 38278
rect 50660 38330 50716 38332
rect 50660 38278 50662 38330
rect 50662 38278 50714 38330
rect 50714 38278 50716 38330
rect 50660 38276 50716 38278
rect 50764 38330 50820 38332
rect 50764 38278 50766 38330
rect 50766 38278 50818 38330
rect 50818 38278 50820 38330
rect 50764 38276 50820 38278
rect 49756 36652 49812 36708
rect 48748 35810 48804 35812
rect 48748 35758 48750 35810
rect 48750 35758 48802 35810
rect 48802 35758 48804 35810
rect 48748 35756 48804 35758
rect 49644 34802 49700 34804
rect 49644 34750 49646 34802
rect 49646 34750 49698 34802
rect 49698 34750 49700 34802
rect 49644 34748 49700 34750
rect 49308 34636 49364 34692
rect 47180 33628 47236 33684
rect 48188 33682 48244 33684
rect 48188 33630 48190 33682
rect 48190 33630 48242 33682
rect 48242 33630 48244 33682
rect 48188 33628 48244 33630
rect 49084 34412 49140 34468
rect 46396 31778 46452 31780
rect 46396 31726 46398 31778
rect 46398 31726 46450 31778
rect 46450 31726 46452 31778
rect 46396 31724 46452 31726
rect 45276 30828 45332 30884
rect 46620 30828 46676 30884
rect 47180 31890 47236 31892
rect 47180 31838 47182 31890
rect 47182 31838 47234 31890
rect 47234 31838 47236 31890
rect 47180 31836 47236 31838
rect 47516 31836 47572 31892
rect 46956 31724 47012 31780
rect 46732 31612 46788 31668
rect 45948 30770 46004 30772
rect 45948 30718 45950 30770
rect 45950 30718 46002 30770
rect 46002 30718 46004 30770
rect 45948 30716 46004 30718
rect 47964 31778 48020 31780
rect 47964 31726 47966 31778
rect 47966 31726 48018 31778
rect 48018 31726 48020 31778
rect 47964 31724 48020 31726
rect 46844 30716 46900 30772
rect 46060 30044 46116 30100
rect 45612 28700 45668 28756
rect 45164 28530 45220 28532
rect 45164 28478 45166 28530
rect 45166 28478 45218 28530
rect 45218 28478 45220 28530
rect 45164 28476 45220 28478
rect 45948 28700 46004 28756
rect 46172 29708 46228 29764
rect 46508 28924 46564 28980
rect 45276 27804 45332 27860
rect 46060 27634 46116 27636
rect 46060 27582 46062 27634
rect 46062 27582 46114 27634
rect 46114 27582 46116 27634
rect 46060 27580 46116 27582
rect 43932 26348 43988 26404
rect 43932 23884 43988 23940
rect 44828 26460 44884 26516
rect 45500 26514 45556 26516
rect 45500 26462 45502 26514
rect 45502 26462 45554 26514
rect 45554 26462 45556 26514
rect 45500 26460 45556 26462
rect 45836 26124 45892 26180
rect 45948 25564 46004 25620
rect 44828 23938 44884 23940
rect 44828 23886 44830 23938
rect 44830 23886 44882 23938
rect 44882 23886 44884 23938
rect 44828 23884 44884 23886
rect 45276 23996 45332 24052
rect 43596 23548 43652 23604
rect 45724 23826 45780 23828
rect 45724 23774 45726 23826
rect 45726 23774 45778 23826
rect 45778 23774 45780 23826
rect 45724 23772 45780 23774
rect 46172 25900 46228 25956
rect 46284 25730 46340 25732
rect 46284 25678 46286 25730
rect 46286 25678 46338 25730
rect 46338 25678 46340 25730
rect 46284 25676 46340 25678
rect 48636 32732 48692 32788
rect 48748 31500 48804 31556
rect 48748 30604 48804 30660
rect 48300 30546 48356 30548
rect 48300 30494 48302 30546
rect 48302 30494 48354 30546
rect 48354 30494 48356 30546
rect 48300 30492 48356 30494
rect 48636 30380 48692 30436
rect 48188 29650 48244 29652
rect 48188 29598 48190 29650
rect 48190 29598 48242 29650
rect 48242 29598 48244 29650
rect 48188 29596 48244 29598
rect 48188 28700 48244 28756
rect 48748 28588 48804 28644
rect 47068 28476 47124 28532
rect 47740 28476 47796 28532
rect 46620 27858 46676 27860
rect 46620 27806 46622 27858
rect 46622 27806 46674 27858
rect 46674 27806 46676 27858
rect 46620 27804 46676 27806
rect 50204 36876 50260 36932
rect 51996 42028 52052 42084
rect 51996 41580 52052 41636
rect 52780 42028 52836 42084
rect 53340 42642 53396 42644
rect 53340 42590 53342 42642
rect 53342 42590 53394 42642
rect 53394 42590 53396 42642
rect 53340 42588 53396 42590
rect 53116 41970 53172 41972
rect 53116 41918 53118 41970
rect 53118 41918 53170 41970
rect 53170 41918 53172 41970
rect 53116 41916 53172 41918
rect 53788 42140 53844 42196
rect 54348 41858 54404 41860
rect 54348 41806 54350 41858
rect 54350 41806 54402 41858
rect 54402 41806 54404 41858
rect 54348 41804 54404 41806
rect 53788 40124 53844 40180
rect 53228 39954 53284 39956
rect 53228 39902 53230 39954
rect 53230 39902 53282 39954
rect 53282 39902 53284 39954
rect 53228 39900 53284 39902
rect 51996 39788 52052 39844
rect 53004 39842 53060 39844
rect 53004 39790 53006 39842
rect 53006 39790 53058 39842
rect 53058 39790 53060 39842
rect 53004 39788 53060 39790
rect 51772 38668 51828 38724
rect 51548 37826 51604 37828
rect 51548 37774 51550 37826
rect 51550 37774 51602 37826
rect 51602 37774 51604 37826
rect 51548 37772 51604 37774
rect 51436 36988 51492 37044
rect 50316 36818 50372 36820
rect 50316 36766 50318 36818
rect 50318 36766 50370 36818
rect 50370 36766 50372 36818
rect 50316 36764 50372 36766
rect 51212 36876 51268 36932
rect 51324 36764 51380 36820
rect 50540 36706 50596 36708
rect 50540 36654 50542 36706
rect 50542 36654 50594 36706
rect 50594 36654 50596 36706
rect 50540 36652 50596 36654
rect 50876 36706 50932 36708
rect 50876 36654 50878 36706
rect 50878 36654 50930 36706
rect 50930 36654 50932 36706
rect 50876 36652 50932 36654
rect 50556 36314 50612 36316
rect 50556 36262 50558 36314
rect 50558 36262 50610 36314
rect 50610 36262 50612 36314
rect 50556 36260 50612 36262
rect 50660 36314 50716 36316
rect 50660 36262 50662 36314
rect 50662 36262 50714 36314
rect 50714 36262 50716 36314
rect 50660 36260 50716 36262
rect 50764 36314 50820 36316
rect 50764 36262 50766 36314
rect 50766 36262 50818 36314
rect 50818 36262 50820 36314
rect 50764 36260 50820 36262
rect 50092 35756 50148 35812
rect 49644 34524 49700 34580
rect 49420 33628 49476 33684
rect 49420 31836 49476 31892
rect 48972 30604 49028 30660
rect 49308 30658 49364 30660
rect 49308 30606 49310 30658
rect 49310 30606 49362 30658
rect 49362 30606 49364 30658
rect 49308 30604 49364 30606
rect 49084 28588 49140 28644
rect 47740 27634 47796 27636
rect 47740 27582 47742 27634
rect 47742 27582 47794 27634
rect 47794 27582 47796 27634
rect 47740 27580 47796 27582
rect 49084 27580 49140 27636
rect 46956 27522 47012 27524
rect 46956 27470 46958 27522
rect 46958 27470 47010 27522
rect 47010 27470 47012 27522
rect 46956 27468 47012 27470
rect 48412 27468 48468 27524
rect 46508 25564 46564 25620
rect 46732 27356 46788 27412
rect 46060 23772 46116 23828
rect 45276 23548 45332 23604
rect 49084 27356 49140 27412
rect 48412 24780 48468 24836
rect 48524 26402 48580 26404
rect 48524 26350 48526 26402
rect 48526 26350 48578 26402
rect 48578 26350 48580 26402
rect 48524 26348 48580 26350
rect 46844 23772 46900 23828
rect 44604 21698 44660 21700
rect 44604 21646 44606 21698
rect 44606 21646 44658 21698
rect 44658 21646 44660 21698
rect 44604 21644 44660 21646
rect 45052 21644 45108 21700
rect 44156 21586 44212 21588
rect 44156 21534 44158 21586
rect 44158 21534 44210 21586
rect 44210 21534 44212 21586
rect 44156 21532 44212 21534
rect 42252 20636 42308 20692
rect 41804 19740 41860 19796
rect 43484 20524 43540 20580
rect 42700 20300 42756 20356
rect 43372 20412 43428 20468
rect 42700 19404 42756 19460
rect 43596 20412 43652 20468
rect 43484 20188 43540 20244
rect 45164 21532 45220 21588
rect 45724 21644 45780 21700
rect 44156 20188 44212 20244
rect 45500 21532 45556 21588
rect 46396 20690 46452 20692
rect 46396 20638 46398 20690
rect 46398 20638 46450 20690
rect 46450 20638 46452 20690
rect 46396 20636 46452 20638
rect 45948 20578 46004 20580
rect 45948 20526 45950 20578
rect 45950 20526 46002 20578
rect 46002 20526 46004 20578
rect 45948 20524 46004 20526
rect 45724 20412 45780 20468
rect 44268 19458 44324 19460
rect 44268 19406 44270 19458
rect 44270 19406 44322 19458
rect 44322 19406 44324 19458
rect 44268 19404 44324 19406
rect 41692 15820 41748 15876
rect 41580 15708 41636 15764
rect 45612 18508 45668 18564
rect 43484 18396 43540 18452
rect 42924 17778 42980 17780
rect 42924 17726 42926 17778
rect 42926 17726 42978 17778
rect 42978 17726 42980 17778
rect 42924 17724 42980 17726
rect 42924 16828 42980 16884
rect 43932 17666 43988 17668
rect 43932 17614 43934 17666
rect 43934 17614 43986 17666
rect 43986 17614 43988 17666
rect 43932 17612 43988 17614
rect 43036 16658 43092 16660
rect 43036 16606 43038 16658
rect 43038 16606 43090 16658
rect 43090 16606 43092 16658
rect 43036 16604 43092 16606
rect 42364 15874 42420 15876
rect 42364 15822 42366 15874
rect 42366 15822 42418 15874
rect 42418 15822 42420 15874
rect 42364 15820 42420 15822
rect 41692 15372 41748 15428
rect 42364 15372 42420 15428
rect 41468 15036 41524 15092
rect 40236 14754 40292 14756
rect 40236 14702 40238 14754
rect 40238 14702 40290 14754
rect 40290 14702 40292 14754
rect 40236 14700 40292 14702
rect 41356 13858 41412 13860
rect 41356 13806 41358 13858
rect 41358 13806 41410 13858
rect 41410 13806 41412 13858
rect 41356 13804 41412 13806
rect 40348 13692 40404 13748
rect 39900 13468 39956 13524
rect 38108 12796 38164 12852
rect 37324 12572 37380 12628
rect 38668 12572 38724 12628
rect 39004 12626 39060 12628
rect 39004 12574 39006 12626
rect 39006 12574 39058 12626
rect 39058 12574 39060 12626
rect 39004 12572 39060 12574
rect 39340 12626 39396 12628
rect 39340 12574 39342 12626
rect 39342 12574 39394 12626
rect 39394 12574 39396 12626
rect 39340 12572 39396 12574
rect 39676 12796 39732 12852
rect 40012 12572 40068 12628
rect 37212 9324 37268 9380
rect 37324 10556 37380 10612
rect 38332 10610 38388 10612
rect 38332 10558 38334 10610
rect 38334 10558 38386 10610
rect 38386 10558 38388 10610
rect 38332 10556 38388 10558
rect 37324 9548 37380 9604
rect 35644 8652 35700 8708
rect 36204 8706 36260 8708
rect 36204 8654 36206 8706
rect 36206 8654 36258 8706
rect 36258 8654 36260 8706
rect 36204 8652 36260 8654
rect 39228 10556 39284 10612
rect 39676 10610 39732 10612
rect 39676 10558 39678 10610
rect 39678 10558 39730 10610
rect 39730 10558 39732 10610
rect 39676 10556 39732 10558
rect 39452 10444 39508 10500
rect 37660 9436 37716 9492
rect 35308 8092 35364 8148
rect 36652 8092 36708 8148
rect 37660 8316 37716 8372
rect 38780 8428 38836 8484
rect 41020 13746 41076 13748
rect 41020 13694 41022 13746
rect 41022 13694 41074 13746
rect 41074 13694 41076 13746
rect 41020 13692 41076 13694
rect 42700 15036 42756 15092
rect 42364 13804 42420 13860
rect 42140 12460 42196 12516
rect 40012 8652 40068 8708
rect 40348 10556 40404 10612
rect 40124 10444 40180 10500
rect 40236 9602 40292 9604
rect 40236 9550 40238 9602
rect 40238 9550 40290 9602
rect 40290 9550 40292 9602
rect 40236 9548 40292 9550
rect 40908 9602 40964 9604
rect 40908 9550 40910 9602
rect 40910 9550 40962 9602
rect 40962 9550 40964 9602
rect 40908 9548 40964 9550
rect 41244 9324 41300 9380
rect 40460 8652 40516 8708
rect 40236 8428 40292 8484
rect 40124 8316 40180 8372
rect 41020 8540 41076 8596
rect 38780 8092 38836 8148
rect 41916 9826 41972 9828
rect 41916 9774 41918 9826
rect 41918 9774 41970 9826
rect 41970 9774 41972 9826
rect 41916 9772 41972 9774
rect 45724 18450 45780 18452
rect 45724 18398 45726 18450
rect 45726 18398 45778 18450
rect 45778 18398 45780 18450
rect 45724 18396 45780 18398
rect 45276 17612 45332 17668
rect 45948 17666 46004 17668
rect 45948 17614 45950 17666
rect 45950 17614 46002 17666
rect 46002 17614 46004 17666
rect 45948 17612 46004 17614
rect 43932 16492 43988 16548
rect 44716 16380 44772 16436
rect 44828 16716 44884 16772
rect 46284 18396 46340 18452
rect 46396 20188 46452 20244
rect 46732 20076 46788 20132
rect 43484 15762 43540 15764
rect 43484 15710 43486 15762
rect 43486 15710 43538 15762
rect 43538 15710 43540 15762
rect 43484 15708 43540 15710
rect 44940 15708 44996 15764
rect 43260 12796 43316 12852
rect 43820 14754 43876 14756
rect 43820 14702 43822 14754
rect 43822 14702 43874 14754
rect 43874 14702 43876 14754
rect 43820 14700 43876 14702
rect 43484 14476 43540 14532
rect 42924 12514 42980 12516
rect 42924 12462 42926 12514
rect 42926 12462 42978 12514
rect 42978 12462 42980 12514
rect 42924 12460 42980 12462
rect 46060 16434 46116 16436
rect 46060 16382 46062 16434
rect 46062 16382 46114 16434
rect 46114 16382 46116 16434
rect 46060 16380 46116 16382
rect 46956 19740 47012 19796
rect 46620 17836 46676 17892
rect 46732 18396 46788 18452
rect 47068 18562 47124 18564
rect 47068 18510 47070 18562
rect 47070 18510 47122 18562
rect 47122 18510 47124 18562
rect 47068 18508 47124 18510
rect 47740 23996 47796 24052
rect 47516 23938 47572 23940
rect 47516 23886 47518 23938
rect 47518 23886 47570 23938
rect 47570 23886 47572 23938
rect 47516 23884 47572 23886
rect 48188 24332 48244 24388
rect 49308 29596 49364 29652
rect 50876 34636 50932 34692
rect 53564 39788 53620 39844
rect 54012 39842 54068 39844
rect 54012 39790 54014 39842
rect 54014 39790 54066 39842
rect 54066 39790 54068 39842
rect 54012 39788 54068 39790
rect 54572 39954 54628 39956
rect 54572 39902 54574 39954
rect 54574 39902 54626 39954
rect 54626 39902 54628 39954
rect 54572 39900 54628 39902
rect 54684 40348 54740 40404
rect 54348 39676 54404 39732
rect 55580 40348 55636 40404
rect 55356 39842 55412 39844
rect 55356 39790 55358 39842
rect 55358 39790 55410 39842
rect 55410 39790 55412 39842
rect 55356 39788 55412 39790
rect 53676 38780 53732 38836
rect 53676 37436 53732 37492
rect 51996 36764 52052 36820
rect 51660 36428 51716 36484
rect 51884 36540 51940 36596
rect 51100 34748 51156 34804
rect 50764 34578 50820 34580
rect 50764 34526 50766 34578
rect 50766 34526 50818 34578
rect 50818 34526 50820 34578
rect 50764 34524 50820 34526
rect 50876 34466 50932 34468
rect 50876 34414 50878 34466
rect 50878 34414 50930 34466
rect 50930 34414 50932 34466
rect 50876 34412 50932 34414
rect 50556 34298 50612 34300
rect 50556 34246 50558 34298
rect 50558 34246 50610 34298
rect 50610 34246 50612 34298
rect 50556 34244 50612 34246
rect 50660 34298 50716 34300
rect 50660 34246 50662 34298
rect 50662 34246 50714 34298
rect 50714 34246 50716 34298
rect 50660 34244 50716 34246
rect 50764 34298 50820 34300
rect 50764 34246 50766 34298
rect 50766 34246 50818 34298
rect 50818 34246 50820 34298
rect 50764 34244 50820 34246
rect 50316 33516 50372 33572
rect 51548 34860 51604 34916
rect 51324 34690 51380 34692
rect 51324 34638 51326 34690
rect 51326 34638 51378 34690
rect 51378 34638 51380 34690
rect 51324 34636 51380 34638
rect 54348 37490 54404 37492
rect 54348 37438 54350 37490
rect 54350 37438 54402 37490
rect 54402 37438 54404 37490
rect 54348 37436 54404 37438
rect 53788 36988 53844 37044
rect 53452 36428 53508 36484
rect 52332 36034 52388 36036
rect 52332 35982 52334 36034
rect 52334 35982 52386 36034
rect 52386 35982 52388 36034
rect 52332 35980 52388 35982
rect 52780 35980 52836 36036
rect 56140 39788 56196 39844
rect 56476 39676 56532 39732
rect 57148 39730 57204 39732
rect 57148 39678 57150 39730
rect 57150 39678 57202 39730
rect 57202 39678 57204 39730
rect 57148 39676 57204 39678
rect 56700 38556 56756 38612
rect 57036 38610 57092 38612
rect 57036 38558 57038 38610
rect 57038 38558 57090 38610
rect 57090 38558 57092 38610
rect 57036 38556 57092 38558
rect 55356 36988 55412 37044
rect 54460 36876 54516 36932
rect 55132 36706 55188 36708
rect 55132 36654 55134 36706
rect 55134 36654 55186 36706
rect 55186 36654 55188 36706
rect 55132 36652 55188 36654
rect 55356 36652 55412 36708
rect 55580 37714 55636 37716
rect 55580 37662 55582 37714
rect 55582 37662 55634 37714
rect 55634 37662 55636 37714
rect 55580 37660 55636 37662
rect 54012 36594 54068 36596
rect 54012 36542 54014 36594
rect 54014 36542 54066 36594
rect 54066 36542 54068 36594
rect 54012 36540 54068 36542
rect 55244 36428 55300 36484
rect 53676 35810 53732 35812
rect 53676 35758 53678 35810
rect 53678 35758 53730 35810
rect 53730 35758 53732 35810
rect 53676 35756 53732 35758
rect 53452 35308 53508 35364
rect 53004 34802 53060 34804
rect 53004 34750 53006 34802
rect 53006 34750 53058 34802
rect 53058 34750 53060 34802
rect 53004 34748 53060 34750
rect 53452 34802 53508 34804
rect 53452 34750 53454 34802
rect 53454 34750 53506 34802
rect 53506 34750 53508 34802
rect 53452 34748 53508 34750
rect 53228 34636 53284 34692
rect 50556 32282 50612 32284
rect 50556 32230 50558 32282
rect 50558 32230 50610 32282
rect 50610 32230 50612 32282
rect 50556 32228 50612 32230
rect 50660 32282 50716 32284
rect 50660 32230 50662 32282
rect 50662 32230 50714 32282
rect 50714 32230 50716 32282
rect 50660 32228 50716 32230
rect 50764 32282 50820 32284
rect 50764 32230 50766 32282
rect 50766 32230 50818 32282
rect 50818 32230 50820 32282
rect 50764 32228 50820 32230
rect 50204 31836 50260 31892
rect 50204 31666 50260 31668
rect 50204 31614 50206 31666
rect 50206 31614 50258 31666
rect 50258 31614 50260 31666
rect 50204 31612 50260 31614
rect 49532 31500 49588 31556
rect 50316 30716 50372 30772
rect 49980 30546 50036 30548
rect 49980 30494 49982 30546
rect 49982 30494 50034 30546
rect 50034 30494 50036 30546
rect 49980 30492 50036 30494
rect 49644 29874 49700 29876
rect 49644 29822 49646 29874
rect 49646 29822 49698 29874
rect 49698 29822 49700 29874
rect 49644 29820 49700 29822
rect 49868 29708 49924 29764
rect 49756 28812 49812 28868
rect 50316 28700 50372 28756
rect 50556 30266 50612 30268
rect 50556 30214 50558 30266
rect 50558 30214 50610 30266
rect 50610 30214 50612 30266
rect 50556 30212 50612 30214
rect 50660 30266 50716 30268
rect 50660 30214 50662 30266
rect 50662 30214 50714 30266
rect 50714 30214 50716 30266
rect 50660 30212 50716 30214
rect 50764 30266 50820 30268
rect 50764 30214 50766 30266
rect 50766 30214 50818 30266
rect 50818 30214 50820 30266
rect 50764 30212 50820 30214
rect 50988 30268 51044 30324
rect 50876 29820 50932 29876
rect 52108 31836 52164 31892
rect 52444 31724 52500 31780
rect 51548 31500 51604 31556
rect 51660 31612 51716 31668
rect 51324 30380 51380 30436
rect 54236 35980 54292 36036
rect 54572 35810 54628 35812
rect 54572 35758 54574 35810
rect 54574 35758 54626 35810
rect 54626 35758 54628 35810
rect 54572 35756 54628 35758
rect 57036 37660 57092 37716
rect 57596 37714 57652 37716
rect 57596 37662 57598 37714
rect 57598 37662 57650 37714
rect 57650 37662 57652 37714
rect 57596 37660 57652 37662
rect 56700 36652 56756 36708
rect 55580 35756 55636 35812
rect 55020 35420 55076 35476
rect 54348 33964 54404 34020
rect 55580 35474 55636 35476
rect 55580 35422 55582 35474
rect 55582 35422 55634 35474
rect 55634 35422 55636 35474
rect 55580 35420 55636 35422
rect 56588 36594 56644 36596
rect 56588 36542 56590 36594
rect 56590 36542 56642 36594
rect 56642 36542 56644 36594
rect 56588 36540 56644 36542
rect 57148 36988 57204 37044
rect 57484 36988 57540 37044
rect 56924 35756 56980 35812
rect 55916 35308 55972 35364
rect 55804 34018 55860 34020
rect 55804 33966 55806 34018
rect 55806 33966 55858 34018
rect 55858 33966 55860 34018
rect 55804 33964 55860 33966
rect 55580 33740 55636 33796
rect 53676 32732 53732 32788
rect 53900 33516 53956 33572
rect 55692 33628 55748 33684
rect 55132 32732 55188 32788
rect 52780 31612 52836 31668
rect 53676 31836 53732 31892
rect 53452 31778 53508 31780
rect 53452 31726 53454 31778
rect 53454 31726 53506 31778
rect 53506 31726 53508 31778
rect 53452 31724 53508 31726
rect 53340 31500 53396 31556
rect 52556 30434 52612 30436
rect 52556 30382 52558 30434
rect 52558 30382 52610 30434
rect 52610 30382 52612 30434
rect 52556 30380 52612 30382
rect 52444 30268 52500 30324
rect 53564 30658 53620 30660
rect 53564 30606 53566 30658
rect 53566 30606 53618 30658
rect 53618 30606 53620 30658
rect 53564 30604 53620 30606
rect 54236 30658 54292 30660
rect 54236 30606 54238 30658
rect 54238 30606 54290 30658
rect 54290 30606 54292 30658
rect 54236 30604 54292 30606
rect 53004 30268 53060 30324
rect 54236 30268 54292 30324
rect 52780 29874 52836 29876
rect 52780 29822 52782 29874
rect 52782 29822 52834 29874
rect 52834 29822 52836 29874
rect 52780 29820 52836 29822
rect 50540 28700 50596 28756
rect 50988 28588 51044 28644
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 49308 26514 49364 26516
rect 49308 26462 49310 26514
rect 49310 26462 49362 26514
rect 49362 26462 49364 26514
rect 49308 26460 49364 26462
rect 49308 25954 49364 25956
rect 49308 25902 49310 25954
rect 49310 25902 49362 25954
rect 49362 25902 49364 25954
rect 49308 25900 49364 25902
rect 48748 23996 48804 24052
rect 48636 23884 48692 23940
rect 50428 26908 50484 26964
rect 50204 26460 50260 26516
rect 49644 24332 49700 24388
rect 51324 27916 51380 27972
rect 53452 29762 53508 29764
rect 53452 29710 53454 29762
rect 53454 29710 53506 29762
rect 53506 29710 53508 29762
rect 53452 29708 53508 29710
rect 52780 28812 52836 28868
rect 54012 28866 54068 28868
rect 54012 28814 54014 28866
rect 54014 28814 54066 28866
rect 54066 28814 54068 28866
rect 54012 28812 54068 28814
rect 52780 28642 52836 28644
rect 52780 28590 52782 28642
rect 52782 28590 52834 28642
rect 52834 28590 52836 28642
rect 52780 28588 52836 28590
rect 51324 27468 51380 27524
rect 50540 26460 50596 26516
rect 49980 24050 50036 24052
rect 49980 23998 49982 24050
rect 49982 23998 50034 24050
rect 50034 23998 50036 24050
rect 49980 23996 50036 23998
rect 49532 23884 49588 23940
rect 48972 23772 49028 23828
rect 49644 23548 49700 23604
rect 50556 26234 50612 26236
rect 50556 26182 50558 26234
rect 50558 26182 50610 26234
rect 50610 26182 50612 26234
rect 50556 26180 50612 26182
rect 50660 26234 50716 26236
rect 50660 26182 50662 26234
rect 50662 26182 50714 26234
rect 50714 26182 50716 26234
rect 50660 26180 50716 26182
rect 50764 26234 50820 26236
rect 50764 26182 50766 26234
rect 50766 26182 50818 26234
rect 50818 26182 50820 26234
rect 50764 26180 50820 26182
rect 51100 26460 51156 26516
rect 51436 26684 51492 26740
rect 51996 27692 52052 27748
rect 50764 25900 50820 25956
rect 50876 25676 50932 25732
rect 50556 24218 50612 24220
rect 50556 24166 50558 24218
rect 50558 24166 50610 24218
rect 50610 24166 50612 24218
rect 50556 24164 50612 24166
rect 50660 24218 50716 24220
rect 50660 24166 50662 24218
rect 50662 24166 50714 24218
rect 50714 24166 50716 24218
rect 50660 24164 50716 24166
rect 50764 24218 50820 24220
rect 50764 24166 50766 24218
rect 50766 24166 50818 24218
rect 50818 24166 50820 24218
rect 50764 24164 50820 24166
rect 50204 23660 50260 23716
rect 48524 21644 48580 21700
rect 47628 20578 47684 20580
rect 47628 20526 47630 20578
rect 47630 20526 47682 20578
rect 47682 20526 47684 20578
rect 47628 20524 47684 20526
rect 47516 20188 47572 20244
rect 47628 19740 47684 19796
rect 48076 20690 48132 20692
rect 48076 20638 48078 20690
rect 48078 20638 48130 20690
rect 48130 20638 48132 20690
rect 48076 20636 48132 20638
rect 47740 20412 47796 20468
rect 48636 20300 48692 20356
rect 49084 21756 49140 21812
rect 48860 21698 48916 21700
rect 48860 21646 48862 21698
rect 48862 21646 48914 21698
rect 48914 21646 48916 21698
rect 48860 21644 48916 21646
rect 50428 23602 50484 23604
rect 50428 23550 50430 23602
rect 50430 23550 50482 23602
rect 50482 23550 50484 23602
rect 50428 23548 50484 23550
rect 49756 21420 49812 21476
rect 49532 20412 49588 20468
rect 47404 17948 47460 18004
rect 47740 18508 47796 18564
rect 47180 17612 47236 17668
rect 49084 18732 49140 18788
rect 48860 18674 48916 18676
rect 48860 18622 48862 18674
rect 48862 18622 48914 18674
rect 48914 18622 48916 18674
rect 48860 18620 48916 18622
rect 47964 18562 48020 18564
rect 47964 18510 47966 18562
rect 47966 18510 48018 18562
rect 48018 18510 48020 18562
rect 47964 18508 48020 18510
rect 48188 17890 48244 17892
rect 48188 17838 48190 17890
rect 48190 17838 48242 17890
rect 48242 17838 48244 17890
rect 48188 17836 48244 17838
rect 47516 16604 47572 16660
rect 47740 16716 47796 16772
rect 47180 15820 47236 15876
rect 47068 15650 47124 15652
rect 47068 15598 47070 15650
rect 47070 15598 47122 15650
rect 47122 15598 47124 15650
rect 47068 15596 47124 15598
rect 45836 14754 45892 14756
rect 45836 14702 45838 14754
rect 45838 14702 45890 14754
rect 45890 14702 45892 14754
rect 45836 14700 45892 14702
rect 45388 14642 45444 14644
rect 45388 14590 45390 14642
rect 45390 14590 45442 14642
rect 45442 14590 45444 14642
rect 45388 14588 45444 14590
rect 44940 14530 44996 14532
rect 44940 14478 44942 14530
rect 44942 14478 44994 14530
rect 44994 14478 44996 14530
rect 44940 14476 44996 14478
rect 46396 14476 46452 14532
rect 44268 14418 44324 14420
rect 44268 14366 44270 14418
rect 44270 14366 44322 14418
rect 44322 14366 44324 14418
rect 44268 14364 44324 14366
rect 45612 14364 45668 14420
rect 46732 14418 46788 14420
rect 46732 14366 46734 14418
rect 46734 14366 46786 14418
rect 46786 14366 46788 14418
rect 46732 14364 46788 14366
rect 43820 12796 43876 12852
rect 46284 12796 46340 12852
rect 43484 12460 43540 12516
rect 44492 12572 44548 12628
rect 43596 10444 43652 10500
rect 44044 11730 44100 11732
rect 44044 11678 44046 11730
rect 44046 11678 44098 11730
rect 44098 11678 44100 11730
rect 44044 11676 44100 11678
rect 44940 12514 44996 12516
rect 44940 12462 44942 12514
rect 44942 12462 44994 12514
rect 44994 12462 44996 12514
rect 44940 12460 44996 12462
rect 49756 19628 49812 19684
rect 49868 20636 49924 20692
rect 49420 18562 49476 18564
rect 49420 18510 49422 18562
rect 49422 18510 49474 18562
rect 49474 18510 49476 18562
rect 49420 18508 49476 18510
rect 49532 17836 49588 17892
rect 49980 19682 50036 19684
rect 49980 19630 49982 19682
rect 49982 19630 50034 19682
rect 50034 19630 50036 19682
rect 49980 19628 50036 19630
rect 50988 24780 51044 24836
rect 51212 24444 51268 24500
rect 51324 23772 51380 23828
rect 51100 23548 51156 23604
rect 50556 22202 50612 22204
rect 50556 22150 50558 22202
rect 50558 22150 50610 22202
rect 50610 22150 50612 22202
rect 50556 22148 50612 22150
rect 50660 22202 50716 22204
rect 50660 22150 50662 22202
rect 50662 22150 50714 22202
rect 50714 22150 50716 22202
rect 50660 22148 50716 22150
rect 50764 22202 50820 22204
rect 50764 22150 50766 22202
rect 50766 22150 50818 22202
rect 50818 22150 50820 22202
rect 50764 22148 50820 22150
rect 50876 21756 50932 21812
rect 50988 21698 51044 21700
rect 50988 21646 50990 21698
rect 50990 21646 51042 21698
rect 51042 21646 51044 21698
rect 50988 21644 51044 21646
rect 50540 20690 50596 20692
rect 50540 20638 50542 20690
rect 50542 20638 50594 20690
rect 50594 20638 50596 20690
rect 50540 20636 50596 20638
rect 50204 20300 50260 20356
rect 50556 20186 50612 20188
rect 50556 20134 50558 20186
rect 50558 20134 50610 20186
rect 50610 20134 50612 20186
rect 50556 20132 50612 20134
rect 50660 20186 50716 20188
rect 50660 20134 50662 20186
rect 50662 20134 50714 20186
rect 50714 20134 50716 20186
rect 50660 20132 50716 20134
rect 50764 20186 50820 20188
rect 50764 20134 50766 20186
rect 50766 20134 50818 20186
rect 50818 20134 50820 20186
rect 50764 20132 50820 20134
rect 50988 20412 51044 20468
rect 50876 19628 50932 19684
rect 49980 18844 50036 18900
rect 50092 18674 50148 18676
rect 50092 18622 50094 18674
rect 50094 18622 50146 18674
rect 50146 18622 50148 18674
rect 50092 18620 50148 18622
rect 50876 18732 50932 18788
rect 50556 18170 50612 18172
rect 50556 18118 50558 18170
rect 50558 18118 50610 18170
rect 50610 18118 50612 18170
rect 50556 18116 50612 18118
rect 50660 18170 50716 18172
rect 50660 18118 50662 18170
rect 50662 18118 50714 18170
rect 50714 18118 50716 18170
rect 50660 18116 50716 18118
rect 50764 18170 50820 18172
rect 50764 18118 50766 18170
rect 50766 18118 50818 18170
rect 50818 18118 50820 18170
rect 50764 18116 50820 18118
rect 50540 17948 50596 18004
rect 51212 23660 51268 23716
rect 51436 23436 51492 23492
rect 51548 24780 51604 24836
rect 52444 27580 52500 27636
rect 53116 27970 53172 27972
rect 53116 27918 53118 27970
rect 53118 27918 53170 27970
rect 53170 27918 53172 27970
rect 53116 27916 53172 27918
rect 52780 27746 52836 27748
rect 52780 27694 52782 27746
rect 52782 27694 52834 27746
rect 52834 27694 52836 27746
rect 52780 27692 52836 27694
rect 53116 27580 53172 27636
rect 52668 26796 52724 26852
rect 52780 26514 52836 26516
rect 52780 26462 52782 26514
rect 52782 26462 52834 26514
rect 52834 26462 52836 26514
rect 52780 26460 52836 26462
rect 51660 23772 51716 23828
rect 53564 26908 53620 26964
rect 53788 26908 53844 26964
rect 53564 26738 53620 26740
rect 53564 26686 53566 26738
rect 53566 26686 53618 26738
rect 53618 26686 53620 26738
rect 53564 26684 53620 26686
rect 53676 26460 53732 26516
rect 55020 32674 55076 32676
rect 55020 32622 55022 32674
rect 55022 32622 55074 32674
rect 55074 32622 55076 32674
rect 55020 32620 55076 32622
rect 55020 31836 55076 31892
rect 54684 30658 54740 30660
rect 54684 30606 54686 30658
rect 54686 30606 54738 30658
rect 54738 30606 54740 30658
rect 54684 30604 54740 30606
rect 57932 36706 57988 36708
rect 57932 36654 57934 36706
rect 57934 36654 57986 36706
rect 57986 36654 57988 36706
rect 57932 36652 57988 36654
rect 56700 33794 56756 33796
rect 56700 33742 56702 33794
rect 56702 33742 56754 33794
rect 56754 33742 56756 33794
rect 56700 33740 56756 33742
rect 56364 32898 56420 32900
rect 56364 32846 56366 32898
rect 56366 32846 56418 32898
rect 56418 32846 56420 32898
rect 56364 32844 56420 32846
rect 56924 32844 56980 32900
rect 57148 33852 57204 33908
rect 56252 32562 56308 32564
rect 56252 32510 56254 32562
rect 56254 32510 56306 32562
rect 56306 32510 56308 32562
rect 56252 32508 56308 32510
rect 55580 31948 55636 32004
rect 56028 31836 56084 31892
rect 54348 29820 54404 29876
rect 54796 28812 54852 28868
rect 54012 26684 54068 26740
rect 55132 28588 55188 28644
rect 56812 32674 56868 32676
rect 56812 32622 56814 32674
rect 56814 32622 56866 32674
rect 56866 32622 56868 32674
rect 56812 32620 56868 32622
rect 57708 33906 57764 33908
rect 57708 33854 57710 33906
rect 57710 33854 57762 33906
rect 57762 33854 57764 33906
rect 57708 33852 57764 33854
rect 57372 33682 57428 33684
rect 57372 33630 57374 33682
rect 57374 33630 57426 33682
rect 57426 33630 57428 33682
rect 57372 33628 57428 33630
rect 57708 32898 57764 32900
rect 57708 32846 57710 32898
rect 57710 32846 57762 32898
rect 57762 32846 57764 32898
rect 57708 32844 57764 32846
rect 56924 31836 56980 31892
rect 57036 31948 57092 32004
rect 56700 31666 56756 31668
rect 56700 31614 56702 31666
rect 56702 31614 56754 31666
rect 56754 31614 56756 31666
rect 56700 31612 56756 31614
rect 56700 30268 56756 30324
rect 55804 28476 55860 28532
rect 56924 28476 56980 28532
rect 57148 31666 57204 31668
rect 57148 31614 57150 31666
rect 57150 31614 57202 31666
rect 57202 31614 57204 31666
rect 57148 31612 57204 31614
rect 54908 27858 54964 27860
rect 54908 27806 54910 27858
rect 54910 27806 54962 27858
rect 54962 27806 54964 27858
rect 54908 27804 54964 27806
rect 55692 27746 55748 27748
rect 55692 27694 55694 27746
rect 55694 27694 55746 27746
rect 55746 27694 55748 27746
rect 55692 27692 55748 27694
rect 56588 27746 56644 27748
rect 56588 27694 56590 27746
rect 56590 27694 56642 27746
rect 56642 27694 56644 27746
rect 56588 27692 56644 27694
rect 54012 25842 54068 25844
rect 54012 25790 54014 25842
rect 54014 25790 54066 25842
rect 54066 25790 54068 25842
rect 54012 25788 54068 25790
rect 54460 25900 54516 25956
rect 55804 26738 55860 26740
rect 55804 26686 55806 26738
rect 55806 26686 55858 26738
rect 55858 26686 55860 26738
rect 55804 26684 55860 26686
rect 54572 25788 54628 25844
rect 51660 23436 51716 23492
rect 52668 23772 52724 23828
rect 51324 21308 51380 21364
rect 52780 23660 52836 23716
rect 54124 24498 54180 24500
rect 54124 24446 54126 24498
rect 54126 24446 54178 24498
rect 54178 24446 54180 24498
rect 54124 24444 54180 24446
rect 55356 25954 55412 25956
rect 55356 25902 55358 25954
rect 55358 25902 55410 25954
rect 55410 25902 55412 25954
rect 55356 25900 55412 25902
rect 55580 25618 55636 25620
rect 55580 25566 55582 25618
rect 55582 25566 55634 25618
rect 55634 25566 55636 25618
rect 55580 25564 55636 25566
rect 56028 25618 56084 25620
rect 56028 25566 56030 25618
rect 56030 25566 56082 25618
rect 56082 25566 56084 25618
rect 56028 25564 56084 25566
rect 56924 27858 56980 27860
rect 56924 27806 56926 27858
rect 56926 27806 56978 27858
rect 56978 27806 56980 27858
rect 56924 27804 56980 27806
rect 58156 27746 58212 27748
rect 58156 27694 58158 27746
rect 58158 27694 58210 27746
rect 58210 27694 58212 27746
rect 58156 27692 58212 27694
rect 57260 26908 57316 26964
rect 56700 25618 56756 25620
rect 56700 25566 56702 25618
rect 56702 25566 56754 25618
rect 56754 25566 56756 25618
rect 56700 25564 56756 25566
rect 55356 24556 55412 24612
rect 56812 24610 56868 24612
rect 56812 24558 56814 24610
rect 56814 24558 56866 24610
rect 56866 24558 56868 24610
rect 56812 24556 56868 24558
rect 54684 23772 54740 23828
rect 54460 23548 54516 23604
rect 55132 23548 55188 23604
rect 53452 22540 53508 22596
rect 51884 22428 51940 22484
rect 51772 21644 51828 21700
rect 53228 21756 53284 21812
rect 52892 21308 52948 21364
rect 52220 20636 52276 20692
rect 53116 20636 53172 20692
rect 51548 19682 51604 19684
rect 51548 19630 51550 19682
rect 51550 19630 51602 19682
rect 51602 19630 51604 19682
rect 51548 19628 51604 19630
rect 52556 18844 52612 18900
rect 53340 20412 53396 20468
rect 54348 22594 54404 22596
rect 54348 22542 54350 22594
rect 54350 22542 54402 22594
rect 54402 22542 54404 22594
rect 54348 22540 54404 22542
rect 54684 22482 54740 22484
rect 54684 22430 54686 22482
rect 54686 22430 54738 22482
rect 54738 22430 54740 22482
rect 54684 22428 54740 22430
rect 56476 22482 56532 22484
rect 56476 22430 56478 22482
rect 56478 22430 56530 22482
rect 56530 22430 56532 22482
rect 56476 22428 56532 22430
rect 57148 22482 57204 22484
rect 57148 22430 57150 22482
rect 57150 22430 57202 22482
rect 57202 22430 57204 22482
rect 57148 22428 57204 22430
rect 54908 21868 54964 21924
rect 54124 21698 54180 21700
rect 54124 21646 54126 21698
rect 54126 21646 54178 21698
rect 54178 21646 54180 21698
rect 54124 21644 54180 21646
rect 54124 20748 54180 20804
rect 54908 20802 54964 20804
rect 54908 20750 54910 20802
rect 54910 20750 54962 20802
rect 54962 20750 54964 20802
rect 54908 20748 54964 20750
rect 55244 21810 55300 21812
rect 55244 21758 55246 21810
rect 55246 21758 55298 21810
rect 55298 21758 55300 21810
rect 55244 21756 55300 21758
rect 56700 21810 56756 21812
rect 56700 21758 56702 21810
rect 56702 21758 56754 21810
rect 56754 21758 56756 21810
rect 56700 21756 56756 21758
rect 53788 20690 53844 20692
rect 53788 20638 53790 20690
rect 53790 20638 53842 20690
rect 53842 20638 53844 20690
rect 53788 20636 53844 20638
rect 53228 19628 53284 19684
rect 56028 21420 56084 21476
rect 57036 21532 57092 21588
rect 56252 20802 56308 20804
rect 56252 20750 56254 20802
rect 56254 20750 56306 20802
rect 56306 20750 56308 20802
rect 56252 20748 56308 20750
rect 57708 21756 57764 21812
rect 57148 21420 57204 21476
rect 57036 20748 57092 20804
rect 55804 20690 55860 20692
rect 55804 20638 55806 20690
rect 55806 20638 55858 20690
rect 55858 20638 55860 20690
rect 55804 20636 55860 20638
rect 47964 15650 48020 15652
rect 47964 15598 47966 15650
rect 47966 15598 48018 15650
rect 48018 15598 48020 15650
rect 47964 15596 48020 15598
rect 49308 16716 49364 16772
rect 48972 16658 49028 16660
rect 48972 16606 48974 16658
rect 48974 16606 49026 16658
rect 49026 16606 49028 16658
rect 48972 16604 49028 16606
rect 49756 16716 49812 16772
rect 49756 15650 49812 15652
rect 49756 15598 49758 15650
rect 49758 15598 49810 15650
rect 49810 15598 49812 15650
rect 49756 15596 49812 15598
rect 47180 14476 47236 14532
rect 50316 16604 50372 16660
rect 50204 16268 50260 16324
rect 50764 16268 50820 16324
rect 50876 16604 50932 16660
rect 50556 16154 50612 16156
rect 50556 16102 50558 16154
rect 50558 16102 50610 16154
rect 50610 16102 50612 16154
rect 50556 16100 50612 16102
rect 50660 16154 50716 16156
rect 50660 16102 50662 16154
rect 50662 16102 50714 16154
rect 50714 16102 50716 16154
rect 50660 16100 50716 16102
rect 50764 16154 50820 16156
rect 50764 16102 50766 16154
rect 50766 16102 50818 16154
rect 50818 16102 50820 16154
rect 50764 16100 50820 16102
rect 49980 15148 50036 15204
rect 48860 14364 48916 14420
rect 47740 12850 47796 12852
rect 47740 12798 47742 12850
rect 47742 12798 47794 12850
rect 47794 12798 47796 12850
rect 47740 12796 47796 12798
rect 50540 15260 50596 15316
rect 50764 15148 50820 15204
rect 51660 16380 51716 16436
rect 51772 16268 51828 16324
rect 51212 15874 51268 15876
rect 51212 15822 51214 15874
rect 51214 15822 51266 15874
rect 51266 15822 51268 15874
rect 51212 15820 51268 15822
rect 52556 16658 52612 16660
rect 52556 16606 52558 16658
rect 52558 16606 52610 16658
rect 52610 16606 52612 16658
rect 52556 16604 52612 16606
rect 52556 16434 52612 16436
rect 52556 16382 52558 16434
rect 52558 16382 52610 16434
rect 52610 16382 52612 16434
rect 52556 16380 52612 16382
rect 52892 15820 52948 15876
rect 53228 16380 53284 16436
rect 51772 15708 51828 15764
rect 52780 15708 52836 15764
rect 50988 15596 51044 15652
rect 50988 14754 51044 14756
rect 50988 14702 50990 14754
rect 50990 14702 51042 14754
rect 51042 14702 51044 14754
rect 50988 14700 51044 14702
rect 51660 15260 51716 15316
rect 52108 14754 52164 14756
rect 52108 14702 52110 14754
rect 52110 14702 52162 14754
rect 52162 14702 52164 14754
rect 52108 14700 52164 14702
rect 50092 14418 50148 14420
rect 50092 14366 50094 14418
rect 50094 14366 50146 14418
rect 50146 14366 50148 14418
rect 50092 14364 50148 14366
rect 52556 14588 52612 14644
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 51212 13858 51268 13860
rect 51212 13806 51214 13858
rect 51214 13806 51266 13858
rect 51266 13806 51268 13858
rect 51212 13804 51268 13806
rect 54908 16434 54964 16436
rect 54908 16382 54910 16434
rect 54910 16382 54962 16434
rect 54962 16382 54964 16434
rect 54908 16380 54964 16382
rect 54572 15708 54628 15764
rect 54236 15650 54292 15652
rect 54236 15598 54238 15650
rect 54238 15598 54290 15650
rect 54290 15598 54292 15650
rect 54236 15596 54292 15598
rect 53340 15260 53396 15316
rect 53228 14642 53284 14644
rect 53228 14590 53230 14642
rect 53230 14590 53282 14642
rect 53282 14590 53284 14642
rect 53228 14588 53284 14590
rect 52444 13804 52500 13860
rect 49980 12626 50036 12628
rect 49980 12574 49982 12626
rect 49982 12574 50034 12626
rect 50034 12574 50036 12626
rect 49980 12572 50036 12574
rect 47068 12460 47124 12516
rect 47964 12460 48020 12516
rect 50556 12122 50612 12124
rect 50556 12070 50558 12122
rect 50558 12070 50610 12122
rect 50610 12070 50612 12122
rect 50556 12068 50612 12070
rect 50660 12122 50716 12124
rect 50660 12070 50662 12122
rect 50662 12070 50714 12122
rect 50714 12070 50716 12122
rect 50660 12068 50716 12070
rect 50764 12122 50820 12124
rect 50764 12070 50766 12122
rect 50766 12070 50818 12122
rect 50818 12070 50820 12122
rect 50764 12068 50820 12070
rect 46620 11730 46676 11732
rect 46620 11678 46622 11730
rect 46622 11678 46674 11730
rect 46674 11678 46676 11730
rect 46620 11676 46676 11678
rect 48076 10444 48132 10500
rect 42028 8706 42084 8708
rect 42028 8654 42030 8706
rect 42030 8654 42082 8706
rect 42082 8654 42084 8706
rect 42028 8652 42084 8654
rect 50556 10106 50612 10108
rect 50556 10054 50558 10106
rect 50558 10054 50610 10106
rect 50610 10054 50612 10106
rect 50556 10052 50612 10054
rect 50660 10106 50716 10108
rect 50660 10054 50662 10106
rect 50662 10054 50714 10106
rect 50714 10054 50716 10106
rect 50660 10052 50716 10054
rect 50764 10106 50820 10108
rect 50764 10054 50766 10106
rect 50766 10054 50818 10106
rect 50818 10054 50820 10106
rect 50764 10052 50820 10054
rect 43260 8594 43316 8596
rect 43260 8542 43262 8594
rect 43262 8542 43314 8594
rect 43314 8542 43316 8594
rect 43260 8540 43316 8542
rect 41468 8428 41524 8484
rect 41916 8316 41972 8372
rect 50556 8090 50612 8092
rect 50556 8038 50558 8090
rect 50558 8038 50610 8090
rect 50610 8038 50612 8090
rect 50556 8036 50612 8038
rect 50660 8090 50716 8092
rect 50660 8038 50662 8090
rect 50662 8038 50714 8090
rect 50714 8038 50716 8090
rect 50660 8036 50716 8038
rect 50764 8090 50820 8092
rect 50764 8038 50766 8090
rect 50766 8038 50818 8090
rect 50818 8038 50820 8090
rect 50764 8036 50820 8038
rect 33740 7586 33796 7588
rect 33740 7534 33742 7586
rect 33742 7534 33794 7586
rect 33794 7534 33796 7586
rect 33740 7532 33796 7534
rect 33628 6578 33684 6580
rect 33628 6526 33630 6578
rect 33630 6526 33682 6578
rect 33682 6526 33684 6578
rect 33628 6524 33684 6526
rect 33852 6636 33908 6692
rect 34972 6466 35028 6468
rect 34972 6414 34974 6466
rect 34974 6414 35026 6466
rect 35026 6414 35028 6466
rect 34972 6412 35028 6414
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 50556 6074 50612 6076
rect 50556 6022 50558 6074
rect 50558 6022 50610 6074
rect 50610 6022 50612 6074
rect 50556 6020 50612 6022
rect 50660 6074 50716 6076
rect 50660 6022 50662 6074
rect 50662 6022 50714 6074
rect 50714 6022 50716 6074
rect 50660 6020 50716 6022
rect 50764 6074 50820 6076
rect 50764 6022 50766 6074
rect 50766 6022 50818 6074
rect 50818 6022 50820 6074
rect 50764 6020 50820 6022
rect 35196 5404 35252 5460
rect 36092 5458 36148 5460
rect 36092 5406 36094 5458
rect 36094 5406 36146 5458
rect 36146 5406 36148 5458
rect 36092 5404 36148 5406
rect 35196 5066 35252 5068
rect 35196 5014 35198 5066
rect 35198 5014 35250 5066
rect 35250 5014 35252 5066
rect 35196 5012 35252 5014
rect 35300 5066 35356 5068
rect 35300 5014 35302 5066
rect 35302 5014 35354 5066
rect 35354 5014 35356 5066
rect 35300 5012 35356 5014
rect 35404 5066 35460 5068
rect 35404 5014 35406 5066
rect 35406 5014 35458 5066
rect 35458 5014 35460 5066
rect 35404 5012 35460 5014
rect 19836 4058 19892 4060
rect 19836 4006 19838 4058
rect 19838 4006 19890 4058
rect 19890 4006 19892 4058
rect 19836 4004 19892 4006
rect 19940 4058 19996 4060
rect 19940 4006 19942 4058
rect 19942 4006 19994 4058
rect 19994 4006 19996 4058
rect 19940 4004 19996 4006
rect 20044 4058 20100 4060
rect 20044 4006 20046 4058
rect 20046 4006 20098 4058
rect 20098 4006 20100 4058
rect 20044 4004 20100 4006
rect 50556 4058 50612 4060
rect 50556 4006 50558 4058
rect 50558 4006 50610 4058
rect 50610 4006 50612 4058
rect 50556 4004 50612 4006
rect 50660 4058 50716 4060
rect 50660 4006 50662 4058
rect 50662 4006 50714 4058
rect 50714 4006 50716 4058
rect 50660 4004 50716 4006
rect 50764 4058 50820 4060
rect 50764 4006 50766 4058
rect 50766 4006 50818 4058
rect 50818 4006 50820 4058
rect 50764 4004 50820 4006
<< metal3 >>
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 4466 55412 4476 55468
rect 4532 55412 4580 55468
rect 4636 55412 4684 55468
rect 4740 55412 4750 55468
rect 35186 55412 35196 55468
rect 35252 55412 35300 55468
rect 35356 55412 35404 55468
rect 35460 55412 35470 55468
rect 19826 54404 19836 54460
rect 19892 54404 19940 54460
rect 19996 54404 20044 54460
rect 20100 54404 20110 54460
rect 50546 54404 50556 54460
rect 50612 54404 50660 54460
rect 50716 54404 50764 54460
rect 50820 54404 50830 54460
rect 59200 53844 60000 53872
rect 55234 53788 55244 53844
rect 55300 53788 60000 53844
rect 59200 53760 60000 53788
rect 4466 53396 4476 53452
rect 4532 53396 4580 53452
rect 4636 53396 4684 53452
rect 4740 53396 4750 53452
rect 35186 53396 35196 53452
rect 35252 53396 35300 53452
rect 35356 53396 35404 53452
rect 35460 53396 35470 53452
rect 19826 52388 19836 52444
rect 19892 52388 19940 52444
rect 19996 52388 20044 52444
rect 20100 52388 20110 52444
rect 50546 52388 50556 52444
rect 50612 52388 50660 52444
rect 50716 52388 50764 52444
rect 50820 52388 50830 52444
rect 3388 52108 5852 52164
rect 5908 52108 5918 52164
rect 0 51828 800 51856
rect 3388 51828 3444 52108
rect 0 51772 3444 51828
rect 0 51744 800 51772
rect 4466 51380 4476 51436
rect 4532 51380 4580 51436
rect 4636 51380 4684 51436
rect 4740 51380 4750 51436
rect 35186 51380 35196 51436
rect 35252 51380 35300 51436
rect 35356 51380 35404 51436
rect 35460 51380 35470 51436
rect 19826 50372 19836 50428
rect 19892 50372 19940 50428
rect 19996 50372 20044 50428
rect 20100 50372 20110 50428
rect 50546 50372 50556 50428
rect 50612 50372 50660 50428
rect 50716 50372 50764 50428
rect 50820 50372 50830 50428
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 36978 48972 36988 49028
rect 37044 48972 37436 49028
rect 37492 48972 40348 49028
rect 40404 48972 41692 49028
rect 41748 48972 42364 49028
rect 42420 48972 43708 49028
rect 31266 48860 31276 48916
rect 31332 48860 32732 48916
rect 32788 48860 32798 48916
rect 41234 48860 41244 48916
rect 41300 48860 41804 48916
rect 41860 48860 42140 48916
rect 42196 48860 43484 48916
rect 43540 48860 43550 48916
rect 43652 48860 43708 48972
rect 43764 48860 43774 48916
rect 30818 48748 30828 48804
rect 30884 48748 31948 48804
rect 32004 48748 32014 48804
rect 40348 48748 40796 48804
rect 40852 48748 41356 48804
rect 41412 48748 42812 48804
rect 42868 48748 42878 48804
rect 40348 48692 40404 48748
rect 40002 48636 40012 48692
rect 40068 48636 40404 48692
rect 19826 48356 19836 48412
rect 19892 48356 19940 48412
rect 19996 48356 20044 48412
rect 20100 48356 20110 48412
rect 50546 48356 50556 48412
rect 50612 48356 50660 48412
rect 50716 48356 50764 48412
rect 50820 48356 50830 48412
rect 24658 47740 24668 47796
rect 24724 47740 26572 47796
rect 26628 47740 26638 47796
rect 36306 47740 36316 47796
rect 36372 47740 37100 47796
rect 37156 47740 38108 47796
rect 38164 47740 38174 47796
rect 4466 47348 4476 47404
rect 4532 47348 4580 47404
rect 4636 47348 4684 47404
rect 4740 47348 4750 47404
rect 35186 47348 35196 47404
rect 35252 47348 35300 47404
rect 35356 47348 35404 47404
rect 35460 47348 35470 47404
rect 26562 47068 26572 47124
rect 26628 47068 26852 47124
rect 26796 47012 26852 47068
rect 3938 46956 3948 47012
rect 4004 46956 4508 47012
rect 4564 46956 5628 47012
rect 5684 46956 5694 47012
rect 26796 46956 27580 47012
rect 27636 46956 27646 47012
rect 38994 46844 39004 46900
rect 39060 46844 40236 46900
rect 40292 46844 41132 46900
rect 41188 46844 41198 46900
rect 27794 46620 27804 46676
rect 27860 46620 29708 46676
rect 29764 46620 31500 46676
rect 31556 46620 32620 46676
rect 32676 46620 32686 46676
rect 39890 46620 39900 46676
rect 39956 46620 40684 46676
rect 40740 46620 41244 46676
rect 41300 46620 41580 46676
rect 41636 46620 41646 46676
rect 43026 46508 43036 46564
rect 43092 46508 44044 46564
rect 44100 46508 44110 46564
rect 19826 46340 19836 46396
rect 19892 46340 19940 46396
rect 19996 46340 20044 46396
rect 20100 46340 20110 46396
rect 50546 46340 50556 46396
rect 50612 46340 50660 46396
rect 50716 46340 50764 46396
rect 50820 46340 50830 46396
rect 40114 46172 40124 46228
rect 40180 46172 40908 46228
rect 40964 46172 40974 46228
rect 27570 45948 27580 46004
rect 27636 45948 28588 46004
rect 28644 45948 28654 46004
rect 35074 45836 35084 45892
rect 35140 45836 35980 45892
rect 36036 45836 36046 45892
rect 4162 45724 4172 45780
rect 4228 45724 6188 45780
rect 6244 45724 7196 45780
rect 7252 45724 9660 45780
rect 9716 45724 9726 45780
rect 24994 45724 25004 45780
rect 25060 45724 26460 45780
rect 26516 45724 29260 45780
rect 29316 45724 29326 45780
rect 31938 45724 31948 45780
rect 32004 45724 33292 45780
rect 33348 45724 34636 45780
rect 34692 45724 35868 45780
rect 35924 45724 36092 45780
rect 36148 45724 36158 45780
rect 8764 45668 8820 45724
rect 5730 45612 5740 45668
rect 5796 45612 7644 45668
rect 7700 45612 7710 45668
rect 8754 45612 8764 45668
rect 8820 45612 8830 45668
rect 6066 45500 6076 45556
rect 6132 45500 8316 45556
rect 8372 45500 8382 45556
rect 30930 45388 30940 45444
rect 30996 45388 31948 45444
rect 38444 45388 39004 45444
rect 39060 45388 39070 45444
rect 4466 45332 4476 45388
rect 4532 45332 4580 45388
rect 4636 45332 4684 45388
rect 4740 45332 4750 45388
rect 31892 45332 31948 45388
rect 35186 45332 35196 45388
rect 35252 45332 35300 45388
rect 35356 45332 35404 45388
rect 35460 45332 35470 45388
rect 38444 45332 38500 45388
rect 1698 45276 1708 45332
rect 1764 45276 3052 45332
rect 3108 45276 4172 45332
rect 4228 45276 4238 45332
rect 30258 45276 30268 45332
rect 30324 45276 31276 45332
rect 31332 45276 31342 45332
rect 31892 45276 33180 45332
rect 33236 45276 33246 45332
rect 38322 45276 38332 45332
rect 38388 45276 38500 45332
rect 41458 45276 41468 45332
rect 41524 45276 42924 45332
rect 42980 45276 42990 45332
rect 11666 45052 11676 45108
rect 11732 45052 12796 45108
rect 12852 45052 12862 45108
rect 9538 44940 9548 44996
rect 9604 44940 10220 44996
rect 10276 44940 11564 44996
rect 11620 44940 11630 44996
rect 22194 44940 22204 44996
rect 22260 44940 26404 44996
rect 35970 44940 35980 44996
rect 36036 44940 37660 44996
rect 37716 44940 38780 44996
rect 38836 44940 38846 44996
rect 26348 44884 26404 44940
rect 6626 44828 6636 44884
rect 6692 44828 9660 44884
rect 9716 44828 9726 44884
rect 22754 44828 22764 44884
rect 22820 44828 23436 44884
rect 23492 44828 23502 44884
rect 26338 44828 26348 44884
rect 26404 44828 27804 44884
rect 27860 44828 27870 44884
rect 28130 44828 28140 44884
rect 28196 44828 29484 44884
rect 29540 44828 29932 44884
rect 29988 44828 31948 44884
rect 32004 44828 32014 44884
rect 2370 44604 2380 44660
rect 2436 44604 3388 44660
rect 3444 44604 6076 44660
rect 6132 44604 6142 44660
rect 9202 44604 9212 44660
rect 9268 44604 10332 44660
rect 10388 44604 10398 44660
rect 35634 44604 35644 44660
rect 35700 44604 36428 44660
rect 36484 44604 36494 44660
rect 37202 44604 37212 44660
rect 37268 44604 41132 44660
rect 41188 44604 45164 44660
rect 45220 44604 45500 44660
rect 45556 44604 45566 44660
rect 0 44436 800 44464
rect 0 44380 1820 44436
rect 1876 44380 1886 44436
rect 0 44352 800 44380
rect 19826 44324 19836 44380
rect 19892 44324 19940 44380
rect 19996 44324 20044 44380
rect 20100 44324 20110 44380
rect 50546 44324 50556 44380
rect 50612 44324 50660 44380
rect 50716 44324 50764 44380
rect 50820 44324 50830 44380
rect 8530 44044 8540 44100
rect 8596 44044 9884 44100
rect 9940 44044 12348 44100
rect 12404 44044 12414 44100
rect 23986 44044 23996 44100
rect 24052 44044 24668 44100
rect 24724 44044 27244 44100
rect 27300 44044 28644 44100
rect 33170 44044 33180 44100
rect 33236 44044 34412 44100
rect 34468 44044 35644 44100
rect 35700 44044 35710 44100
rect 28588 43988 28644 44044
rect 10882 43932 10892 43988
rect 10948 43932 14476 43988
rect 14532 43932 14542 43988
rect 27682 43932 27692 43988
rect 27748 43932 28140 43988
rect 28196 43932 28206 43988
rect 28578 43932 28588 43988
rect 28644 43932 28812 43988
rect 28868 43932 29932 43988
rect 29988 43932 29998 43988
rect 12786 43820 12796 43876
rect 12852 43820 14588 43876
rect 14644 43820 14654 43876
rect 22194 43820 22204 43876
rect 22260 43820 23548 43876
rect 23604 43820 23614 43876
rect 31892 43820 33516 43876
rect 33572 43820 35532 43876
rect 35588 43820 35598 43876
rect 36754 43820 36764 43876
rect 36820 43820 37996 43876
rect 38052 43820 39004 43876
rect 39060 43820 39070 43876
rect 40002 43820 40012 43876
rect 40068 43820 41244 43876
rect 41300 43820 41310 43876
rect 31892 43764 31948 43820
rect 20178 43708 20188 43764
rect 20244 43708 21644 43764
rect 21700 43708 22540 43764
rect 22596 43708 22606 43764
rect 23874 43708 23884 43764
rect 23940 43708 26684 43764
rect 26740 43708 26750 43764
rect 31266 43708 31276 43764
rect 31332 43708 31948 43764
rect 32274 43708 32284 43764
rect 32340 43708 33180 43764
rect 33236 43708 33246 43764
rect 36082 43708 36092 43764
rect 36148 43708 37100 43764
rect 37156 43708 37166 43764
rect 43138 43708 43148 43764
rect 43204 43708 45724 43764
rect 45780 43708 46508 43764
rect 46564 43708 46574 43764
rect 12338 43596 12348 43652
rect 12404 43596 13468 43652
rect 13524 43596 13534 43652
rect 23090 43596 23100 43652
rect 23156 43596 24668 43652
rect 24724 43596 24734 43652
rect 45490 43596 45500 43652
rect 45556 43596 46732 43652
rect 46788 43596 47292 43652
rect 47348 43596 47358 43652
rect 22530 43484 22540 43540
rect 22596 43484 23884 43540
rect 23940 43484 23950 43540
rect 46050 43484 46060 43540
rect 46116 43484 47404 43540
rect 47460 43484 47964 43540
rect 48020 43484 48030 43540
rect 4466 43316 4476 43372
rect 4532 43316 4580 43372
rect 4636 43316 4684 43372
rect 4740 43316 4750 43372
rect 35186 43316 35196 43372
rect 35252 43316 35300 43372
rect 35356 43316 35404 43372
rect 35460 43316 35470 43372
rect 1922 43148 1932 43204
rect 1988 43148 2716 43204
rect 2772 43148 5628 43204
rect 5684 43148 5694 43204
rect 10770 43148 10780 43204
rect 10836 43148 11452 43204
rect 11508 43148 13468 43204
rect 13524 43148 13534 43204
rect 4946 42812 4956 42868
rect 5012 42812 6188 42868
rect 6244 42812 6254 42868
rect 27794 42812 27804 42868
rect 27860 42812 28588 42868
rect 28644 42812 28654 42868
rect 47954 42812 47964 42868
rect 48020 42812 49420 42868
rect 49476 42812 49486 42868
rect 20132 42700 22316 42756
rect 22372 42700 23100 42756
rect 23156 42700 23436 42756
rect 23492 42700 23502 42756
rect 31892 42700 33292 42756
rect 33348 42700 35308 42756
rect 35364 42700 35374 42756
rect 47506 42700 47516 42756
rect 47572 42700 48860 42756
rect 48916 42700 48926 42756
rect 13346 42588 13356 42644
rect 13412 42588 16716 42644
rect 16772 42588 16782 42644
rect 20132 42532 20188 42700
rect 31892 42644 31948 42700
rect 21410 42588 21420 42644
rect 21476 42588 22204 42644
rect 22260 42588 22764 42644
rect 22820 42588 22830 42644
rect 28018 42588 28028 42644
rect 28084 42588 29820 42644
rect 29876 42588 31948 42644
rect 51650 42588 51660 42644
rect 51716 42588 53340 42644
rect 53396 42588 53406 42644
rect 17836 42476 19852 42532
rect 19908 42476 20188 42532
rect 17836 42420 17892 42476
rect 17826 42364 17836 42420
rect 17892 42364 17902 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 45378 42140 45388 42196
rect 45444 42140 46732 42196
rect 46788 42140 47740 42196
rect 47796 42140 49084 42196
rect 49140 42140 49756 42196
rect 49812 42140 52108 42196
rect 52164 42140 53788 42196
rect 53844 42140 53854 42196
rect 20132 42028 21420 42084
rect 21476 42028 21486 42084
rect 26898 42028 26908 42084
rect 26964 42028 28028 42084
rect 28084 42028 28094 42084
rect 48850 42028 48860 42084
rect 48916 42028 49308 42084
rect 49364 42028 49868 42084
rect 49924 42028 51660 42084
rect 51716 42028 51726 42084
rect 51986 42028 51996 42084
rect 52052 42028 52780 42084
rect 52836 42028 52846 42084
rect 20132 41972 20188 42028
rect 2370 41916 2380 41972
rect 2436 41916 3388 41972
rect 3444 41916 3454 41972
rect 18498 41916 18508 41972
rect 18564 41916 20188 41972
rect 20514 41916 20524 41972
rect 20580 41916 21980 41972
rect 22036 41916 22046 41972
rect 23538 41916 23548 41972
rect 23604 41916 23614 41972
rect 23762 41916 23772 41972
rect 23828 41916 26124 41972
rect 26180 41916 26190 41972
rect 26338 41916 26348 41972
rect 26404 41916 27132 41972
rect 27188 41916 27198 41972
rect 32050 41916 32060 41972
rect 32116 41916 33404 41972
rect 33460 41916 33470 41972
rect 34626 41916 34636 41972
rect 34692 41916 41132 41972
rect 41188 41916 42588 41972
rect 42644 41916 42654 41972
rect 43922 41916 43932 41972
rect 43988 41916 44380 41972
rect 44436 41916 44446 41972
rect 44706 41916 44716 41972
rect 44772 41916 45388 41972
rect 45444 41916 45454 41972
rect 50866 41916 50876 41972
rect 50932 41916 53116 41972
rect 53172 41916 53182 41972
rect 23548 41860 23604 41916
rect 33404 41860 33460 41916
rect 23548 41804 30044 41860
rect 30100 41804 30110 41860
rect 33404 41804 37436 41860
rect 37492 41804 40012 41860
rect 40068 41804 40078 41860
rect 40898 41804 40908 41860
rect 40964 41804 44268 41860
rect 44324 41804 44940 41860
rect 44996 41804 45006 41860
rect 47506 41804 47516 41860
rect 47572 41804 48636 41860
rect 48692 41804 49196 41860
rect 49252 41804 49262 41860
rect 51090 41804 51100 41860
rect 51156 41804 54348 41860
rect 54404 41804 54414 41860
rect 40908 41748 40964 41804
rect 26786 41692 26796 41748
rect 26852 41692 30492 41748
rect 30548 41692 30558 41748
rect 38658 41692 38668 41748
rect 38724 41692 39900 41748
rect 39956 41692 40964 41748
rect 44482 41692 44492 41748
rect 44548 41692 45612 41748
rect 45668 41692 45678 41748
rect 50866 41692 50876 41748
rect 50932 41692 51212 41748
rect 51268 41692 51278 41748
rect 5730 41580 5740 41636
rect 5796 41580 6972 41636
rect 7028 41580 7038 41636
rect 9650 41580 9660 41636
rect 9716 41580 11340 41636
rect 11396 41580 14364 41636
rect 14420 41580 14430 41636
rect 26002 41580 26012 41636
rect 26068 41580 27020 41636
rect 27076 41580 27086 41636
rect 37538 41580 37548 41636
rect 37604 41580 38892 41636
rect 38948 41580 41580 41636
rect 41636 41580 43484 41636
rect 43540 41580 43550 41636
rect 49410 41580 49420 41636
rect 49476 41580 51996 41636
rect 52052 41580 52062 41636
rect 1810 41468 1820 41524
rect 1876 41468 4396 41524
rect 4452 41468 5628 41524
rect 5684 41468 5694 41524
rect 4466 41300 4476 41356
rect 4532 41300 4580 41356
rect 4636 41300 4684 41356
rect 4740 41300 4750 41356
rect 35186 41300 35196 41356
rect 35252 41300 35300 41356
rect 35356 41300 35404 41356
rect 35460 41300 35470 41356
rect 32722 41132 32732 41188
rect 32788 41132 34972 41188
rect 35028 41132 35038 41188
rect 18956 41020 21308 41076
rect 21364 41020 21374 41076
rect 1698 40908 1708 40964
rect 1764 40908 2380 40964
rect 2436 40908 6076 40964
rect 6132 40908 6142 40964
rect 18956 40852 19012 41020
rect 30370 40908 30380 40964
rect 30436 40908 37324 40964
rect 37380 40908 37390 40964
rect 37874 40908 37884 40964
rect 37940 40908 40348 40964
rect 40404 40908 43036 40964
rect 43092 40908 43932 40964
rect 43988 40908 43998 40964
rect 17602 40796 17612 40852
rect 17668 40796 17948 40852
rect 18004 40796 18172 40852
rect 18228 40796 18956 40852
rect 19012 40796 19022 40852
rect 20178 40796 20188 40852
rect 20244 40796 20748 40852
rect 20804 40796 29484 40852
rect 29540 40796 34468 40852
rect 43474 40796 43484 40852
rect 43540 40796 43708 40852
rect 44034 40796 44044 40852
rect 44100 40796 45388 40852
rect 45444 40796 45454 40852
rect 46722 40796 46732 40852
rect 46788 40796 47516 40852
rect 47572 40796 47582 40852
rect 34412 40740 34468 40796
rect 10210 40684 10220 40740
rect 10276 40684 10780 40740
rect 10836 40684 13468 40740
rect 13524 40684 13534 40740
rect 22530 40684 22540 40740
rect 22596 40684 23100 40740
rect 23156 40684 23884 40740
rect 23940 40684 23950 40740
rect 29810 40684 29820 40740
rect 29876 40684 31164 40740
rect 31220 40684 32508 40740
rect 32564 40684 32574 40740
rect 34402 40684 34412 40740
rect 34468 40684 36764 40740
rect 36820 40684 38556 40740
rect 38612 40684 41244 40740
rect 41300 40684 42700 40740
rect 42756 40684 42766 40740
rect 43652 40628 43708 40796
rect 44044 40628 44100 40796
rect 4946 40572 4956 40628
rect 5012 40572 6188 40628
rect 6244 40572 6254 40628
rect 8372 40572 9324 40628
rect 9380 40572 10444 40628
rect 10500 40572 10510 40628
rect 12786 40572 12796 40628
rect 12852 40572 13580 40628
rect 13636 40572 13646 40628
rect 25106 40572 25116 40628
rect 25172 40572 29372 40628
rect 29428 40572 29438 40628
rect 43652 40572 44100 40628
rect 1810 40348 1820 40404
rect 1876 40348 3052 40404
rect 3108 40348 4060 40404
rect 4116 40348 4126 40404
rect 8372 40292 8428 40572
rect 21410 40460 21420 40516
rect 21476 40460 29260 40516
rect 29316 40460 30716 40516
rect 30772 40460 37100 40516
rect 37156 40460 37660 40516
rect 37716 40460 37726 40516
rect 26562 40348 26572 40404
rect 26628 40348 27020 40404
rect 27076 40348 27086 40404
rect 29810 40348 29820 40404
rect 29876 40348 34076 40404
rect 34132 40348 34142 40404
rect 54674 40348 54684 40404
rect 54740 40348 55580 40404
rect 55636 40348 55646 40404
rect 19826 40292 19836 40348
rect 19892 40292 19940 40348
rect 19996 40292 20044 40348
rect 20100 40292 20110 40348
rect 50546 40292 50556 40348
rect 50612 40292 50660 40348
rect 50716 40292 50764 40348
rect 50820 40292 50830 40348
rect 6850 40236 6860 40292
rect 6916 40236 8428 40292
rect 30258 40236 30268 40292
rect 30324 40236 31612 40292
rect 31668 40236 32508 40292
rect 32564 40236 33068 40292
rect 33124 40236 33134 40292
rect 46722 40124 46732 40180
rect 46788 40124 53788 40180
rect 53844 40124 53854 40180
rect 24658 40012 24668 40068
rect 24724 40012 25452 40068
rect 25508 40012 25518 40068
rect 27122 40012 27132 40068
rect 27188 40012 28476 40068
rect 28532 40012 28542 40068
rect 39890 40012 39900 40068
rect 39956 40012 40908 40068
rect 40964 40012 40974 40068
rect 42354 40012 42364 40068
rect 42420 40012 43708 40068
rect 43764 40012 43774 40068
rect 3826 39900 3836 39956
rect 3892 39900 4956 39956
rect 5012 39900 5022 39956
rect 24210 39900 24220 39956
rect 24276 39900 25116 39956
rect 25172 39900 25182 39956
rect 27682 39900 27692 39956
rect 27748 39900 29260 39956
rect 29316 39900 29326 39956
rect 44930 39900 44940 39956
rect 44996 39900 45724 39956
rect 45780 39900 45790 39956
rect 46620 39900 48748 39956
rect 48804 39900 49196 39956
rect 49252 39900 49868 39956
rect 49924 39900 50988 39956
rect 51044 39900 51054 39956
rect 53218 39900 53228 39956
rect 53284 39900 54572 39956
rect 54628 39900 54638 39956
rect 46620 39844 46676 39900
rect 11330 39788 11340 39844
rect 11396 39788 11676 39844
rect 11732 39788 12684 39844
rect 12740 39788 12750 39844
rect 21634 39788 21644 39844
rect 21700 39788 22652 39844
rect 22708 39788 22718 39844
rect 26450 39788 26460 39844
rect 26516 39788 27580 39844
rect 27636 39788 27646 39844
rect 35522 39788 35532 39844
rect 35588 39788 41916 39844
rect 41972 39788 41982 39844
rect 44482 39788 44492 39844
rect 44548 39788 45388 39844
rect 45444 39788 46676 39844
rect 46834 39788 46844 39844
rect 46900 39788 50540 39844
rect 50596 39788 50606 39844
rect 51986 39788 51996 39844
rect 52052 39788 53004 39844
rect 53060 39788 53070 39844
rect 53554 39788 53564 39844
rect 53620 39788 54012 39844
rect 54068 39788 55356 39844
rect 55412 39788 56140 39844
rect 56196 39788 56206 39844
rect 0 39732 800 39760
rect 44492 39732 44548 39788
rect 0 39676 4284 39732
rect 4340 39676 4350 39732
rect 16482 39676 16492 39732
rect 16548 39676 18396 39732
rect 18452 39676 18462 39732
rect 36418 39676 36428 39732
rect 36484 39676 37884 39732
rect 37940 39676 37950 39732
rect 38210 39676 38220 39732
rect 38276 39676 44548 39732
rect 53004 39732 53060 39788
rect 53004 39676 54348 39732
rect 54404 39676 56476 39732
rect 56532 39676 57148 39732
rect 57204 39676 57214 39732
rect 0 39648 800 39676
rect 12786 39564 12796 39620
rect 12852 39564 13916 39620
rect 13972 39564 13982 39620
rect 35634 39564 35644 39620
rect 35700 39564 36988 39620
rect 37044 39564 37054 39620
rect 4466 39284 4476 39340
rect 4532 39284 4580 39340
rect 4636 39284 4684 39340
rect 4740 39284 4750 39340
rect 35186 39284 35196 39340
rect 35252 39284 35300 39340
rect 35356 39284 35404 39340
rect 35460 39284 35470 39340
rect 27122 39228 27132 39284
rect 27188 39228 28364 39284
rect 28420 39228 28430 39284
rect 4946 39116 4956 39172
rect 5012 39116 8316 39172
rect 8372 39116 8382 39172
rect 0 39060 800 39088
rect 0 39004 17388 39060
rect 17444 39004 17454 39060
rect 18722 39004 18732 39060
rect 18788 39004 20412 39060
rect 20468 39004 21644 39060
rect 21700 39004 21710 39060
rect 39218 39004 39228 39060
rect 39284 39004 40460 39060
rect 40516 39004 41356 39060
rect 41412 39004 41422 39060
rect 0 38976 800 39004
rect 28354 38892 28364 38948
rect 28420 38892 30044 38948
rect 30100 38892 30110 38948
rect 30594 38892 30604 38948
rect 30660 38892 33628 38948
rect 33684 38892 34412 38948
rect 34468 38892 34748 38948
rect 34804 38892 36092 38948
rect 36148 38892 36158 38948
rect 37538 38892 37548 38948
rect 37604 38892 38108 38948
rect 38164 38892 41132 38948
rect 41188 38892 41198 38948
rect 19954 38780 19964 38836
rect 20020 38780 21868 38836
rect 21924 38780 21934 38836
rect 25106 38780 25116 38836
rect 25172 38780 27580 38836
rect 27636 38780 27646 38836
rect 44930 38780 44940 38836
rect 44996 38780 46508 38836
rect 46564 38780 46574 38836
rect 53666 38780 53676 38836
rect 53732 38780 55468 38836
rect 3826 38668 3836 38724
rect 3892 38668 4620 38724
rect 4676 38668 6076 38724
rect 6132 38668 6860 38724
rect 6916 38668 6926 38724
rect 12226 38668 12236 38724
rect 12292 38668 13468 38724
rect 13524 38668 13534 38724
rect 17826 38668 17836 38724
rect 17892 38668 18508 38724
rect 18564 38668 22988 38724
rect 23044 38668 23054 38724
rect 37874 38668 37884 38724
rect 37940 38668 38892 38724
rect 38948 38668 41244 38724
rect 41300 38668 41310 38724
rect 42018 38668 42028 38724
rect 42084 38668 47180 38724
rect 47236 38668 47246 38724
rect 48290 38668 48300 38724
rect 48356 38668 50540 38724
rect 50596 38668 51772 38724
rect 51828 38668 51838 38724
rect 55412 38612 55468 38780
rect 16818 38556 16828 38612
rect 16884 38556 20412 38612
rect 20468 38556 21532 38612
rect 21588 38556 21598 38612
rect 55412 38556 56700 38612
rect 56756 38556 57036 38612
rect 57092 38556 57102 38612
rect 26852 38444 34524 38500
rect 34580 38444 34590 38500
rect 19826 38276 19836 38332
rect 19892 38276 19940 38332
rect 19996 38276 20044 38332
rect 20100 38276 20110 38332
rect 26852 38276 26908 38444
rect 28242 38332 28252 38388
rect 28308 38332 28318 38388
rect 4834 38220 4844 38276
rect 4900 38220 5516 38276
rect 5572 38220 7084 38276
rect 7140 38220 7150 38276
rect 26002 38220 26012 38276
rect 26068 38220 26908 38276
rect 6290 38108 6300 38164
rect 6356 38108 7532 38164
rect 7588 38108 8876 38164
rect 8932 38108 8942 38164
rect 17042 37996 17052 38052
rect 17108 37996 17948 38052
rect 18004 37996 19068 38052
rect 19124 37996 19134 38052
rect 28252 37940 28308 38332
rect 50546 38276 50556 38332
rect 50612 38276 50660 38332
rect 50716 38276 50764 38332
rect 50820 38276 50830 38332
rect 37762 38220 37772 38276
rect 37828 38220 38556 38276
rect 38612 38220 38622 38276
rect 37874 37996 37884 38052
rect 37940 37996 40348 38052
rect 40404 37996 40414 38052
rect 17490 37884 17500 37940
rect 17556 37884 20412 37940
rect 20468 37884 21308 37940
rect 21364 37884 22092 37940
rect 22148 37884 23548 37940
rect 23604 37884 23614 37940
rect 25778 37884 25788 37940
rect 25844 37884 28308 37940
rect 45938 37884 45948 37940
rect 46004 37884 47292 37940
rect 47348 37884 47358 37940
rect 4274 37772 4284 37828
rect 4340 37772 18396 37828
rect 18452 37772 18462 37828
rect 19394 37772 19404 37828
rect 19460 37772 19964 37828
rect 20020 37772 20636 37828
rect 20692 37772 20702 37828
rect 39778 37772 39788 37828
rect 39844 37772 40908 37828
rect 40964 37772 40974 37828
rect 42466 37772 42476 37828
rect 42532 37772 43484 37828
rect 43540 37772 44492 37828
rect 44548 37772 44828 37828
rect 44884 37772 45276 37828
rect 45332 37772 45342 37828
rect 50372 37772 51548 37828
rect 51604 37772 51614 37828
rect 0 37716 800 37744
rect 18396 37716 18452 37772
rect 50372 37716 50428 37772
rect 0 37660 16828 37716
rect 16884 37660 16894 37716
rect 18396 37660 21084 37716
rect 21140 37660 22204 37716
rect 22260 37660 22652 37716
rect 22708 37660 22718 37716
rect 24882 37660 24892 37716
rect 24948 37660 26348 37716
rect 26404 37660 27244 37716
rect 27300 37660 27310 37716
rect 32498 37660 32508 37716
rect 32564 37660 35308 37716
rect 35364 37660 35374 37716
rect 42578 37660 42588 37716
rect 42644 37660 48860 37716
rect 48916 37660 50092 37716
rect 50148 37660 50428 37716
rect 55570 37660 55580 37716
rect 55636 37660 57036 37716
rect 57092 37660 57596 37716
rect 57652 37660 57662 37716
rect 0 37632 800 37660
rect 40338 37548 40348 37604
rect 40404 37548 42252 37604
rect 42308 37548 43036 37604
rect 43092 37548 43102 37604
rect 53666 37436 53676 37492
rect 53732 37436 54348 37492
rect 54404 37436 54414 37492
rect 4466 37268 4476 37324
rect 4532 37268 4580 37324
rect 4636 37268 4684 37324
rect 4740 37268 4750 37324
rect 35186 37268 35196 37324
rect 35252 37268 35300 37324
rect 35356 37268 35404 37324
rect 35460 37268 35470 37324
rect 4498 37100 4508 37156
rect 4564 37100 6636 37156
rect 6692 37100 6702 37156
rect 0 37044 800 37072
rect 0 36988 18844 37044
rect 18900 36988 19964 37044
rect 20020 36988 20412 37044
rect 20468 36988 21756 37044
rect 21812 36988 21822 37044
rect 51426 36988 51436 37044
rect 51492 36988 53788 37044
rect 53844 36988 55356 37044
rect 55412 36988 57148 37044
rect 57204 36988 57484 37044
rect 57540 36988 57550 37044
rect 0 36960 800 36988
rect 21756 36932 21812 36988
rect 7634 36876 7644 36932
rect 7700 36876 8764 36932
rect 8820 36876 8830 36932
rect 13570 36876 13580 36932
rect 13636 36876 14812 36932
rect 14868 36876 14878 36932
rect 19170 36876 19180 36932
rect 19236 36876 20076 36932
rect 20132 36876 21420 36932
rect 21476 36876 21486 36932
rect 21756 36876 21980 36932
rect 22036 36876 22046 36932
rect 50194 36876 50204 36932
rect 50260 36876 51212 36932
rect 51268 36876 54460 36932
rect 54516 36876 54526 36932
rect 14690 36764 14700 36820
rect 14756 36764 15036 36820
rect 15092 36764 15484 36820
rect 15540 36764 15550 36820
rect 19058 36764 19068 36820
rect 19124 36764 29372 36820
rect 29428 36764 30716 36820
rect 30772 36764 30782 36820
rect 44930 36764 44940 36820
rect 44996 36764 46172 36820
rect 46228 36764 47180 36820
rect 47236 36764 47246 36820
rect 48178 36764 48188 36820
rect 48244 36764 50316 36820
rect 50372 36764 51324 36820
rect 51380 36764 51996 36820
rect 52052 36764 52062 36820
rect 17826 36652 17836 36708
rect 17892 36652 18508 36708
rect 18564 36652 18574 36708
rect 21410 36652 21420 36708
rect 21476 36652 21980 36708
rect 22036 36652 22046 36708
rect 22194 36652 22204 36708
rect 22260 36652 22540 36708
rect 22596 36652 25340 36708
rect 25396 36652 25406 36708
rect 27346 36652 27356 36708
rect 27412 36652 29260 36708
rect 29316 36652 29326 36708
rect 43474 36652 43484 36708
rect 43540 36652 44044 36708
rect 44100 36652 46732 36708
rect 46788 36652 46798 36708
rect 47730 36652 47740 36708
rect 47796 36652 49756 36708
rect 49812 36652 50540 36708
rect 50596 36652 50876 36708
rect 50932 36652 50942 36708
rect 55122 36652 55132 36708
rect 55188 36652 55198 36708
rect 55346 36652 55356 36708
rect 55412 36652 56700 36708
rect 56756 36652 57932 36708
rect 57988 36652 57998 36708
rect 55132 36596 55188 36652
rect 4946 36540 4956 36596
rect 5012 36540 6188 36596
rect 6244 36540 6254 36596
rect 8306 36540 8316 36596
rect 8372 36540 11004 36596
rect 11060 36540 11070 36596
rect 15810 36540 15820 36596
rect 15876 36540 18060 36596
rect 18116 36540 18126 36596
rect 21634 36540 21644 36596
rect 21700 36540 23548 36596
rect 23604 36540 24220 36596
rect 24276 36540 25116 36596
rect 25172 36540 25182 36596
rect 36418 36540 36428 36596
rect 36484 36540 37660 36596
rect 37716 36540 37726 36596
rect 43138 36540 43148 36596
rect 43204 36540 43932 36596
rect 43988 36540 43998 36596
rect 51874 36540 51884 36596
rect 51940 36540 54012 36596
rect 54068 36540 54078 36596
rect 55132 36540 56588 36596
rect 56644 36540 56654 36596
rect 9762 36428 9772 36484
rect 9828 36428 13468 36484
rect 13524 36428 13534 36484
rect 51650 36428 51660 36484
rect 51716 36428 53452 36484
rect 53508 36428 55244 36484
rect 55300 36428 55310 36484
rect 0 36372 800 36400
rect 0 36316 4172 36372
rect 4228 36316 4238 36372
rect 0 36288 800 36316
rect 19826 36260 19836 36316
rect 19892 36260 19940 36316
rect 19996 36260 20044 36316
rect 20100 36260 20110 36316
rect 50546 36260 50556 36316
rect 50612 36260 50660 36316
rect 50716 36260 50764 36316
rect 50820 36260 50830 36316
rect 20066 36092 20076 36148
rect 20132 36092 22876 36148
rect 22932 36092 27356 36148
rect 27412 36092 27422 36148
rect 36418 36092 36428 36148
rect 36484 36092 36876 36148
rect 36932 36092 40348 36148
rect 40404 36092 40414 36148
rect 2706 35980 2716 36036
rect 2772 35980 3164 36036
rect 3220 35980 4060 36036
rect 4116 35980 4126 36036
rect 21746 35980 21756 36036
rect 21812 35980 21980 36036
rect 22036 35980 22046 36036
rect 24770 35980 24780 36036
rect 24836 35980 30156 36036
rect 30212 35980 30222 36036
rect 38882 35980 38892 36036
rect 38948 35980 39676 36036
rect 39732 35980 41244 36036
rect 41300 35980 41916 36036
rect 41972 35980 42252 36036
rect 42308 35980 43820 36036
rect 43876 35980 44380 36036
rect 44436 35980 44828 36036
rect 44884 35980 45612 36036
rect 45668 35980 46732 36036
rect 46788 35980 47740 36036
rect 47796 35980 47806 36036
rect 52322 35980 52332 36036
rect 52388 35980 52780 36036
rect 52836 35980 54236 36036
rect 54292 35980 54302 36036
rect 12114 35868 12124 35924
rect 12180 35868 14476 35924
rect 14532 35868 14542 35924
rect 19730 35868 19740 35924
rect 19796 35868 20748 35924
rect 20804 35868 20814 35924
rect 25554 35868 25564 35924
rect 25620 35868 27020 35924
rect 27076 35868 27086 35924
rect 14578 35756 14588 35812
rect 14644 35756 19628 35812
rect 19684 35756 19694 35812
rect 23202 35756 23212 35812
rect 23268 35756 24108 35812
rect 24164 35756 24444 35812
rect 24500 35756 25900 35812
rect 25956 35756 25966 35812
rect 32162 35756 32172 35812
rect 32228 35756 34972 35812
rect 35028 35756 36204 35812
rect 36260 35756 36270 35812
rect 36754 35756 36764 35812
rect 36820 35756 37324 35812
rect 37380 35756 39228 35812
rect 39284 35756 39294 35812
rect 46386 35756 46396 35812
rect 46452 35756 48748 35812
rect 48804 35756 48814 35812
rect 50082 35756 50092 35812
rect 50148 35756 53676 35812
rect 53732 35756 53742 35812
rect 54562 35756 54572 35812
rect 54628 35756 55580 35812
rect 55636 35756 56924 35812
rect 56980 35756 56990 35812
rect 22530 35644 22540 35700
rect 22596 35644 23100 35700
rect 23156 35644 23772 35700
rect 23828 35644 23838 35700
rect 40338 35644 40348 35700
rect 40404 35644 43148 35700
rect 43204 35644 43214 35700
rect 34626 35532 34636 35588
rect 34692 35532 35980 35588
rect 36036 35532 36046 35588
rect 16594 35420 16604 35476
rect 16660 35420 17948 35476
rect 18004 35420 18014 35476
rect 55010 35420 55020 35476
rect 55076 35420 55580 35476
rect 55636 35420 55646 35476
rect 55804 35364 55860 35756
rect 18946 35308 18956 35364
rect 19012 35308 20524 35364
rect 20580 35308 27132 35364
rect 27188 35308 28028 35364
rect 28084 35308 28094 35364
rect 53442 35308 53452 35364
rect 53508 35308 55916 35364
rect 55972 35308 55982 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 4162 34972 4172 35028
rect 4228 34972 19180 35028
rect 19236 34972 20300 35028
rect 20356 34972 22540 35028
rect 22596 34972 22606 35028
rect 2370 34860 2380 34916
rect 2436 34860 3052 34916
rect 3108 34860 5628 34916
rect 5684 34860 5694 34916
rect 16146 34860 16156 34916
rect 16212 34860 19516 34916
rect 19572 34860 19582 34916
rect 35634 34860 35644 34916
rect 35700 34860 37548 34916
rect 37604 34860 39452 34916
rect 39508 34860 39518 34916
rect 40796 34860 42588 34916
rect 42644 34860 43596 34916
rect 43652 34860 43662 34916
rect 50372 34860 51548 34916
rect 51604 34860 51614 34916
rect 40796 34804 40852 34860
rect 50372 34804 50428 34860
rect 22530 34748 22540 34804
rect 22596 34748 23548 34804
rect 23604 34748 23614 34804
rect 32050 34748 32060 34804
rect 32116 34748 32732 34804
rect 32788 34748 32798 34804
rect 36082 34748 36092 34804
rect 36148 34748 37660 34804
rect 37716 34748 40852 34804
rect 41010 34748 41020 34804
rect 41076 34748 41580 34804
rect 41636 34748 42364 34804
rect 42420 34748 44268 34804
rect 44324 34748 45500 34804
rect 45556 34748 45566 34804
rect 46610 34748 46620 34804
rect 46676 34748 47516 34804
rect 47572 34748 49644 34804
rect 49700 34748 50428 34804
rect 51090 34748 51100 34804
rect 51156 34748 53004 34804
rect 53060 34748 53452 34804
rect 53508 34748 53518 34804
rect 4050 34636 4060 34692
rect 4116 34636 4620 34692
rect 4676 34636 5516 34692
rect 5572 34636 5852 34692
rect 5908 34636 8540 34692
rect 8596 34636 9324 34692
rect 9380 34636 9390 34692
rect 9874 34636 9884 34692
rect 9940 34636 12124 34692
rect 12180 34636 13468 34692
rect 13524 34636 13534 34692
rect 22418 34636 22428 34692
rect 22484 34636 23772 34692
rect 23828 34636 23838 34692
rect 35186 34636 35196 34692
rect 35252 34636 37884 34692
rect 37940 34636 37950 34692
rect 40786 34636 40796 34692
rect 40852 34636 41692 34692
rect 41748 34636 42252 34692
rect 42308 34636 42318 34692
rect 42802 34636 42812 34692
rect 42868 34636 45052 34692
rect 45108 34636 45118 34692
rect 49298 34636 49308 34692
rect 49364 34636 50876 34692
rect 50932 34636 50942 34692
rect 51314 34636 51324 34692
rect 51380 34636 53228 34692
rect 53284 34636 53294 34692
rect 42252 34580 42308 34636
rect 4946 34524 4956 34580
rect 5012 34524 5740 34580
rect 5796 34524 5806 34580
rect 8978 34524 8988 34580
rect 9044 34524 10108 34580
rect 10164 34524 10174 34580
rect 23202 34524 23212 34580
rect 23268 34524 25900 34580
rect 25956 34524 25966 34580
rect 28578 34524 28588 34580
rect 28644 34524 29260 34580
rect 29316 34524 29326 34580
rect 32498 34524 32508 34580
rect 32564 34524 32732 34580
rect 32788 34524 33404 34580
rect 33460 34524 34412 34580
rect 34468 34524 34478 34580
rect 42252 34524 43260 34580
rect 43316 34524 43326 34580
rect 49634 34524 49644 34580
rect 49700 34524 50764 34580
rect 50820 34524 50830 34580
rect 9426 34412 9436 34468
rect 9492 34412 10332 34468
rect 10388 34412 10398 34468
rect 11890 34412 11900 34468
rect 11956 34412 12908 34468
rect 12964 34412 12974 34468
rect 0 34356 800 34384
rect 0 34300 12572 34356
rect 12628 34300 12638 34356
rect 0 34272 800 34300
rect 19826 34244 19836 34300
rect 19892 34244 19940 34300
rect 19996 34244 20044 34300
rect 20100 34244 20110 34300
rect 10882 34076 10892 34132
rect 10948 34076 12124 34132
rect 12180 34076 13020 34132
rect 13076 34076 13086 34132
rect 15026 33964 15036 34020
rect 15092 33964 16156 34020
rect 16212 33964 16222 34020
rect 13570 33852 13580 33908
rect 13636 33852 18452 33908
rect 18396 33796 18452 33852
rect 25900 33796 25956 34524
rect 28018 34412 28028 34468
rect 28084 34412 29484 34468
rect 29540 34412 29550 34468
rect 49074 34412 49084 34468
rect 49140 34412 50876 34468
rect 50932 34412 50942 34468
rect 50546 34244 50556 34300
rect 50612 34244 50660 34300
rect 50716 34244 50764 34300
rect 50820 34244 50830 34300
rect 40338 34188 40348 34244
rect 40404 34188 40414 34244
rect 40562 34188 40572 34244
rect 40628 34188 41468 34244
rect 41524 34188 41534 34244
rect 40348 34132 40404 34188
rect 38770 34076 38780 34132
rect 38836 34076 41804 34132
rect 41860 34076 41870 34132
rect 26786 33964 26796 34020
rect 26852 33964 27580 34020
rect 27636 33964 27646 34020
rect 35186 33964 35196 34020
rect 35252 33964 35868 34020
rect 35924 33964 36988 34020
rect 37044 33964 37054 34020
rect 39218 33964 39228 34020
rect 39284 33964 40348 34020
rect 40404 33964 41020 34020
rect 41076 33964 41086 34020
rect 54338 33964 54348 34020
rect 54404 33964 55804 34020
rect 55860 33964 55870 34020
rect 26450 33852 26460 33908
rect 26516 33852 27132 33908
rect 27188 33852 27198 33908
rect 33170 33852 33180 33908
rect 33236 33852 34972 33908
rect 35028 33852 44828 33908
rect 44884 33852 46284 33908
rect 46340 33852 47068 33908
rect 47124 33852 47134 33908
rect 57138 33852 57148 33908
rect 57204 33852 57708 33908
rect 57764 33852 57774 33908
rect 14466 33740 14476 33796
rect 14532 33740 15932 33796
rect 15988 33740 15998 33796
rect 18386 33740 18396 33796
rect 18452 33740 18462 33796
rect 22428 33740 23212 33796
rect 23268 33740 23278 33796
rect 25900 33740 27692 33796
rect 27748 33740 28700 33796
rect 28756 33740 28766 33796
rect 32050 33740 32060 33796
rect 32116 33740 32396 33796
rect 32452 33740 32732 33796
rect 32788 33740 32798 33796
rect 33506 33740 33516 33796
rect 33572 33740 34860 33796
rect 34916 33740 34926 33796
rect 35634 33740 35644 33796
rect 35700 33740 43820 33796
rect 43876 33740 43886 33796
rect 55570 33740 55580 33796
rect 55636 33740 56700 33796
rect 56756 33740 56766 33796
rect 22428 33684 22484 33740
rect 4274 33628 4284 33684
rect 4340 33628 5852 33684
rect 5908 33628 5918 33684
rect 12898 33628 12908 33684
rect 12964 33628 14364 33684
rect 14420 33628 14430 33684
rect 20514 33628 20524 33684
rect 20580 33628 21532 33684
rect 21588 33628 21980 33684
rect 22036 33628 22428 33684
rect 22484 33628 22494 33684
rect 22754 33628 22764 33684
rect 22820 33628 24668 33684
rect 24724 33628 25228 33684
rect 25284 33628 25294 33684
rect 29026 33628 29036 33684
rect 29092 33628 30716 33684
rect 30772 33628 30782 33684
rect 34066 33628 34076 33684
rect 34132 33628 35532 33684
rect 35588 33628 35598 33684
rect 38658 33628 38668 33684
rect 38724 33628 41244 33684
rect 41300 33628 42700 33684
rect 42756 33628 43148 33684
rect 43204 33628 43214 33684
rect 47170 33628 47180 33684
rect 47236 33628 48188 33684
rect 48244 33628 49420 33684
rect 49476 33628 49486 33684
rect 55682 33628 55692 33684
rect 55748 33628 57372 33684
rect 57428 33628 57438 33684
rect 10994 33516 11004 33572
rect 11060 33516 12460 33572
rect 12516 33516 12526 33572
rect 32162 33516 32172 33572
rect 32228 33516 39340 33572
rect 39396 33516 39406 33572
rect 50306 33516 50316 33572
rect 50372 33516 53900 33572
rect 53956 33516 53966 33572
rect 32498 33404 32508 33460
rect 32564 33404 33292 33460
rect 33348 33404 33358 33460
rect 34178 33404 34188 33460
rect 34244 33404 34748 33460
rect 34804 33404 35756 33460
rect 35812 33404 35822 33460
rect 37986 33404 37996 33460
rect 38052 33404 39116 33460
rect 39172 33404 39182 33460
rect 25750 33292 25788 33348
rect 25844 33292 25854 33348
rect 4466 33236 4476 33292
rect 4532 33236 4580 33292
rect 4636 33236 4684 33292
rect 4740 33236 4750 33292
rect 35186 33236 35196 33292
rect 35252 33236 35300 33292
rect 35356 33236 35404 33292
rect 35460 33236 35470 33292
rect 2706 33068 2716 33124
rect 2772 33068 3276 33124
rect 3332 33068 4844 33124
rect 4900 33068 4910 33124
rect 27906 33068 27916 33124
rect 27972 33068 28364 33124
rect 28420 33068 45164 33124
rect 45220 33068 45230 33124
rect 0 33012 800 33040
rect 0 32956 14700 33012
rect 14756 32956 14766 33012
rect 19282 32956 19292 33012
rect 19348 32956 20412 33012
rect 20468 32956 21084 33012
rect 21140 32956 21150 33012
rect 37314 32956 37324 33012
rect 37380 32956 38108 33012
rect 38164 32956 39228 33012
rect 39284 32956 39294 33012
rect 44930 32956 44940 33012
rect 44996 32956 46060 33012
rect 46116 32956 46126 33012
rect 0 32928 800 32956
rect 15698 32844 15708 32900
rect 15764 32844 18956 32900
rect 19012 32844 26124 32900
rect 26180 32844 26190 32900
rect 29922 32844 29932 32900
rect 29988 32844 31612 32900
rect 31668 32844 31948 32900
rect 32004 32844 32014 32900
rect 39106 32844 39116 32900
rect 39172 32844 41916 32900
rect 41972 32844 41982 32900
rect 56354 32844 56364 32900
rect 56420 32844 56924 32900
rect 56980 32844 57708 32900
rect 57764 32844 57774 32900
rect 3378 32732 3388 32788
rect 3444 32732 4396 32788
rect 4452 32732 4462 32788
rect 14578 32732 14588 32788
rect 14644 32732 15372 32788
rect 15428 32732 15438 32788
rect 18386 32732 18396 32788
rect 18452 32732 27020 32788
rect 27076 32732 27086 32788
rect 28578 32732 28588 32788
rect 28644 32732 48636 32788
rect 48692 32732 48702 32788
rect 53666 32732 53676 32788
rect 53732 32732 55132 32788
rect 55188 32732 55468 32788
rect 55412 32676 55468 32732
rect 39218 32620 39228 32676
rect 39284 32620 39676 32676
rect 39732 32620 40124 32676
rect 40180 32620 40190 32676
rect 55010 32620 55020 32676
rect 55076 32620 55086 32676
rect 55412 32620 56812 32676
rect 56868 32620 56878 32676
rect 55020 32564 55076 32620
rect 12786 32508 12796 32564
rect 12852 32508 17948 32564
rect 18004 32508 18014 32564
rect 41794 32508 41804 32564
rect 41860 32508 42812 32564
rect 42868 32508 43484 32564
rect 43540 32508 44156 32564
rect 44212 32508 45164 32564
rect 45220 32508 45230 32564
rect 55020 32508 56252 32564
rect 56308 32508 56318 32564
rect 10770 32396 10780 32452
rect 10836 32396 11788 32452
rect 11844 32396 11854 32452
rect 26852 32396 27692 32452
rect 27748 32396 27758 32452
rect 0 32340 800 32368
rect 26852 32340 26908 32396
rect 0 32284 16044 32340
rect 16100 32284 16110 32340
rect 23874 32284 23884 32340
rect 23940 32284 24780 32340
rect 24836 32284 26908 32340
rect 0 32256 800 32284
rect 19826 32228 19836 32284
rect 19892 32228 19940 32284
rect 19996 32228 20044 32284
rect 20100 32228 20110 32284
rect 50546 32228 50556 32284
rect 50612 32228 50660 32284
rect 50716 32228 50764 32284
rect 50820 32228 50830 32284
rect 27010 32172 27020 32228
rect 27076 32172 27580 32228
rect 27636 32172 27646 32228
rect 32610 32172 32620 32228
rect 32676 32172 33068 32228
rect 33124 32172 33134 32228
rect 31612 32060 31836 32116
rect 31892 32060 31902 32116
rect 24210 31948 24220 32004
rect 24276 31948 25340 32004
rect 25396 31948 25406 32004
rect 27346 31948 27356 32004
rect 27412 31948 28364 32004
rect 28420 31948 28430 32004
rect 31612 31892 31668 32060
rect 43250 31948 43260 32004
rect 43316 31948 44380 32004
rect 44436 31948 44446 32004
rect 55570 31948 55580 32004
rect 55636 31948 57036 32004
rect 57092 31948 57102 32004
rect 4946 31836 4956 31892
rect 5012 31836 5852 31892
rect 5908 31836 5918 31892
rect 11330 31836 11340 31892
rect 11396 31836 14364 31892
rect 14420 31836 14430 31892
rect 20178 31836 20188 31892
rect 20244 31836 20972 31892
rect 21028 31836 21038 31892
rect 21858 31836 21868 31892
rect 21924 31836 24108 31892
rect 24164 31836 24174 31892
rect 26422 31836 26460 31892
rect 26516 31836 26526 31892
rect 30930 31836 30940 31892
rect 30996 31836 31668 31892
rect 31826 31836 31836 31892
rect 31892 31836 35644 31892
rect 35700 31836 35710 31892
rect 37762 31836 37772 31892
rect 37828 31836 39900 31892
rect 39956 31836 39966 31892
rect 40226 31836 40236 31892
rect 40292 31836 41804 31892
rect 41860 31836 42812 31892
rect 42868 31836 42878 31892
rect 44034 31836 44044 31892
rect 44100 31836 47180 31892
rect 47236 31836 47246 31892
rect 47506 31836 47516 31892
rect 47572 31836 49420 31892
rect 49476 31836 50204 31892
rect 50260 31836 50270 31892
rect 52098 31836 52108 31892
rect 52164 31836 53676 31892
rect 53732 31836 55020 31892
rect 55076 31836 56028 31892
rect 56084 31836 56924 31892
rect 56980 31836 56990 31892
rect 39900 31780 39956 31836
rect 47180 31780 47236 31836
rect 13906 31724 13916 31780
rect 13972 31724 14476 31780
rect 14532 31724 15372 31780
rect 15428 31724 15438 31780
rect 16370 31724 16380 31780
rect 16436 31724 20860 31780
rect 20916 31724 20926 31780
rect 21410 31724 21420 31780
rect 21476 31724 23212 31780
rect 23268 31724 23278 31780
rect 25228 31724 26012 31780
rect 26068 31724 27468 31780
rect 27524 31724 27534 31780
rect 29810 31724 29820 31780
rect 29876 31724 33628 31780
rect 33684 31724 33694 31780
rect 34738 31724 34748 31780
rect 34804 31724 35532 31780
rect 35588 31724 35598 31780
rect 35746 31724 35756 31780
rect 35812 31724 36988 31780
rect 37044 31724 37054 31780
rect 39900 31724 44268 31780
rect 44324 31724 44334 31780
rect 45154 31724 45164 31780
rect 45220 31724 46396 31780
rect 46452 31724 46956 31780
rect 47012 31724 47022 31780
rect 47180 31724 47964 31780
rect 48020 31724 48030 31780
rect 52434 31724 52444 31780
rect 52500 31724 53452 31780
rect 53508 31724 53518 31780
rect 0 31668 800 31696
rect 25228 31668 25284 31724
rect 32732 31668 32788 31724
rect 43820 31668 43876 31724
rect 0 31612 14924 31668
rect 14980 31612 14990 31668
rect 22754 31612 22764 31668
rect 22820 31612 25228 31668
rect 25284 31612 25294 31668
rect 25778 31612 25788 31668
rect 25844 31612 27020 31668
rect 27076 31612 27086 31668
rect 32722 31612 32732 31668
rect 32788 31612 32798 31668
rect 40338 31612 40348 31668
rect 40404 31612 40908 31668
rect 40964 31612 40974 31668
rect 43810 31612 43820 31668
rect 43876 31612 43886 31668
rect 44930 31612 44940 31668
rect 44996 31612 45388 31668
rect 45444 31612 46732 31668
rect 46788 31612 46798 31668
rect 50194 31612 50204 31668
rect 50260 31612 51660 31668
rect 51716 31612 52780 31668
rect 52836 31612 52846 31668
rect 56690 31612 56700 31668
rect 56756 31612 57148 31668
rect 57204 31612 57214 31668
rect 0 31584 800 31612
rect 40908 31556 40964 31612
rect 17826 31500 17836 31556
rect 17892 31500 20748 31556
rect 20804 31500 21756 31556
rect 21812 31500 21822 31556
rect 22866 31500 22876 31556
rect 22932 31500 24108 31556
rect 24164 31500 24174 31556
rect 24994 31500 25004 31556
rect 25060 31500 26348 31556
rect 26404 31500 26414 31556
rect 40908 31500 48748 31556
rect 48804 31500 49532 31556
rect 49588 31500 49598 31556
rect 51538 31500 51548 31556
rect 51604 31500 53340 31556
rect 53396 31500 53406 31556
rect 20850 31388 20860 31444
rect 20916 31388 23772 31444
rect 23828 31388 23838 31444
rect 26898 31388 26908 31444
rect 26964 31388 27132 31444
rect 27188 31388 27198 31444
rect 36530 31388 36540 31444
rect 36596 31388 37660 31444
rect 37716 31388 38668 31444
rect 38612 31332 38668 31388
rect 13458 31276 13468 31332
rect 13524 31276 16828 31332
rect 16884 31276 20188 31332
rect 20244 31276 20254 31332
rect 38612 31276 40348 31332
rect 40404 31276 40414 31332
rect 4466 31220 4476 31276
rect 4532 31220 4580 31276
rect 4636 31220 4684 31276
rect 4740 31220 4750 31276
rect 35186 31220 35196 31276
rect 35252 31220 35300 31276
rect 35356 31220 35404 31276
rect 35460 31220 35470 31276
rect 15922 31052 15932 31108
rect 15988 31052 25116 31108
rect 25172 31052 25182 31108
rect 26674 31052 26684 31108
rect 26740 31052 27580 31108
rect 27636 31052 27646 31108
rect 40562 31052 40572 31108
rect 40628 31052 41132 31108
rect 41188 31052 41692 31108
rect 41748 31052 41758 31108
rect 0 30996 800 31024
rect 0 30940 15036 30996
rect 15092 30940 15102 30996
rect 0 30912 800 30940
rect 2370 30828 2380 30884
rect 2436 30828 2716 30884
rect 2772 30828 5628 30884
rect 5684 30828 5694 30884
rect 19170 30828 19180 30884
rect 19236 30828 25788 30884
rect 25844 30828 25854 30884
rect 26226 30828 26236 30884
rect 26292 30828 28252 30884
rect 28308 30828 28318 30884
rect 41906 30828 41916 30884
rect 41972 30828 44044 30884
rect 44100 30828 45276 30884
rect 45332 30828 46620 30884
rect 46676 30828 46686 30884
rect 23986 30716 23996 30772
rect 24052 30716 25900 30772
rect 25956 30716 25966 30772
rect 27906 30716 27916 30772
rect 27972 30716 29708 30772
rect 29764 30716 29774 30772
rect 29932 30716 34692 30772
rect 35746 30716 35756 30772
rect 35812 30716 37324 30772
rect 37380 30716 37390 30772
rect 39218 30716 39228 30772
rect 39284 30716 39900 30772
rect 39956 30716 41356 30772
rect 41412 30716 41422 30772
rect 43698 30716 43708 30772
rect 43764 30716 45948 30772
rect 46004 30716 46844 30772
rect 46900 30716 46910 30772
rect 49308 30716 50316 30772
rect 50372 30716 50382 30772
rect 29932 30660 29988 30716
rect 34636 30660 34692 30716
rect 49308 30660 49364 30716
rect 13906 30604 13916 30660
rect 13972 30604 15484 30660
rect 15540 30604 15550 30660
rect 24994 30604 25004 30660
rect 25060 30604 25564 30660
rect 25620 30604 25630 30660
rect 26338 30604 26348 30660
rect 26404 30604 26908 30660
rect 26964 30604 26974 30660
rect 29138 30604 29148 30660
rect 29204 30604 29988 30660
rect 30818 30604 30828 30660
rect 30884 30604 32060 30660
rect 32116 30604 34412 30660
rect 34468 30604 34478 30660
rect 34636 30604 38220 30660
rect 38276 30604 38286 30660
rect 48738 30604 48748 30660
rect 48804 30604 48972 30660
rect 49028 30604 49308 30660
rect 49364 30604 49374 30660
rect 53554 30604 53564 30660
rect 53620 30604 54236 30660
rect 54292 30604 54684 30660
rect 54740 30604 54750 30660
rect 4946 30492 4956 30548
rect 5012 30492 5740 30548
rect 5796 30492 5806 30548
rect 9314 30492 9324 30548
rect 9380 30492 10444 30548
rect 10500 30492 12460 30548
rect 12516 30492 13468 30548
rect 13524 30492 13534 30548
rect 14578 30492 14588 30548
rect 14644 30492 17724 30548
rect 17780 30492 17790 30548
rect 22642 30492 22652 30548
rect 22708 30492 26684 30548
rect 26740 30492 26750 30548
rect 32946 30492 32956 30548
rect 33012 30492 33628 30548
rect 33684 30492 33694 30548
rect 35522 30492 35532 30548
rect 35588 30492 38444 30548
rect 38500 30492 39676 30548
rect 39732 30492 40348 30548
rect 40404 30492 40414 30548
rect 48290 30492 48300 30548
rect 48356 30492 49980 30548
rect 50036 30492 50046 30548
rect 6738 30380 6748 30436
rect 6804 30380 13580 30436
rect 13636 30380 13646 30436
rect 16034 30380 16044 30436
rect 16100 30380 18284 30436
rect 18340 30380 26460 30436
rect 26516 30380 26526 30436
rect 28578 30380 28588 30436
rect 28644 30380 29260 30436
rect 29316 30380 48636 30436
rect 48692 30380 48702 30436
rect 51314 30380 51324 30436
rect 51380 30380 52556 30436
rect 52612 30380 52622 30436
rect 0 30324 800 30352
rect 0 30268 4228 30324
rect 4722 30268 4732 30324
rect 4788 30268 6076 30324
rect 6132 30268 6142 30324
rect 26002 30268 26012 30324
rect 26068 30268 26796 30324
rect 26852 30268 26862 30324
rect 27346 30268 27356 30324
rect 27412 30268 29036 30324
rect 29092 30268 29102 30324
rect 35970 30268 35980 30324
rect 36036 30268 36652 30324
rect 36708 30268 37996 30324
rect 38052 30268 38062 30324
rect 38210 30268 38220 30324
rect 38276 30268 40124 30324
rect 40180 30268 40190 30324
rect 50978 30268 50988 30324
rect 51044 30268 52444 30324
rect 52500 30268 53004 30324
rect 53060 30268 54236 30324
rect 54292 30268 56700 30324
rect 56756 30268 56766 30324
rect 0 30240 800 30268
rect 4172 30212 4228 30268
rect 19826 30212 19836 30268
rect 19892 30212 19940 30268
rect 19996 30212 20044 30268
rect 20100 30212 20110 30268
rect 50546 30212 50556 30268
rect 50612 30212 50660 30268
rect 50716 30212 50764 30268
rect 50820 30212 50830 30268
rect 4172 30156 14252 30212
rect 14308 30156 14318 30212
rect 25778 30156 25788 30212
rect 25844 30156 29596 30212
rect 29652 30156 29662 30212
rect 31378 30156 31388 30212
rect 31444 30156 31454 30212
rect 34850 30156 34860 30212
rect 34916 30156 36540 30212
rect 36596 30156 43932 30212
rect 43988 30156 43998 30212
rect 1810 30044 1820 30100
rect 1876 30044 3836 30100
rect 3892 30044 3902 30100
rect 9650 30044 9660 30100
rect 9716 30044 10332 30100
rect 10388 30044 10398 30100
rect 17714 30044 17724 30100
rect 17780 30044 25564 30100
rect 25620 30044 25630 30100
rect 27010 30044 27020 30100
rect 27076 30044 28140 30100
rect 28196 30044 28206 30100
rect 31388 29988 31444 30156
rect 32610 30044 32620 30100
rect 32676 30044 35532 30100
rect 35588 30044 35598 30100
rect 39442 30044 39452 30100
rect 39508 30044 43484 30100
rect 43540 30044 46060 30100
rect 46116 30044 46126 30100
rect 8530 29932 8540 29988
rect 8596 29932 9324 29988
rect 9380 29932 9390 29988
rect 23090 29932 23100 29988
rect 23156 29932 24332 29988
rect 24388 29932 24398 29988
rect 24546 29932 24556 29988
rect 24612 29932 25788 29988
rect 25844 29932 25854 29988
rect 31388 29932 43372 29988
rect 43428 29932 43438 29988
rect 6178 29820 6188 29876
rect 6244 29820 6972 29876
rect 7028 29820 7308 29876
rect 7364 29820 7374 29876
rect 15250 29820 15260 29876
rect 15316 29820 19180 29876
rect 19236 29820 19246 29876
rect 19618 29820 19628 29876
rect 19684 29820 24444 29876
rect 24500 29820 24510 29876
rect 25554 29820 25564 29876
rect 25620 29820 27132 29876
rect 27188 29820 27198 29876
rect 33506 29820 33516 29876
rect 33572 29820 34188 29876
rect 34244 29820 36204 29876
rect 36260 29820 36988 29876
rect 37044 29820 37054 29876
rect 49634 29820 49644 29876
rect 49700 29820 50876 29876
rect 50932 29820 50942 29876
rect 52770 29820 52780 29876
rect 52836 29820 54348 29876
rect 54404 29820 54414 29876
rect 1922 29708 1932 29764
rect 1988 29708 3724 29764
rect 3780 29708 3790 29764
rect 9986 29708 9996 29764
rect 10052 29708 12908 29764
rect 12964 29708 12974 29764
rect 24322 29708 24332 29764
rect 24388 29708 25004 29764
rect 25060 29708 25676 29764
rect 25732 29708 26572 29764
rect 26628 29708 26638 29764
rect 27682 29708 27692 29764
rect 27748 29708 29260 29764
rect 29316 29708 29326 29764
rect 29922 29708 29932 29764
rect 29988 29708 33180 29764
rect 33236 29708 33246 29764
rect 33730 29708 33740 29764
rect 33796 29708 35420 29764
rect 35476 29708 35486 29764
rect 44482 29708 44492 29764
rect 44548 29708 46172 29764
rect 46228 29708 46238 29764
rect 49858 29708 49868 29764
rect 49924 29708 53452 29764
rect 53508 29708 53518 29764
rect 0 29652 800 29680
rect 0 29596 13916 29652
rect 13972 29596 13982 29652
rect 27458 29596 27468 29652
rect 27524 29596 28476 29652
rect 28532 29596 28924 29652
rect 28980 29596 31612 29652
rect 31668 29596 31678 29652
rect 31826 29596 31836 29652
rect 31892 29596 32172 29652
rect 32228 29596 32238 29652
rect 34514 29596 34524 29652
rect 34580 29596 37100 29652
rect 37156 29596 48188 29652
rect 48244 29596 49308 29652
rect 49364 29596 49374 29652
rect 0 29568 800 29596
rect 3378 29484 3388 29540
rect 3444 29484 8764 29540
rect 8820 29484 8830 29540
rect 23874 29484 23884 29540
rect 23940 29484 25228 29540
rect 25284 29484 27020 29540
rect 27076 29484 27086 29540
rect 31266 29484 31276 29540
rect 31332 29484 34860 29540
rect 34916 29484 35196 29540
rect 35252 29484 37212 29540
rect 37268 29484 37548 29540
rect 37604 29484 37614 29540
rect 3266 29372 3276 29428
rect 3332 29372 5068 29428
rect 5124 29372 5134 29428
rect 7858 29372 7868 29428
rect 7924 29372 8876 29428
rect 8932 29372 10108 29428
rect 10164 29372 10174 29428
rect 29026 29372 29036 29428
rect 29092 29372 40796 29428
rect 40852 29372 40862 29428
rect 32162 29260 32172 29316
rect 32228 29260 34636 29316
rect 34692 29260 34702 29316
rect 4466 29204 4476 29260
rect 4532 29204 4580 29260
rect 4636 29204 4684 29260
rect 4740 29204 4750 29260
rect 35186 29204 35196 29260
rect 35252 29204 35300 29260
rect 35356 29204 35404 29260
rect 35460 29204 35470 29260
rect 24210 29148 24220 29204
rect 24276 29148 29820 29204
rect 29876 29148 29886 29204
rect 4274 29036 4284 29092
rect 4340 29036 5516 29092
rect 5572 29036 5582 29092
rect 9650 29036 9660 29092
rect 9716 29036 11340 29092
rect 11396 29036 13468 29092
rect 13524 29036 13534 29092
rect 30034 29036 30044 29092
rect 30100 29036 31276 29092
rect 31332 29036 31342 29092
rect 31714 29036 31724 29092
rect 31780 29036 34580 29092
rect 0 28980 800 29008
rect 34524 28980 34580 29036
rect 0 28924 3668 28980
rect 3826 28924 3836 28980
rect 3892 28924 4508 28980
rect 4564 28924 4574 28980
rect 6738 28924 6748 28980
rect 6804 28924 6814 28980
rect 10434 28924 10444 28980
rect 10500 28924 12796 28980
rect 12852 28924 14028 28980
rect 14084 28924 14094 28980
rect 24210 28924 24220 28980
rect 24276 28924 25004 28980
rect 25060 28924 25070 28980
rect 26898 28924 26908 28980
rect 26964 28924 30716 28980
rect 30772 28924 30782 28980
rect 33282 28924 33292 28980
rect 33348 28924 33516 28980
rect 33572 28924 33582 28980
rect 34514 28924 34524 28980
rect 34580 28924 36092 28980
rect 36148 28924 46508 28980
rect 46564 28924 46574 28980
rect 0 28896 800 28924
rect 3612 28868 3668 28924
rect 6748 28868 6804 28924
rect 3612 28812 6804 28868
rect 15092 28812 19628 28868
rect 19684 28812 19694 28868
rect 26338 28812 26348 28868
rect 26404 28812 27580 28868
rect 27636 28812 27646 28868
rect 29474 28812 29484 28868
rect 29540 28812 30380 28868
rect 30436 28812 30446 28868
rect 31490 28812 31500 28868
rect 31556 28812 32620 28868
rect 32676 28812 32686 28868
rect 39890 28812 39900 28868
rect 39956 28812 41244 28868
rect 41300 28812 41310 28868
rect 49746 28812 49756 28868
rect 49812 28812 52780 28868
rect 52836 28812 52846 28868
rect 54002 28812 54012 28868
rect 54068 28812 54796 28868
rect 54852 28812 54862 28868
rect 5058 28700 5068 28756
rect 5124 28700 6188 28756
rect 6244 28700 6254 28756
rect 12898 28700 12908 28756
rect 12964 28700 14476 28756
rect 14532 28700 14542 28756
rect 8978 28588 8988 28644
rect 9044 28588 12796 28644
rect 12852 28588 14700 28644
rect 14756 28588 14766 28644
rect 15026 28588 15036 28644
rect 15092 28588 15148 28812
rect 19506 28700 19516 28756
rect 19572 28700 20300 28756
rect 20356 28700 21308 28756
rect 21364 28700 22316 28756
rect 22372 28700 22988 28756
rect 23044 28700 23054 28756
rect 25106 28700 25116 28756
rect 25172 28700 29148 28756
rect 29204 28700 29214 28756
rect 30146 28700 30156 28756
rect 30212 28700 32956 28756
rect 33012 28700 33022 28756
rect 45602 28700 45612 28756
rect 45668 28700 45948 28756
rect 46004 28700 48188 28756
rect 48244 28700 50316 28756
rect 50372 28700 50540 28756
rect 50596 28700 50606 28756
rect 17826 28588 17836 28644
rect 17892 28588 20748 28644
rect 20804 28588 21756 28644
rect 21812 28588 21822 28644
rect 31042 28588 31052 28644
rect 31108 28588 34076 28644
rect 34132 28588 34142 28644
rect 38322 28588 38332 28644
rect 38388 28588 38556 28644
rect 38612 28588 39116 28644
rect 39172 28588 39182 28644
rect 48636 28588 48748 28644
rect 48804 28588 49084 28644
rect 49140 28588 50988 28644
rect 51044 28588 51054 28644
rect 52770 28588 52780 28644
rect 52836 28588 55132 28644
rect 55188 28588 55198 28644
rect 48636 28532 48692 28588
rect 8418 28476 8428 28532
rect 8484 28476 9100 28532
rect 9156 28476 9166 28532
rect 24994 28476 25004 28532
rect 25060 28476 25900 28532
rect 25956 28476 26572 28532
rect 26628 28476 26638 28532
rect 32610 28476 32620 28532
rect 32676 28476 38780 28532
rect 38836 28476 45164 28532
rect 45220 28476 45230 28532
rect 47058 28476 47068 28532
rect 47124 28476 47740 28532
rect 47796 28476 48692 28532
rect 55794 28476 55804 28532
rect 55860 28476 56924 28532
rect 56980 28476 56990 28532
rect 26114 28364 26124 28420
rect 26180 28364 26460 28420
rect 26516 28364 27020 28420
rect 27076 28364 31836 28420
rect 31892 28364 31902 28420
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 33506 28140 33516 28196
rect 33572 28140 35196 28196
rect 35252 28140 35262 28196
rect 34626 28028 34636 28084
rect 34692 28028 35532 28084
rect 35588 28028 35598 28084
rect 24882 27916 24892 27972
rect 24948 27916 25228 27972
rect 25284 27916 25294 27972
rect 29810 27916 29820 27972
rect 29876 27916 30828 27972
rect 30884 27916 30894 27972
rect 51314 27916 51324 27972
rect 51380 27916 53116 27972
rect 53172 27916 53182 27972
rect 1810 27804 1820 27860
rect 1876 27804 2380 27860
rect 2436 27804 2940 27860
rect 2996 27804 3388 27860
rect 3444 27804 4284 27860
rect 4340 27804 5068 27860
rect 5124 27804 5740 27860
rect 5796 27804 5806 27860
rect 32610 27804 32620 27860
rect 32676 27804 33516 27860
rect 33572 27804 33582 27860
rect 33842 27804 33852 27860
rect 33908 27804 34524 27860
rect 34580 27804 34590 27860
rect 45266 27804 45276 27860
rect 45332 27804 46620 27860
rect 46676 27804 46686 27860
rect 54898 27804 54908 27860
rect 54964 27804 56924 27860
rect 56980 27804 56990 27860
rect 20850 27692 20860 27748
rect 20916 27692 22204 27748
rect 22260 27692 22270 27748
rect 23650 27692 23660 27748
rect 23716 27692 24444 27748
rect 24500 27692 24510 27748
rect 24658 27692 24668 27748
rect 24724 27692 26348 27748
rect 26404 27692 26908 27748
rect 32162 27692 32172 27748
rect 32228 27692 34188 27748
rect 34244 27692 34254 27748
rect 35074 27692 35084 27748
rect 35140 27692 35644 27748
rect 35700 27692 35710 27748
rect 51986 27692 51996 27748
rect 52052 27692 52780 27748
rect 52836 27692 52846 27748
rect 55682 27692 55692 27748
rect 55748 27692 56588 27748
rect 56644 27692 58156 27748
rect 58212 27692 58222 27748
rect 26852 27636 26908 27692
rect 26852 27580 29708 27636
rect 29764 27580 31500 27636
rect 31556 27580 31566 27636
rect 46050 27580 46060 27636
rect 46116 27580 47740 27636
rect 47796 27580 47806 27636
rect 49074 27580 49084 27636
rect 49140 27580 52444 27636
rect 52500 27580 53116 27636
rect 53172 27580 53182 27636
rect 33170 27468 33180 27524
rect 33236 27468 35084 27524
rect 35140 27468 35150 27524
rect 46946 27468 46956 27524
rect 47012 27468 48412 27524
rect 48468 27468 51324 27524
rect 51380 27468 51390 27524
rect 21634 27356 21644 27412
rect 21700 27356 22876 27412
rect 22932 27356 22942 27412
rect 46722 27356 46732 27412
rect 46788 27356 49084 27412
rect 49140 27356 49150 27412
rect 4466 27188 4476 27244
rect 4532 27188 4580 27244
rect 4636 27188 4684 27244
rect 4740 27188 4750 27244
rect 35186 27188 35196 27244
rect 35252 27188 35300 27244
rect 35356 27188 35404 27244
rect 35460 27188 35470 27244
rect 33590 27132 33628 27188
rect 33684 27132 33694 27188
rect 25218 27020 25228 27076
rect 25284 27020 26348 27076
rect 26404 27020 26414 27076
rect 39330 27020 39340 27076
rect 39396 27020 41020 27076
rect 41076 27020 41086 27076
rect 26002 26908 26012 26964
rect 26068 26908 29596 26964
rect 29652 26908 29662 26964
rect 40338 26908 40348 26964
rect 40404 26908 42140 26964
rect 42196 26908 42206 26964
rect 50418 26908 50428 26964
rect 50484 26908 53564 26964
rect 53620 26908 53630 26964
rect 53778 26908 53788 26964
rect 53844 26908 57260 26964
rect 57316 26908 57326 26964
rect 22530 26796 22540 26852
rect 22596 26796 24556 26852
rect 24612 26796 24622 26852
rect 31602 26796 31612 26852
rect 31668 26796 32284 26852
rect 32340 26796 32350 26852
rect 35522 26796 35532 26852
rect 35588 26796 39452 26852
rect 39508 26796 39518 26852
rect 52658 26796 52668 26852
rect 52724 26796 55468 26852
rect 55412 26740 55468 26796
rect 15922 26684 15932 26740
rect 15988 26684 24668 26740
rect 24724 26684 24734 26740
rect 24994 26684 25004 26740
rect 25060 26684 25676 26740
rect 25732 26684 25742 26740
rect 30594 26684 30604 26740
rect 30660 26684 31948 26740
rect 32004 26684 32014 26740
rect 32498 26684 32508 26740
rect 32564 26684 32574 26740
rect 33282 26684 33292 26740
rect 33348 26684 33358 26740
rect 35858 26684 35868 26740
rect 35924 26684 38220 26740
rect 38276 26684 38286 26740
rect 51426 26684 51436 26740
rect 51492 26684 53564 26740
rect 53620 26684 54012 26740
rect 54068 26684 54078 26740
rect 55412 26684 55804 26740
rect 55860 26684 55870 26740
rect 32508 26628 32564 26684
rect 17042 26572 17052 26628
rect 17108 26572 17948 26628
rect 18004 26572 21868 26628
rect 21924 26572 21934 26628
rect 23538 26572 23548 26628
rect 23604 26572 24556 26628
rect 24612 26572 24622 26628
rect 31714 26572 31724 26628
rect 31780 26572 32564 26628
rect 31724 26516 31780 26572
rect 20738 26460 20748 26516
rect 20804 26460 22092 26516
rect 22148 26460 22158 26516
rect 23314 26460 23324 26516
rect 23380 26460 23772 26516
rect 23828 26460 24612 26516
rect 25554 26460 25564 26516
rect 25620 26460 27356 26516
rect 27412 26460 27422 26516
rect 31378 26460 31388 26516
rect 31444 26460 31780 26516
rect 32050 26460 32060 26516
rect 32116 26460 32956 26516
rect 33012 26460 33022 26516
rect 24556 26404 24612 26460
rect 33292 26404 33348 26684
rect 34178 26572 34188 26628
rect 34244 26572 36540 26628
rect 36596 26572 36606 26628
rect 37650 26572 37660 26628
rect 37716 26572 38780 26628
rect 38836 26572 38846 26628
rect 33842 26460 33852 26516
rect 33908 26460 35196 26516
rect 35252 26460 35868 26516
rect 35924 26460 35934 26516
rect 42018 26460 42028 26516
rect 42084 26460 44828 26516
rect 44884 26460 45500 26516
rect 45556 26460 45566 26516
rect 49298 26460 49308 26516
rect 49364 26460 50204 26516
rect 50260 26460 50540 26516
rect 50596 26460 51100 26516
rect 51156 26460 51166 26516
rect 52770 26460 52780 26516
rect 52836 26460 53676 26516
rect 53732 26460 53742 26516
rect 18946 26348 18956 26404
rect 19012 26348 19852 26404
rect 19908 26348 20972 26404
rect 21028 26348 21038 26404
rect 23202 26348 23212 26404
rect 23268 26348 24332 26404
rect 24388 26348 24398 26404
rect 24556 26348 33348 26404
rect 43922 26348 43932 26404
rect 43988 26348 48524 26404
rect 48580 26348 48590 26404
rect 22530 26236 22540 26292
rect 22596 26236 24220 26292
rect 24276 26236 29484 26292
rect 29540 26236 30604 26292
rect 30660 26236 31724 26292
rect 31780 26236 31790 26292
rect 32498 26236 32508 26292
rect 32564 26236 33516 26292
rect 33572 26236 33582 26292
rect 37986 26236 37996 26292
rect 38052 26236 38668 26292
rect 38724 26236 38734 26292
rect 19826 26180 19836 26236
rect 19892 26180 19940 26236
rect 19996 26180 20044 26236
rect 20100 26180 20110 26236
rect 50546 26180 50556 26236
rect 50612 26180 50660 26236
rect 50716 26180 50764 26236
rect 50820 26180 50830 26236
rect 30146 26124 30156 26180
rect 30212 26124 45836 26180
rect 45892 26124 45902 26180
rect 17714 26012 17724 26068
rect 17780 26012 21420 26068
rect 21476 26012 21486 26068
rect 21858 26012 21868 26068
rect 21924 26012 22764 26068
rect 22820 26012 22830 26068
rect 24434 26012 24444 26068
rect 24500 26012 25116 26068
rect 25172 26012 25182 26068
rect 26898 26012 26908 26068
rect 26964 26012 29932 26068
rect 29988 26012 29998 26068
rect 16706 25900 16716 25956
rect 16772 25900 18172 25956
rect 18228 25900 18238 25956
rect 26114 25900 26124 25956
rect 26180 25900 26572 25956
rect 26628 25900 26908 25956
rect 27906 25900 27916 25956
rect 27972 25900 28588 25956
rect 28644 25900 29372 25956
rect 29428 25900 31388 25956
rect 31444 25900 31454 25956
rect 34402 25900 34412 25956
rect 34468 25900 35532 25956
rect 35588 25900 35598 25956
rect 38612 25900 42252 25956
rect 42308 25900 42318 25956
rect 46162 25900 46172 25956
rect 46228 25900 49308 25956
rect 49364 25900 50764 25956
rect 50820 25900 50830 25956
rect 54450 25900 54460 25956
rect 54516 25900 55356 25956
rect 55412 25900 55422 25956
rect 26852 25844 26908 25900
rect 38612 25844 38668 25900
rect 14578 25788 14588 25844
rect 14644 25788 17612 25844
rect 17668 25788 17678 25844
rect 23426 25788 23436 25844
rect 23492 25788 26684 25844
rect 26740 25788 26750 25844
rect 26852 25788 27020 25844
rect 27076 25788 27086 25844
rect 30818 25788 30828 25844
rect 30884 25788 38668 25844
rect 54002 25788 54012 25844
rect 54068 25788 54572 25844
rect 54628 25788 55468 25844
rect 21410 25676 21420 25732
rect 21476 25676 22428 25732
rect 22484 25676 22494 25732
rect 24882 25676 24892 25732
rect 24948 25676 25900 25732
rect 25956 25676 25966 25732
rect 31714 25676 31724 25732
rect 31780 25676 32172 25732
rect 32228 25676 32238 25732
rect 32610 25676 32620 25732
rect 32676 25676 33852 25732
rect 33908 25676 33918 25732
rect 36418 25676 36428 25732
rect 36484 25676 36876 25732
rect 36932 25676 37548 25732
rect 37604 25676 37996 25732
rect 38052 25676 38062 25732
rect 38658 25676 38668 25732
rect 38724 25676 39676 25732
rect 39732 25676 40348 25732
rect 40404 25676 41244 25732
rect 41300 25676 41310 25732
rect 46274 25676 46284 25732
rect 46340 25676 50876 25732
rect 50932 25676 50942 25732
rect 55412 25620 55468 25788
rect 24546 25564 24556 25620
rect 24612 25564 25564 25620
rect 25620 25564 26572 25620
rect 26628 25564 26638 25620
rect 27682 25564 27692 25620
rect 27748 25564 28028 25620
rect 28084 25564 28588 25620
rect 28644 25564 29596 25620
rect 29652 25564 31164 25620
rect 31220 25564 32844 25620
rect 32900 25564 32910 25620
rect 33394 25564 33404 25620
rect 33460 25564 34972 25620
rect 35028 25564 35038 25620
rect 35634 25564 35644 25620
rect 35700 25564 37436 25620
rect 37492 25564 37772 25620
rect 37828 25564 37838 25620
rect 45938 25564 45948 25620
rect 46004 25564 46508 25620
rect 46564 25564 46574 25620
rect 55412 25564 55580 25620
rect 55636 25564 56028 25620
rect 56084 25564 56700 25620
rect 56756 25564 56766 25620
rect 25330 25452 25340 25508
rect 25396 25452 30156 25508
rect 30212 25452 30222 25508
rect 32050 25452 32060 25508
rect 32116 25452 35868 25508
rect 35924 25452 35934 25508
rect 36082 25452 36092 25508
rect 36148 25452 37548 25508
rect 37604 25452 37614 25508
rect 18610 25340 18620 25396
rect 18676 25340 20188 25396
rect 25218 25340 25228 25396
rect 25284 25340 26348 25396
rect 26404 25340 26908 25396
rect 26964 25340 27244 25396
rect 27300 25340 27310 25396
rect 34962 25340 34972 25396
rect 35028 25340 36204 25396
rect 36260 25340 36270 25396
rect 20132 25284 20188 25340
rect 20132 25228 25788 25284
rect 25844 25228 25854 25284
rect 4466 25172 4476 25228
rect 4532 25172 4580 25228
rect 4636 25172 4684 25228
rect 4740 25172 4750 25228
rect 35186 25172 35196 25228
rect 35252 25172 35300 25228
rect 35356 25172 35404 25228
rect 35460 25172 35470 25228
rect 26786 25004 26796 25060
rect 26852 25004 30716 25060
rect 30772 25004 30782 25060
rect 30034 24892 30044 24948
rect 30100 24892 30828 24948
rect 30884 24892 30894 24948
rect 19394 24780 19404 24836
rect 19460 24780 21644 24836
rect 21700 24780 21710 24836
rect 21980 24780 22092 24836
rect 22148 24780 24724 24836
rect 36642 24780 36652 24836
rect 36708 24780 37884 24836
rect 37940 24780 37950 24836
rect 48402 24780 48412 24836
rect 48468 24780 50988 24836
rect 51044 24780 51548 24836
rect 51604 24780 51614 24836
rect 20132 24556 20188 24780
rect 21980 24724 22036 24780
rect 24668 24724 24724 24780
rect 21074 24668 21084 24724
rect 21140 24668 22036 24724
rect 22194 24668 22204 24724
rect 22260 24668 23324 24724
rect 23380 24668 23390 24724
rect 24658 24668 24668 24724
rect 24724 24668 25452 24724
rect 25508 24668 25620 24724
rect 26114 24668 26124 24724
rect 26180 24668 26460 24724
rect 26516 24668 26526 24724
rect 38882 24668 38892 24724
rect 38948 24668 39788 24724
rect 39844 24668 39854 24724
rect 25564 24612 25620 24668
rect 20244 24556 20254 24612
rect 22306 24556 22316 24612
rect 22372 24556 23884 24612
rect 23940 24556 23950 24612
rect 24546 24556 24556 24612
rect 24612 24556 25340 24612
rect 25396 24556 25406 24612
rect 25564 24556 27468 24612
rect 27524 24556 28924 24612
rect 28980 24556 29260 24612
rect 29316 24556 29326 24612
rect 30258 24556 30268 24612
rect 30324 24556 31948 24612
rect 32004 24556 34748 24612
rect 34804 24556 34814 24612
rect 55346 24556 55356 24612
rect 55412 24556 56812 24612
rect 56868 24556 56878 24612
rect 23884 24500 23940 24556
rect 21746 24444 21756 24500
rect 21812 24444 22876 24500
rect 22932 24444 22942 24500
rect 23884 24444 25676 24500
rect 25732 24444 26460 24500
rect 26516 24444 27580 24500
rect 27636 24444 27646 24500
rect 29586 24444 29596 24500
rect 29652 24444 30604 24500
rect 30660 24444 31500 24500
rect 31556 24444 31566 24500
rect 35522 24444 35532 24500
rect 35588 24444 35980 24500
rect 36036 24444 36876 24500
rect 36932 24444 36942 24500
rect 51202 24444 51212 24500
rect 51268 24444 54124 24500
rect 54180 24444 54190 24500
rect 20290 24332 20300 24388
rect 20356 24332 22652 24388
rect 22708 24332 23548 24388
rect 23604 24332 27692 24388
rect 27748 24332 27758 24388
rect 29810 24332 29820 24388
rect 29876 24332 33628 24388
rect 33684 24332 33694 24388
rect 40562 24332 40572 24388
rect 40628 24332 41468 24388
rect 41524 24332 41534 24388
rect 48178 24332 48188 24388
rect 48244 24332 49644 24388
rect 49700 24332 49710 24388
rect 19826 24164 19836 24220
rect 19892 24164 19940 24220
rect 19996 24164 20044 24220
rect 20100 24164 20110 24220
rect 50546 24164 50556 24220
rect 50612 24164 50660 24220
rect 50716 24164 50764 24220
rect 50820 24164 50830 24220
rect 25778 23996 25788 24052
rect 25844 23996 26348 24052
rect 26404 23996 26414 24052
rect 29362 23996 29372 24052
rect 29428 23996 30604 24052
rect 30660 23996 30670 24052
rect 45266 23996 45276 24052
rect 45332 23996 47740 24052
rect 47796 23996 48748 24052
rect 48804 23996 49980 24052
rect 50036 23996 50046 24052
rect 20738 23884 20748 23940
rect 20804 23884 21532 23940
rect 21588 23884 22540 23940
rect 22596 23884 23548 23940
rect 23604 23884 23996 23940
rect 24052 23884 26684 23940
rect 26740 23884 26750 23940
rect 27234 23884 27244 23940
rect 27300 23884 27468 23940
rect 27524 23884 27534 23940
rect 31154 23884 31164 23940
rect 31220 23884 31388 23940
rect 31444 23884 31454 23940
rect 40562 23884 40572 23940
rect 40628 23884 41020 23940
rect 41076 23884 41356 23940
rect 41412 23884 41422 23940
rect 43652 23884 43932 23940
rect 43988 23884 43998 23940
rect 44818 23884 44828 23940
rect 44884 23884 47516 23940
rect 47572 23884 48636 23940
rect 48692 23884 49532 23940
rect 49588 23884 49598 23940
rect 43652 23828 43708 23884
rect 19170 23772 19180 23828
rect 19236 23772 21868 23828
rect 21924 23772 22316 23828
rect 22372 23772 23100 23828
rect 23156 23772 23166 23828
rect 24322 23772 24332 23828
rect 24388 23772 25788 23828
rect 25844 23772 27580 23828
rect 27636 23772 28028 23828
rect 28084 23772 28094 23828
rect 31714 23772 31724 23828
rect 31780 23772 33180 23828
rect 33236 23772 34188 23828
rect 34244 23772 34254 23828
rect 38770 23772 38780 23828
rect 38836 23772 39900 23828
rect 39956 23772 42812 23828
rect 42868 23772 43708 23828
rect 45714 23772 45724 23828
rect 45780 23772 46060 23828
rect 46116 23772 46844 23828
rect 46900 23772 48972 23828
rect 49028 23772 51324 23828
rect 51380 23772 51660 23828
rect 51716 23772 52668 23828
rect 52724 23772 54684 23828
rect 54740 23772 54750 23828
rect 11666 23660 11676 23716
rect 11732 23660 13468 23716
rect 13524 23660 15148 23716
rect 15204 23660 17500 23716
rect 17556 23660 18844 23716
rect 18900 23660 18910 23716
rect 23650 23660 23660 23716
rect 23716 23660 23996 23716
rect 24052 23660 24062 23716
rect 24434 23660 24444 23716
rect 24500 23660 25228 23716
rect 25284 23660 25294 23716
rect 25788 23660 32060 23716
rect 32116 23660 33068 23716
rect 33124 23660 33134 23716
rect 41458 23660 41468 23716
rect 41524 23660 42140 23716
rect 42196 23660 42206 23716
rect 50194 23660 50204 23716
rect 50260 23660 51212 23716
rect 51268 23660 52780 23716
rect 52836 23660 52846 23716
rect 25788 23604 25844 23660
rect 23202 23548 23212 23604
rect 23268 23548 25788 23604
rect 25844 23548 25854 23604
rect 26674 23548 26684 23604
rect 26740 23548 30772 23604
rect 31490 23548 31500 23604
rect 31556 23548 31948 23604
rect 32004 23548 33516 23604
rect 33572 23548 33582 23604
rect 34626 23548 34636 23604
rect 34692 23548 35532 23604
rect 35588 23548 36428 23604
rect 36484 23548 36494 23604
rect 41234 23548 41244 23604
rect 41300 23548 43596 23604
rect 43652 23548 45276 23604
rect 45332 23548 45342 23604
rect 49634 23548 49644 23604
rect 49700 23548 50428 23604
rect 50484 23548 50494 23604
rect 51090 23548 51100 23604
rect 51156 23548 54460 23604
rect 54516 23548 55132 23604
rect 55188 23548 55198 23604
rect 30716 23492 30772 23548
rect 50428 23492 50484 23548
rect 24658 23436 24668 23492
rect 24724 23436 26348 23492
rect 26404 23436 26414 23492
rect 30706 23436 30716 23492
rect 30772 23436 30782 23492
rect 32498 23436 32508 23492
rect 32564 23436 32844 23492
rect 32900 23436 32910 23492
rect 40002 23436 40012 23492
rect 40068 23436 40796 23492
rect 40852 23436 40862 23492
rect 50428 23436 51436 23492
rect 51492 23436 51660 23492
rect 51716 23436 51726 23492
rect 4466 23156 4476 23212
rect 4532 23156 4580 23212
rect 4636 23156 4684 23212
rect 4740 23156 4750 23212
rect 35186 23156 35196 23212
rect 35252 23156 35300 23212
rect 35356 23156 35404 23212
rect 35460 23156 35470 23212
rect 39330 22988 39340 23044
rect 39396 22988 40124 23044
rect 40180 22988 40190 23044
rect 26786 22876 26796 22932
rect 26852 22876 27468 22932
rect 27524 22876 27534 22932
rect 31154 22764 31164 22820
rect 31220 22764 33964 22820
rect 34020 22764 35532 22820
rect 35588 22764 36204 22820
rect 36260 22764 36270 22820
rect 24658 22540 24668 22596
rect 24724 22540 25116 22596
rect 25172 22540 25182 22596
rect 25554 22540 25564 22596
rect 25620 22540 26908 22596
rect 26964 22540 26974 22596
rect 30034 22540 30044 22596
rect 30100 22540 31164 22596
rect 31220 22540 31612 22596
rect 31668 22540 31678 22596
rect 37986 22540 37996 22596
rect 38052 22540 40572 22596
rect 40628 22540 41020 22596
rect 41076 22540 41244 22596
rect 41300 22540 41310 22596
rect 53442 22540 53452 22596
rect 53508 22540 54348 22596
rect 54404 22540 54414 22596
rect 30146 22428 30156 22484
rect 30212 22428 32284 22484
rect 32340 22428 32350 22484
rect 51874 22428 51884 22484
rect 51940 22428 54684 22484
rect 54740 22428 54750 22484
rect 56466 22428 56476 22484
rect 56532 22428 57148 22484
rect 57204 22428 57214 22484
rect 30706 22316 30716 22372
rect 30772 22316 31836 22372
rect 31892 22316 32620 22372
rect 32676 22316 32686 22372
rect 19826 22148 19836 22204
rect 19892 22148 19940 22204
rect 19996 22148 20044 22204
rect 20100 22148 20110 22204
rect 50546 22148 50556 22204
rect 50612 22148 50660 22204
rect 50716 22148 50764 22204
rect 50820 22148 50830 22204
rect 20132 21868 20300 21924
rect 20356 21868 20366 21924
rect 35970 21868 35980 21924
rect 36036 21868 36046 21924
rect 41346 21868 41356 21924
rect 41412 21868 41916 21924
rect 41972 21868 41982 21924
rect 54898 21868 54908 21924
rect 54964 21868 55468 21924
rect 20132 21700 20188 21868
rect 35980 21812 36036 21868
rect 55412 21812 55468 21868
rect 25666 21756 25676 21812
rect 25732 21756 26348 21812
rect 26404 21756 27356 21812
rect 27412 21756 28140 21812
rect 28196 21756 28700 21812
rect 28756 21756 31052 21812
rect 31108 21756 31118 21812
rect 34402 21756 34412 21812
rect 34468 21756 34972 21812
rect 35028 21756 35644 21812
rect 35700 21756 35710 21812
rect 35980 21756 37100 21812
rect 37156 21756 37166 21812
rect 41458 21756 41468 21812
rect 41524 21756 41804 21812
rect 41860 21756 42364 21812
rect 42420 21756 43708 21812
rect 49074 21756 49084 21812
rect 49140 21756 50876 21812
rect 50932 21756 51828 21812
rect 53218 21756 53228 21812
rect 53284 21756 55244 21812
rect 55300 21756 55310 21812
rect 55412 21756 56700 21812
rect 56756 21756 57708 21812
rect 57764 21756 57774 21812
rect 43652 21700 43708 21756
rect 51772 21700 51828 21756
rect 19842 21644 19852 21700
rect 19908 21644 20188 21700
rect 23202 21644 23212 21700
rect 23268 21644 23278 21700
rect 26450 21644 26460 21700
rect 26516 21644 26908 21700
rect 28578 21644 28588 21700
rect 28644 21644 30268 21700
rect 30324 21644 30334 21700
rect 41010 21644 41020 21700
rect 41076 21644 41580 21700
rect 41636 21644 41646 21700
rect 43652 21644 44604 21700
rect 44660 21644 45052 21700
rect 45108 21644 45724 21700
rect 45780 21644 45790 21700
rect 48514 21644 48524 21700
rect 48580 21644 48860 21700
rect 48916 21644 50988 21700
rect 51044 21644 51054 21700
rect 51762 21644 51772 21700
rect 51828 21644 54124 21700
rect 54180 21644 54190 21700
rect 23212 21588 23268 21644
rect 26852 21588 26908 21644
rect 55244 21588 55300 21756
rect 23212 21532 24668 21588
rect 24724 21532 25452 21588
rect 25508 21532 25518 21588
rect 26852 21532 27804 21588
rect 27860 21532 34076 21588
rect 34132 21532 34142 21588
rect 44146 21532 44156 21588
rect 44212 21532 45164 21588
rect 45220 21532 45500 21588
rect 45556 21532 45566 21588
rect 55244 21532 57036 21588
rect 57092 21532 57102 21588
rect 35074 21420 35084 21476
rect 35140 21420 36204 21476
rect 36260 21420 49756 21476
rect 49812 21420 49822 21476
rect 56018 21420 56028 21476
rect 56084 21420 57148 21476
rect 57204 21420 57214 21476
rect 51314 21308 51324 21364
rect 51380 21308 52892 21364
rect 52948 21308 52958 21364
rect 24210 21196 24220 21252
rect 24276 21196 25116 21252
rect 25172 21196 26796 21252
rect 26852 21196 28588 21252
rect 28644 21196 28654 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 26226 20972 26236 21028
rect 26292 20972 35196 21028
rect 35252 20972 35262 21028
rect 29810 20860 29820 20916
rect 29876 20860 30268 20916
rect 30324 20860 30334 20916
rect 23762 20748 23772 20804
rect 23828 20748 24668 20804
rect 24724 20748 24734 20804
rect 36306 20748 36316 20804
rect 36372 20748 37212 20804
rect 37268 20748 38332 20804
rect 38388 20748 38398 20804
rect 54114 20748 54124 20804
rect 54180 20748 54908 20804
rect 54964 20748 54974 20804
rect 56242 20748 56252 20804
rect 56308 20748 57036 20804
rect 57092 20748 57102 20804
rect 18498 20636 18508 20692
rect 18564 20636 20300 20692
rect 20356 20636 20366 20692
rect 30482 20636 30492 20692
rect 30548 20636 30828 20692
rect 30884 20636 32284 20692
rect 32340 20636 33068 20692
rect 33124 20636 34300 20692
rect 34356 20636 34366 20692
rect 41570 20636 41580 20692
rect 41636 20636 42252 20692
rect 42308 20636 42318 20692
rect 46386 20636 46396 20692
rect 46452 20636 48076 20692
rect 48132 20636 48142 20692
rect 49858 20636 49868 20692
rect 49924 20636 50540 20692
rect 50596 20636 52220 20692
rect 52276 20636 53116 20692
rect 53172 20636 53182 20692
rect 53778 20636 53788 20692
rect 53844 20636 55804 20692
rect 55860 20636 55870 20692
rect 19282 20524 19292 20580
rect 19348 20524 21532 20580
rect 21588 20524 21598 20580
rect 22082 20524 22092 20580
rect 22148 20524 22158 20580
rect 41458 20524 41468 20580
rect 41524 20524 43484 20580
rect 43540 20524 43550 20580
rect 45938 20524 45948 20580
rect 46004 20524 47628 20580
rect 47684 20524 47694 20580
rect 22092 20468 22148 20524
rect 19730 20412 19740 20468
rect 19796 20412 22148 20468
rect 27234 20412 27244 20468
rect 27300 20412 28476 20468
rect 28532 20412 28542 20468
rect 29474 20412 29484 20468
rect 29540 20412 30380 20468
rect 30436 20412 30828 20468
rect 30884 20412 31276 20468
rect 31332 20412 33516 20468
rect 33572 20412 37100 20468
rect 37156 20412 38332 20468
rect 38388 20412 38398 20468
rect 43362 20412 43372 20468
rect 43428 20412 43596 20468
rect 43652 20412 43662 20468
rect 45714 20412 45724 20468
rect 45780 20412 47740 20468
rect 47796 20412 49532 20468
rect 49588 20412 49598 20468
rect 50978 20412 50988 20468
rect 51044 20412 53340 20468
rect 53396 20412 53406 20468
rect 19842 20300 19852 20356
rect 19908 20300 20244 20356
rect 29138 20300 29148 20356
rect 29204 20300 29820 20356
rect 29876 20300 31836 20356
rect 31892 20300 33852 20356
rect 33908 20300 35196 20356
rect 35252 20300 38668 20356
rect 38724 20300 40012 20356
rect 40068 20300 40796 20356
rect 40852 20300 42700 20356
rect 42756 20300 46676 20356
rect 19826 20132 19836 20188
rect 19892 20132 19940 20188
rect 19996 20132 20044 20188
rect 20100 20132 20110 20188
rect 20188 20132 20244 20300
rect 46620 20244 46676 20300
rect 47516 20300 48636 20356
rect 48692 20300 50204 20356
rect 50260 20300 50270 20356
rect 47516 20244 47572 20300
rect 20738 20188 20748 20244
rect 20804 20188 22764 20244
rect 22820 20188 24108 20244
rect 24164 20188 25340 20244
rect 25396 20188 25406 20244
rect 27458 20188 27468 20244
rect 27524 20188 27804 20244
rect 27860 20188 27870 20244
rect 40898 20188 40908 20244
rect 40964 20188 41580 20244
rect 41636 20188 41646 20244
rect 43474 20188 43484 20244
rect 43540 20188 44156 20244
rect 44212 20188 44222 20244
rect 46386 20188 46396 20244
rect 46452 20188 46676 20244
rect 46620 20132 46676 20188
rect 47012 20188 47516 20244
rect 47572 20188 47582 20244
rect 47012 20132 47068 20188
rect 50546 20132 50556 20188
rect 50612 20132 50660 20188
rect 50716 20132 50764 20188
rect 50820 20132 50830 20188
rect 20188 20076 20636 20132
rect 20692 20076 22316 20132
rect 22372 20076 22876 20132
rect 22932 20076 22942 20132
rect 33394 20076 33404 20132
rect 33460 20076 33964 20132
rect 34020 20076 34030 20132
rect 46620 20076 46732 20132
rect 46788 20076 47068 20132
rect 22194 19852 22204 19908
rect 22260 19852 26012 19908
rect 26068 19852 29260 19908
rect 29316 19852 30380 19908
rect 30436 19852 30446 19908
rect 20178 19740 20188 19796
rect 20244 19740 21084 19796
rect 21140 19740 21756 19796
rect 21812 19740 21822 19796
rect 27346 19740 27356 19796
rect 27412 19740 29596 19796
rect 29652 19740 32060 19796
rect 32116 19740 32844 19796
rect 32900 19740 32910 19796
rect 41346 19740 41356 19796
rect 41412 19740 41804 19796
rect 41860 19740 41870 19796
rect 46946 19740 46956 19796
rect 47012 19740 47628 19796
rect 47684 19740 47694 19796
rect 30258 19628 30268 19684
rect 30324 19628 31052 19684
rect 31108 19628 31724 19684
rect 31780 19628 32284 19684
rect 32340 19628 32350 19684
rect 49746 19628 49756 19684
rect 49812 19628 49980 19684
rect 50036 19628 50876 19684
rect 50932 19628 51548 19684
rect 51604 19628 53228 19684
rect 53284 19628 53294 19684
rect 24546 19516 24556 19572
rect 24612 19516 26908 19572
rect 26964 19516 26974 19572
rect 40226 19404 40236 19460
rect 40292 19404 41244 19460
rect 41300 19404 41310 19460
rect 42690 19404 42700 19460
rect 42756 19404 44268 19460
rect 44324 19404 44334 19460
rect 35634 19292 35644 19348
rect 35700 19292 41580 19348
rect 41636 19292 41646 19348
rect 29586 19180 29596 19236
rect 29652 19180 29932 19236
rect 29988 19180 29998 19236
rect 4466 19124 4476 19180
rect 4532 19124 4580 19180
rect 4636 19124 4684 19180
rect 4740 19124 4750 19180
rect 35186 19124 35196 19180
rect 35252 19124 35300 19180
rect 35356 19124 35404 19180
rect 35460 19124 35470 19180
rect 18386 19068 18396 19124
rect 18452 19068 19516 19124
rect 19572 19068 20188 19124
rect 20244 19068 20254 19124
rect 20290 18956 20300 19012
rect 20356 18956 21420 19012
rect 21476 18956 21486 19012
rect 23202 18844 23212 18900
rect 23268 18844 25228 18900
rect 25284 18844 26684 18900
rect 26740 18844 26750 18900
rect 49970 18844 49980 18900
rect 50036 18844 52556 18900
rect 52612 18844 52622 18900
rect 20132 18732 21420 18788
rect 21476 18732 21486 18788
rect 28018 18732 28028 18788
rect 28084 18732 28588 18788
rect 28644 18732 29484 18788
rect 29540 18732 29550 18788
rect 49074 18732 49084 18788
rect 49140 18732 50876 18788
rect 50932 18732 50942 18788
rect 20132 18676 20188 18732
rect 17490 18620 17500 18676
rect 17556 18620 18284 18676
rect 18340 18620 18350 18676
rect 19730 18620 19740 18676
rect 19796 18620 20188 18676
rect 35970 18620 35980 18676
rect 36036 18620 36316 18676
rect 36372 18620 37660 18676
rect 37716 18620 38332 18676
rect 38388 18620 39340 18676
rect 39396 18620 41356 18676
rect 41412 18620 41422 18676
rect 48850 18620 48860 18676
rect 48916 18620 50092 18676
rect 50148 18620 50158 18676
rect 16594 18508 16604 18564
rect 16660 18508 17724 18564
rect 17780 18508 18508 18564
rect 18564 18508 18956 18564
rect 19012 18508 19022 18564
rect 20738 18508 20748 18564
rect 20804 18508 22876 18564
rect 22932 18508 22942 18564
rect 36194 18508 36204 18564
rect 36260 18508 37548 18564
rect 37604 18508 37614 18564
rect 38546 18508 38556 18564
rect 38612 18508 40908 18564
rect 40964 18508 40974 18564
rect 45602 18508 45612 18564
rect 45668 18508 47068 18564
rect 47124 18508 47740 18564
rect 47796 18508 47964 18564
rect 48020 18508 49420 18564
rect 49476 18508 49486 18564
rect 18274 18396 18284 18452
rect 18340 18396 19180 18452
rect 19236 18396 19246 18452
rect 25666 18396 25676 18452
rect 25732 18396 29820 18452
rect 29876 18396 29886 18452
rect 34738 18396 34748 18452
rect 34804 18396 35308 18452
rect 35364 18396 35374 18452
rect 40786 18396 40796 18452
rect 40852 18396 41244 18452
rect 41300 18396 41310 18452
rect 43474 18396 43484 18452
rect 43540 18396 45724 18452
rect 45780 18396 46284 18452
rect 46340 18396 46732 18452
rect 46788 18396 46798 18452
rect 34748 18340 34804 18396
rect 28802 18284 28812 18340
rect 28868 18284 34804 18340
rect 36418 18284 36428 18340
rect 36484 18284 38108 18340
rect 38164 18284 38174 18340
rect 19826 18116 19836 18172
rect 19892 18116 19940 18172
rect 19996 18116 20044 18172
rect 20100 18116 20110 18172
rect 50546 18116 50556 18172
rect 50612 18116 50660 18172
rect 50716 18116 50764 18172
rect 50820 18116 50830 18172
rect 47394 17948 47404 18004
rect 47460 17948 50540 18004
rect 50596 17948 50606 18004
rect 20132 17836 23548 17892
rect 23604 17836 23614 17892
rect 24434 17836 24444 17892
rect 24500 17836 26348 17892
rect 26404 17836 26414 17892
rect 30818 17836 30828 17892
rect 30884 17836 46620 17892
rect 46676 17836 46686 17892
rect 48178 17836 48188 17892
rect 48244 17836 49532 17892
rect 49588 17836 49598 17892
rect 20132 17668 20188 17836
rect 26562 17724 26572 17780
rect 26628 17724 26638 17780
rect 41346 17724 41356 17780
rect 41412 17724 42924 17780
rect 42980 17724 42990 17780
rect 19954 17612 19964 17668
rect 20020 17612 20188 17668
rect 20402 17612 20412 17668
rect 20468 17612 20478 17668
rect 20412 17556 20468 17612
rect 26572 17556 26628 17724
rect 43922 17612 43932 17668
rect 43988 17612 45276 17668
rect 45332 17612 45948 17668
rect 46004 17612 47180 17668
rect 47236 17612 47246 17668
rect 16818 17500 16828 17556
rect 16884 17500 18284 17556
rect 18340 17500 18350 17556
rect 18722 17500 18732 17556
rect 18788 17500 20468 17556
rect 25330 17500 25340 17556
rect 25396 17500 27356 17556
rect 27412 17500 27692 17556
rect 27748 17500 27758 17556
rect 4466 17108 4476 17164
rect 4532 17108 4580 17164
rect 4636 17108 4684 17164
rect 4740 17108 4750 17164
rect 35186 17108 35196 17164
rect 35252 17108 35300 17164
rect 35356 17108 35404 17164
rect 35460 17108 35470 17164
rect 28802 16828 28812 16884
rect 28868 16828 29372 16884
rect 29428 16828 29438 16884
rect 42914 16828 42924 16884
rect 42980 16828 43708 16884
rect 43652 16772 43708 16828
rect 19282 16716 19292 16772
rect 19348 16716 20076 16772
rect 20132 16716 21980 16772
rect 22036 16716 23772 16772
rect 23828 16716 23838 16772
rect 24994 16716 25004 16772
rect 25060 16716 27244 16772
rect 27300 16716 29260 16772
rect 29316 16716 29326 16772
rect 34962 16716 34972 16772
rect 35028 16716 36764 16772
rect 36820 16716 36830 16772
rect 37426 16716 37436 16772
rect 37492 16716 39676 16772
rect 39732 16716 39742 16772
rect 43652 16716 44828 16772
rect 44884 16716 44894 16772
rect 47730 16716 47740 16772
rect 47796 16716 49308 16772
rect 49364 16716 49756 16772
rect 49812 16716 49822 16772
rect 25004 16660 25060 16716
rect 15026 16604 15036 16660
rect 15092 16604 17612 16660
rect 17668 16604 18620 16660
rect 18676 16604 20244 16660
rect 20514 16604 20524 16660
rect 20580 16604 21308 16660
rect 21364 16604 25060 16660
rect 28018 16604 28028 16660
rect 28084 16604 30492 16660
rect 30548 16604 30558 16660
rect 38210 16604 38220 16660
rect 38276 16604 43036 16660
rect 43092 16604 43102 16660
rect 47506 16604 47516 16660
rect 47572 16604 48972 16660
rect 49028 16604 50316 16660
rect 50372 16604 50382 16660
rect 50866 16604 50876 16660
rect 50932 16604 52556 16660
rect 52612 16604 52622 16660
rect 20188 16436 20244 16604
rect 37762 16492 37772 16548
rect 37828 16492 39452 16548
rect 39508 16492 43932 16548
rect 43988 16492 43998 16548
rect 20178 16380 20188 16436
rect 20244 16380 21868 16436
rect 21924 16380 22988 16436
rect 23044 16380 23054 16436
rect 44706 16380 44716 16436
rect 44772 16380 46060 16436
rect 46116 16380 46126 16436
rect 51650 16380 51660 16436
rect 51716 16380 52556 16436
rect 52612 16380 52622 16436
rect 53218 16380 53228 16436
rect 53284 16380 54908 16436
rect 54964 16380 54974 16436
rect 19170 16268 19180 16324
rect 19236 16268 21084 16324
rect 21140 16268 21150 16324
rect 27570 16268 27580 16324
rect 27636 16268 28028 16324
rect 28084 16268 28094 16324
rect 50194 16268 50204 16324
rect 50260 16268 50764 16324
rect 50820 16268 51772 16324
rect 51828 16268 51838 16324
rect 19826 16100 19836 16156
rect 19892 16100 19940 16156
rect 19996 16100 20044 16156
rect 20100 16100 20110 16156
rect 50546 16100 50556 16156
rect 50612 16100 50660 16156
rect 50716 16100 50764 16156
rect 50820 16100 50830 16156
rect 20738 15820 20748 15876
rect 20804 15820 21644 15876
rect 21700 15820 21710 15876
rect 22978 15820 22988 15876
rect 23044 15820 23940 15876
rect 24210 15820 24220 15876
rect 24276 15820 25340 15876
rect 25396 15820 25406 15876
rect 41682 15820 41692 15876
rect 41748 15820 42364 15876
rect 42420 15820 42430 15876
rect 47170 15820 47180 15876
rect 47236 15820 51212 15876
rect 51268 15820 52892 15876
rect 52948 15820 52958 15876
rect 23884 15764 23940 15820
rect 23874 15708 23884 15764
rect 23940 15708 24668 15764
rect 24724 15708 25788 15764
rect 25844 15708 25854 15764
rect 36194 15708 36204 15764
rect 36260 15708 37436 15764
rect 37492 15708 37502 15764
rect 37986 15708 37996 15764
rect 38052 15708 39564 15764
rect 39620 15708 39630 15764
rect 41010 15708 41020 15764
rect 41076 15708 41580 15764
rect 41636 15708 41646 15764
rect 43474 15708 43484 15764
rect 43540 15708 44940 15764
rect 44996 15708 45006 15764
rect 51762 15708 51772 15764
rect 51828 15708 52780 15764
rect 52836 15708 54572 15764
rect 54628 15708 54638 15764
rect 20850 15596 20860 15652
rect 20916 15596 21308 15652
rect 21364 15596 22988 15652
rect 23044 15596 23054 15652
rect 24322 15596 24332 15652
rect 24388 15596 26012 15652
rect 26068 15596 27076 15652
rect 35074 15596 35084 15652
rect 35140 15596 38332 15652
rect 38388 15596 38398 15652
rect 47058 15596 47068 15652
rect 47124 15596 47964 15652
rect 48020 15596 49756 15652
rect 49812 15596 50988 15652
rect 51044 15596 54236 15652
rect 54292 15596 54302 15652
rect 27020 15316 27076 15596
rect 27458 15372 27468 15428
rect 27524 15372 28364 15428
rect 28420 15372 28430 15428
rect 41682 15372 41692 15428
rect 41748 15372 42364 15428
rect 42420 15372 42430 15428
rect 27010 15260 27020 15316
rect 27076 15260 28476 15316
rect 28532 15260 28542 15316
rect 50530 15260 50540 15316
rect 50596 15260 51660 15316
rect 51716 15260 53340 15316
rect 53396 15260 53406 15316
rect 27430 15148 27468 15204
rect 27524 15148 27534 15204
rect 28588 15148 29484 15204
rect 29540 15148 31276 15204
rect 31332 15148 32284 15204
rect 32340 15148 32350 15204
rect 49970 15148 49980 15204
rect 50036 15148 50764 15204
rect 50820 15148 50830 15204
rect 4466 15092 4476 15148
rect 4532 15092 4580 15148
rect 4636 15092 4684 15148
rect 4740 15092 4750 15148
rect 28588 15092 28644 15148
rect 35186 15092 35196 15148
rect 35252 15092 35300 15148
rect 35356 15092 35404 15148
rect 35460 15092 35470 15148
rect 27794 15036 27804 15092
rect 27860 15036 28644 15092
rect 30594 15036 30604 15092
rect 30660 15036 31836 15092
rect 31892 15036 31902 15092
rect 41458 15036 41468 15092
rect 41524 15036 42700 15092
rect 42756 15036 42766 15092
rect 37874 14924 37884 14980
rect 37940 14924 38668 14980
rect 38724 14924 38734 14980
rect 26852 14812 28812 14868
rect 28868 14812 29708 14868
rect 29764 14812 30604 14868
rect 30660 14812 32732 14868
rect 32788 14812 33068 14868
rect 33124 14812 34860 14868
rect 34916 14812 34926 14868
rect 20290 14700 20300 14756
rect 20356 14700 20972 14756
rect 21028 14700 22428 14756
rect 22484 14700 22494 14756
rect 26786 14700 26796 14756
rect 26852 14700 26908 14812
rect 36418 14700 36428 14756
rect 36484 14700 38220 14756
rect 38276 14700 38286 14756
rect 39218 14700 39228 14756
rect 39284 14700 39676 14756
rect 39732 14700 40236 14756
rect 40292 14700 40302 14756
rect 43810 14700 43820 14756
rect 43876 14700 45836 14756
rect 45892 14700 45902 14756
rect 50978 14700 50988 14756
rect 51044 14700 52108 14756
rect 52164 14700 52174 14756
rect 24658 14588 24668 14644
rect 24724 14588 26012 14644
rect 26068 14588 26078 14644
rect 26898 14588 26908 14644
rect 26964 14588 27468 14644
rect 27524 14588 33180 14644
rect 33236 14588 33246 14644
rect 37090 14588 37100 14644
rect 37156 14588 37324 14644
rect 37380 14588 37390 14644
rect 43652 14588 45388 14644
rect 45444 14588 45454 14644
rect 52546 14588 52556 14644
rect 52612 14588 53228 14644
rect 53284 14588 53294 14644
rect 43652 14532 43708 14588
rect 24434 14476 24444 14532
rect 24500 14476 25452 14532
rect 25508 14476 25518 14532
rect 26226 14476 26236 14532
rect 26292 14476 27748 14532
rect 31826 14476 31836 14532
rect 31892 14476 34076 14532
rect 34132 14476 35644 14532
rect 35700 14476 37772 14532
rect 37828 14476 37838 14532
rect 43474 14476 43484 14532
rect 43540 14476 43708 14532
rect 44930 14476 44940 14532
rect 44996 14476 46396 14532
rect 46452 14476 47180 14532
rect 47236 14476 47246 14532
rect 25452 14420 25508 14476
rect 27692 14420 27748 14476
rect 19842 14364 19852 14420
rect 19908 14364 20188 14420
rect 25452 14364 25788 14420
rect 25844 14364 26348 14420
rect 26404 14364 26908 14420
rect 27682 14364 27692 14420
rect 27748 14364 27758 14420
rect 28130 14364 28140 14420
rect 28196 14364 29260 14420
rect 29316 14364 29326 14420
rect 44258 14364 44268 14420
rect 44324 14364 45612 14420
rect 45668 14364 46732 14420
rect 46788 14364 48860 14420
rect 48916 14364 50092 14420
rect 50148 14364 50158 14420
rect 20132 14308 20188 14364
rect 26852 14308 26908 14364
rect 28140 14308 28196 14364
rect 20132 14252 21420 14308
rect 21476 14252 21486 14308
rect 22306 14252 22316 14308
rect 22372 14252 26236 14308
rect 26292 14252 26572 14308
rect 26628 14252 26638 14308
rect 26852 14252 28196 14308
rect 33506 14252 33516 14308
rect 33572 14252 37212 14308
rect 37268 14252 37278 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 21410 13804 21420 13860
rect 21476 13804 23212 13860
rect 23268 13804 24220 13860
rect 24276 13804 24444 13860
rect 24500 13804 24510 13860
rect 25442 13804 25452 13860
rect 25508 13804 26684 13860
rect 26740 13804 26908 13860
rect 29250 13804 29260 13860
rect 29316 13804 30380 13860
rect 30436 13804 32060 13860
rect 32116 13804 37324 13860
rect 37380 13804 37390 13860
rect 41346 13804 41356 13860
rect 41412 13804 42364 13860
rect 42420 13804 42430 13860
rect 51202 13804 51212 13860
rect 51268 13804 52444 13860
rect 52500 13804 52510 13860
rect 21634 13692 21644 13748
rect 21700 13692 22316 13748
rect 22372 13692 22382 13748
rect 26852 13636 26908 13804
rect 33170 13692 33180 13748
rect 33236 13692 33740 13748
rect 33796 13692 33806 13748
rect 40338 13692 40348 13748
rect 40404 13692 41020 13748
rect 41076 13692 41086 13748
rect 26852 13580 28140 13636
rect 28196 13580 28812 13636
rect 28868 13580 30044 13636
rect 30100 13580 30110 13636
rect 32498 13580 32508 13636
rect 32564 13580 33964 13636
rect 34020 13580 34748 13636
rect 34804 13580 38108 13636
rect 38164 13580 38174 13636
rect 17602 13468 17612 13524
rect 17668 13468 18620 13524
rect 18676 13468 19404 13524
rect 19460 13468 19470 13524
rect 28578 13468 28588 13524
rect 28644 13468 30156 13524
rect 30212 13468 30828 13524
rect 30884 13468 33628 13524
rect 33684 13468 33694 13524
rect 34066 13468 34076 13524
rect 34132 13468 34860 13524
rect 34916 13468 34926 13524
rect 38546 13468 38556 13524
rect 38612 13468 39004 13524
rect 39060 13468 39900 13524
rect 39956 13468 39966 13524
rect 27346 13356 27356 13412
rect 27412 13356 28028 13412
rect 28084 13356 32844 13412
rect 32900 13356 32910 13412
rect 4466 13076 4476 13132
rect 4532 13076 4580 13132
rect 4636 13076 4684 13132
rect 4740 13076 4750 13132
rect 35186 13076 35196 13132
rect 35252 13076 35300 13132
rect 35356 13076 35404 13132
rect 35460 13076 35470 13132
rect 28354 12908 28364 12964
rect 28420 12908 31948 12964
rect 32004 12908 32014 12964
rect 36418 12796 36428 12852
rect 36484 12796 37884 12852
rect 37940 12796 37950 12852
rect 38098 12796 38108 12852
rect 38164 12796 39676 12852
rect 39732 12796 43260 12852
rect 43316 12796 43708 12852
rect 43810 12796 43820 12852
rect 43876 12796 46284 12852
rect 46340 12796 47740 12852
rect 47796 12796 47806 12852
rect 32834 12684 32844 12740
rect 32900 12684 34524 12740
rect 34580 12684 34590 12740
rect 43652 12628 43708 12796
rect 37090 12572 37100 12628
rect 37156 12572 37324 12628
rect 37380 12572 38668 12628
rect 38724 12572 39004 12628
rect 39060 12572 39070 12628
rect 39330 12572 39340 12628
rect 39396 12572 40012 12628
rect 40068 12572 40078 12628
rect 43652 12572 44492 12628
rect 44548 12572 49980 12628
rect 50036 12572 50046 12628
rect 42130 12460 42140 12516
rect 42196 12460 42924 12516
rect 42980 12460 43484 12516
rect 43540 12460 43550 12516
rect 44930 12460 44940 12516
rect 44996 12460 47068 12516
rect 47124 12460 47964 12516
rect 48020 12460 48030 12516
rect 18274 12236 18284 12292
rect 18340 12236 21308 12292
rect 21364 12236 21374 12292
rect 19826 12068 19836 12124
rect 19892 12068 19940 12124
rect 19996 12068 20044 12124
rect 20100 12068 20110 12124
rect 50546 12068 50556 12124
rect 50612 12068 50660 12124
rect 50716 12068 50764 12124
rect 50820 12068 50830 12124
rect 22866 11900 22876 11956
rect 22932 11900 24332 11956
rect 24388 11900 25004 11956
rect 25060 11900 25070 11956
rect 26852 11788 27132 11844
rect 27188 11788 27804 11844
rect 27860 11788 28028 11844
rect 28084 11788 28094 11844
rect 32834 11788 32844 11844
rect 32900 11788 32910 11844
rect 26852 11732 26908 11788
rect 23090 11676 23100 11732
rect 23156 11676 25116 11732
rect 25172 11676 25182 11732
rect 25330 11676 25340 11732
rect 25396 11676 26908 11732
rect 32844 11732 32900 11788
rect 32844 11676 34076 11732
rect 34132 11676 34142 11732
rect 44034 11676 44044 11732
rect 44100 11676 46620 11732
rect 46676 11676 46686 11732
rect 25340 11620 25396 11676
rect 22306 11564 22316 11620
rect 22372 11564 23548 11620
rect 23604 11564 23614 11620
rect 24210 11564 24220 11620
rect 24276 11564 25396 11620
rect 20626 11452 20636 11508
rect 20692 11452 23436 11508
rect 23492 11452 23502 11508
rect 24994 11452 25004 11508
rect 25060 11452 26348 11508
rect 26404 11452 26414 11508
rect 21970 11340 21980 11396
rect 22036 11340 23324 11396
rect 23380 11340 23390 11396
rect 4466 11060 4476 11116
rect 4532 11060 4580 11116
rect 4636 11060 4684 11116
rect 4740 11060 4750 11116
rect 35186 11060 35196 11116
rect 35252 11060 35300 11116
rect 35356 11060 35404 11116
rect 35460 11060 35470 11116
rect 20132 10780 20636 10836
rect 20692 10780 21980 10836
rect 22036 10780 22046 10836
rect 20132 10612 20188 10780
rect 28130 10668 28140 10724
rect 28196 10668 30044 10724
rect 30100 10668 30716 10724
rect 30772 10668 30782 10724
rect 19058 10556 19068 10612
rect 19124 10556 19852 10612
rect 19908 10556 20188 10612
rect 21074 10556 21084 10612
rect 21140 10556 21980 10612
rect 22036 10556 22046 10612
rect 37314 10556 37324 10612
rect 37380 10556 38332 10612
rect 38388 10556 39228 10612
rect 39284 10556 39676 10612
rect 39732 10556 40348 10612
rect 40404 10556 40414 10612
rect 20132 10444 21308 10500
rect 21364 10444 21374 10500
rect 28242 10444 28252 10500
rect 28308 10444 29708 10500
rect 29764 10444 31276 10500
rect 31332 10444 31342 10500
rect 32386 10444 32396 10500
rect 32452 10444 33068 10500
rect 33124 10444 33134 10500
rect 39442 10444 39452 10500
rect 39508 10444 40124 10500
rect 40180 10444 40190 10500
rect 43586 10444 43596 10500
rect 43652 10444 48076 10500
rect 48132 10444 48142 10500
rect 20132 10388 20188 10444
rect 19730 10332 19740 10388
rect 19796 10332 20188 10388
rect 22418 10332 22428 10388
rect 22484 10332 24108 10388
rect 24164 10332 24174 10388
rect 32498 10332 32508 10388
rect 32564 10332 33740 10388
rect 33796 10332 33806 10388
rect 16370 10108 16380 10164
rect 16436 10108 17500 10164
rect 17556 10108 18396 10164
rect 18452 10108 18462 10164
rect 22866 10108 22876 10164
rect 22932 10108 27468 10164
rect 27524 10108 27534 10164
rect 19826 10052 19836 10108
rect 19892 10052 19940 10108
rect 19996 10052 20044 10108
rect 20100 10052 20110 10108
rect 50546 10052 50556 10108
rect 50612 10052 50660 10108
rect 50716 10052 50764 10108
rect 50820 10052 50830 10108
rect 16930 9996 16940 10052
rect 16996 9996 18284 10052
rect 18340 9996 18350 10052
rect 24210 9996 24220 10052
rect 24276 9996 25340 10052
rect 25396 9996 27020 10052
rect 27076 9996 27086 10052
rect 32162 9772 32172 9828
rect 32228 9772 41916 9828
rect 41972 9772 41982 9828
rect 28578 9660 28588 9716
rect 28644 9660 29260 9716
rect 29316 9660 29596 9716
rect 29652 9660 30604 9716
rect 30660 9660 30670 9716
rect 19618 9548 19628 9604
rect 19684 9548 20300 9604
rect 20356 9548 20636 9604
rect 20692 9548 20702 9604
rect 32722 9548 32732 9604
rect 32788 9548 34748 9604
rect 34804 9548 36092 9604
rect 36148 9548 37324 9604
rect 37380 9548 37390 9604
rect 40226 9548 40236 9604
rect 40292 9548 40908 9604
rect 40964 9548 40974 9604
rect 18274 9436 18284 9492
rect 18340 9436 18956 9492
rect 19012 9436 20188 9492
rect 20244 9436 20254 9492
rect 35634 9436 35644 9492
rect 35700 9436 36540 9492
rect 36596 9436 37660 9492
rect 37716 9436 37726 9492
rect 37202 9324 37212 9380
rect 37268 9324 41244 9380
rect 41300 9324 41310 9380
rect 4466 9044 4476 9100
rect 4532 9044 4580 9100
rect 4636 9044 4684 9100
rect 4740 9044 4750 9100
rect 35186 9044 35196 9100
rect 35252 9044 35300 9100
rect 35356 9044 35404 9100
rect 35460 9044 35470 9100
rect 19506 8764 19516 8820
rect 19572 8764 20524 8820
rect 20580 8764 23884 8820
rect 23940 8764 24668 8820
rect 24724 8764 24734 8820
rect 19842 8652 19852 8708
rect 19908 8652 20860 8708
rect 20916 8652 21532 8708
rect 21588 8652 21598 8708
rect 29362 8652 29372 8708
rect 29428 8652 30268 8708
rect 30324 8652 30334 8708
rect 30706 8652 30716 8708
rect 30772 8652 32060 8708
rect 32116 8652 33292 8708
rect 33348 8652 35644 8708
rect 35700 8652 35710 8708
rect 36194 8652 36204 8708
rect 36260 8652 40012 8708
rect 40068 8652 40078 8708
rect 40450 8652 40460 8708
rect 40516 8652 42028 8708
rect 42084 8652 42094 8708
rect 40012 8596 40068 8652
rect 20178 8540 20188 8596
rect 20244 8540 20748 8596
rect 20804 8540 20814 8596
rect 23650 8540 23660 8596
rect 23716 8540 25116 8596
rect 25172 8540 25182 8596
rect 27234 8540 27244 8596
rect 27300 8540 29148 8596
rect 29204 8540 29820 8596
rect 29876 8540 31388 8596
rect 31444 8540 31454 8596
rect 40012 8540 41020 8596
rect 41076 8540 43260 8596
rect 43316 8540 43326 8596
rect 18946 8428 18956 8484
rect 19012 8428 19852 8484
rect 19908 8428 20636 8484
rect 20692 8428 22204 8484
rect 22260 8428 22270 8484
rect 31154 8428 31164 8484
rect 31220 8428 32732 8484
rect 32788 8428 32798 8484
rect 38770 8428 38780 8484
rect 38836 8428 40236 8484
rect 40292 8428 41468 8484
rect 41524 8428 41534 8484
rect 37650 8316 37660 8372
rect 37716 8316 40124 8372
rect 40180 8316 41916 8372
rect 41972 8316 41982 8372
rect 33506 8092 33516 8148
rect 33572 8092 35308 8148
rect 35364 8092 36652 8148
rect 36708 8092 38780 8148
rect 38836 8092 38846 8148
rect 19826 8036 19836 8092
rect 19892 8036 19940 8092
rect 19996 8036 20044 8092
rect 20100 8036 20110 8092
rect 50546 8036 50556 8092
rect 50612 8036 50660 8092
rect 50716 8036 50764 8092
rect 50820 8036 50830 8092
rect 24882 7868 24892 7924
rect 24948 7868 30268 7924
rect 30324 7868 30334 7924
rect 27346 7756 27356 7812
rect 27412 7756 34076 7812
rect 34132 7756 34142 7812
rect 22530 7644 22540 7700
rect 22596 7644 23996 7700
rect 24052 7644 24062 7700
rect 21522 7532 21532 7588
rect 21588 7532 22988 7588
rect 23044 7532 23054 7588
rect 24994 7532 25004 7588
rect 25060 7532 26124 7588
rect 26180 7532 26190 7588
rect 32498 7532 32508 7588
rect 32564 7532 33740 7588
rect 33796 7532 33806 7588
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 0 6804 800 6832
rect 0 6748 4620 6804
rect 4676 6748 4686 6804
rect 0 6720 800 6748
rect 20402 6636 20412 6692
rect 20468 6636 21980 6692
rect 22036 6636 22046 6692
rect 25106 6636 25116 6692
rect 25172 6636 27468 6692
rect 27524 6636 28924 6692
rect 28980 6636 30380 6692
rect 30436 6636 30446 6692
rect 32722 6636 32732 6692
rect 32788 6636 33068 6692
rect 33124 6636 33852 6692
rect 33908 6636 33918 6692
rect 21980 6580 22036 6636
rect 19394 6524 19404 6580
rect 19460 6524 20076 6580
rect 20132 6524 21196 6580
rect 21252 6524 21262 6580
rect 21980 6524 24332 6580
rect 24388 6524 24668 6580
rect 24724 6524 25228 6580
rect 25284 6524 25900 6580
rect 25956 6524 27020 6580
rect 27076 6524 27086 6580
rect 28802 6524 28812 6580
rect 28868 6524 29260 6580
rect 29316 6524 29326 6580
rect 31826 6524 31836 6580
rect 31892 6524 33628 6580
rect 33684 6524 33694 6580
rect 20132 6412 20636 6468
rect 20692 6412 20702 6468
rect 31602 6412 31612 6468
rect 31668 6412 32396 6468
rect 32452 6412 34972 6468
rect 35028 6412 35038 6468
rect 20132 6356 20188 6412
rect 4162 6300 4172 6356
rect 4228 6300 4238 6356
rect 18162 6300 18172 6356
rect 18228 6300 20188 6356
rect 20514 6300 20524 6356
rect 20580 6300 22204 6356
rect 22260 6300 22270 6356
rect 24322 6300 24332 6356
rect 24388 6300 25340 6356
rect 25396 6300 25406 6356
rect 0 6132 800 6160
rect 4172 6132 4228 6300
rect 0 6076 4228 6132
rect 0 6048 800 6076
rect 19826 6020 19836 6076
rect 19892 6020 19940 6076
rect 19996 6020 20044 6076
rect 20100 6020 20110 6076
rect 50546 6020 50556 6076
rect 50612 6020 50660 6076
rect 50716 6020 50764 6076
rect 50820 6020 50830 6076
rect 27906 5740 27916 5796
rect 27972 5740 29148 5796
rect 29204 5740 29820 5796
rect 29876 5740 29886 5796
rect 26338 5404 26348 5460
rect 26404 5404 28476 5460
rect 28532 5404 28542 5460
rect 35186 5404 35196 5460
rect 35252 5404 36092 5460
rect 36148 5404 36158 5460
rect 4466 5012 4476 5068
rect 4532 5012 4580 5068
rect 4636 5012 4684 5068
rect 4740 5012 4750 5068
rect 35186 5012 35196 5068
rect 35252 5012 35300 5068
rect 35356 5012 35404 5068
rect 35460 5012 35470 5068
rect 23986 4620 23996 4676
rect 24052 4620 25452 4676
rect 25508 4620 25518 4676
rect 25890 4620 25900 4676
rect 25956 4620 26684 4676
rect 26740 4620 27692 4676
rect 27748 4620 27758 4676
rect 19826 4004 19836 4060
rect 19892 4004 19940 4060
rect 19996 4004 20044 4060
rect 20100 4004 20110 4060
rect 50546 4004 50556 4060
rect 50612 4004 50660 4060
rect 50716 4004 50764 4060
rect 50820 4004 50830 4060
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55412 4532 55468
rect 4580 55412 4636 55468
rect 4684 55412 4740 55468
rect 35196 55412 35252 55468
rect 35300 55412 35356 55468
rect 35404 55412 35460 55468
rect 19836 54404 19892 54460
rect 19940 54404 19996 54460
rect 20044 54404 20100 54460
rect 50556 54404 50612 54460
rect 50660 54404 50716 54460
rect 50764 54404 50820 54460
rect 4476 53396 4532 53452
rect 4580 53396 4636 53452
rect 4684 53396 4740 53452
rect 35196 53396 35252 53452
rect 35300 53396 35356 53452
rect 35404 53396 35460 53452
rect 19836 52388 19892 52444
rect 19940 52388 19996 52444
rect 20044 52388 20100 52444
rect 50556 52388 50612 52444
rect 50660 52388 50716 52444
rect 50764 52388 50820 52444
rect 4476 51380 4532 51436
rect 4580 51380 4636 51436
rect 4684 51380 4740 51436
rect 35196 51380 35252 51436
rect 35300 51380 35356 51436
rect 35404 51380 35460 51436
rect 19836 50372 19892 50428
rect 19940 50372 19996 50428
rect 20044 50372 20100 50428
rect 50556 50372 50612 50428
rect 50660 50372 50716 50428
rect 50764 50372 50820 50428
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48356 19892 48412
rect 19940 48356 19996 48412
rect 20044 48356 20100 48412
rect 50556 48356 50612 48412
rect 50660 48356 50716 48412
rect 50764 48356 50820 48412
rect 4476 47348 4532 47404
rect 4580 47348 4636 47404
rect 4684 47348 4740 47404
rect 35196 47348 35252 47404
rect 35300 47348 35356 47404
rect 35404 47348 35460 47404
rect 19836 46340 19892 46396
rect 19940 46340 19996 46396
rect 20044 46340 20100 46396
rect 50556 46340 50612 46396
rect 50660 46340 50716 46396
rect 50764 46340 50820 46396
rect 4476 45332 4532 45388
rect 4580 45332 4636 45388
rect 4684 45332 4740 45388
rect 35196 45332 35252 45388
rect 35300 45332 35356 45388
rect 35404 45332 35460 45388
rect 19836 44324 19892 44380
rect 19940 44324 19996 44380
rect 20044 44324 20100 44380
rect 50556 44324 50612 44380
rect 50660 44324 50716 44380
rect 50764 44324 50820 44380
rect 23548 43820 23604 43876
rect 4476 43316 4532 43372
rect 4580 43316 4636 43372
rect 4684 43316 4740 43372
rect 35196 43316 35252 43372
rect 35300 43316 35356 43372
rect 35404 43316 35460 43372
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 23548 41916 23604 41972
rect 4476 41300 4532 41356
rect 4580 41300 4636 41356
rect 4684 41300 4740 41356
rect 35196 41300 35252 41356
rect 35300 41300 35356 41356
rect 35404 41300 35460 41356
rect 19836 40292 19892 40348
rect 19940 40292 19996 40348
rect 20044 40292 20100 40348
rect 50556 40292 50612 40348
rect 50660 40292 50716 40348
rect 50764 40292 50820 40348
rect 4476 39284 4532 39340
rect 4580 39284 4636 39340
rect 4684 39284 4740 39340
rect 35196 39284 35252 39340
rect 35300 39284 35356 39340
rect 35404 39284 35460 39340
rect 19836 38276 19892 38332
rect 19940 38276 19996 38332
rect 20044 38276 20100 38332
rect 50556 38276 50612 38332
rect 50660 38276 50716 38332
rect 50764 38276 50820 38332
rect 4476 37268 4532 37324
rect 4580 37268 4636 37324
rect 4684 37268 4740 37324
rect 35196 37268 35252 37324
rect 35300 37268 35356 37324
rect 35404 37268 35460 37324
rect 19836 36260 19892 36316
rect 19940 36260 19996 36316
rect 20044 36260 20100 36316
rect 50556 36260 50612 36316
rect 50660 36260 50716 36316
rect 50764 36260 50820 36316
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34244 19892 34300
rect 19940 34244 19996 34300
rect 20044 34244 20100 34300
rect 50556 34244 50612 34300
rect 50660 34244 50716 34300
rect 50764 34244 50820 34300
rect 25788 33292 25844 33348
rect 4476 33236 4532 33292
rect 4580 33236 4636 33292
rect 4684 33236 4740 33292
rect 35196 33236 35252 33292
rect 35300 33236 35356 33292
rect 35404 33236 35460 33292
rect 19836 32228 19892 32284
rect 19940 32228 19996 32284
rect 20044 32228 20100 32284
rect 50556 32228 50612 32284
rect 50660 32228 50716 32284
rect 50764 32228 50820 32284
rect 26460 31836 26516 31892
rect 25788 31612 25844 31668
rect 4476 31220 4532 31276
rect 4580 31220 4636 31276
rect 4684 31220 4740 31276
rect 35196 31220 35252 31276
rect 35300 31220 35356 31276
rect 35404 31220 35460 31276
rect 38220 30604 38276 30660
rect 38220 30268 38276 30324
rect 19836 30212 19892 30268
rect 19940 30212 19996 30268
rect 20044 30212 20100 30268
rect 50556 30212 50612 30268
rect 50660 30212 50716 30268
rect 50764 30212 50820 30268
rect 4476 29204 4532 29260
rect 4580 29204 4636 29260
rect 4684 29204 4740 29260
rect 35196 29204 35252 29260
rect 35300 29204 35356 29260
rect 35404 29204 35460 29260
rect 26460 28364 26516 28420
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27188 4532 27244
rect 4580 27188 4636 27244
rect 4684 27188 4740 27244
rect 35196 27188 35252 27244
rect 35300 27188 35356 27244
rect 35404 27188 35460 27244
rect 33628 27132 33684 27188
rect 19836 26180 19892 26236
rect 19940 26180 19996 26236
rect 20044 26180 20100 26236
rect 50556 26180 50612 26236
rect 50660 26180 50716 26236
rect 50764 26180 50820 26236
rect 4476 25172 4532 25228
rect 4580 25172 4636 25228
rect 4684 25172 4740 25228
rect 35196 25172 35252 25228
rect 35300 25172 35356 25228
rect 35404 25172 35460 25228
rect 33628 24332 33684 24388
rect 19836 24164 19892 24220
rect 19940 24164 19996 24220
rect 20044 24164 20100 24220
rect 50556 24164 50612 24220
rect 50660 24164 50716 24220
rect 50764 24164 50820 24220
rect 4476 23156 4532 23212
rect 4580 23156 4636 23212
rect 4684 23156 4740 23212
rect 35196 23156 35252 23212
rect 35300 23156 35356 23212
rect 35404 23156 35460 23212
rect 19836 22148 19892 22204
rect 19940 22148 19996 22204
rect 20044 22148 20100 22204
rect 50556 22148 50612 22204
rect 50660 22148 50716 22204
rect 50764 22148 50820 22204
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20132 19892 20188
rect 19940 20132 19996 20188
rect 20044 20132 20100 20188
rect 27468 20188 27524 20244
rect 50556 20132 50612 20188
rect 50660 20132 50716 20188
rect 50764 20132 50820 20188
rect 4476 19124 4532 19180
rect 4580 19124 4636 19180
rect 4684 19124 4740 19180
rect 35196 19124 35252 19180
rect 35300 19124 35356 19180
rect 35404 19124 35460 19180
rect 19836 18116 19892 18172
rect 19940 18116 19996 18172
rect 20044 18116 20100 18172
rect 50556 18116 50612 18172
rect 50660 18116 50716 18172
rect 50764 18116 50820 18172
rect 4476 17108 4532 17164
rect 4580 17108 4636 17164
rect 4684 17108 4740 17164
rect 35196 17108 35252 17164
rect 35300 17108 35356 17164
rect 35404 17108 35460 17164
rect 19836 16100 19892 16156
rect 19940 16100 19996 16156
rect 20044 16100 20100 16156
rect 50556 16100 50612 16156
rect 50660 16100 50716 16156
rect 50764 16100 50820 16156
rect 27468 15148 27524 15204
rect 4476 15092 4532 15148
rect 4580 15092 4636 15148
rect 4684 15092 4740 15148
rect 35196 15092 35252 15148
rect 35300 15092 35356 15148
rect 35404 15092 35460 15148
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13076 4532 13132
rect 4580 13076 4636 13132
rect 4684 13076 4740 13132
rect 35196 13076 35252 13132
rect 35300 13076 35356 13132
rect 35404 13076 35460 13132
rect 19836 12068 19892 12124
rect 19940 12068 19996 12124
rect 20044 12068 20100 12124
rect 50556 12068 50612 12124
rect 50660 12068 50716 12124
rect 50764 12068 50820 12124
rect 4476 11060 4532 11116
rect 4580 11060 4636 11116
rect 4684 11060 4740 11116
rect 35196 11060 35252 11116
rect 35300 11060 35356 11116
rect 35404 11060 35460 11116
rect 19836 10052 19892 10108
rect 19940 10052 19996 10108
rect 20044 10052 20100 10108
rect 50556 10052 50612 10108
rect 50660 10052 50716 10108
rect 50764 10052 50820 10108
rect 4476 9044 4532 9100
rect 4580 9044 4636 9100
rect 4684 9044 4740 9100
rect 35196 9044 35252 9100
rect 35300 9044 35356 9100
rect 35404 9044 35460 9100
rect 19836 8036 19892 8092
rect 19940 8036 19996 8092
rect 20044 8036 20100 8092
rect 50556 8036 50612 8092
rect 50660 8036 50716 8092
rect 50764 8036 50820 8092
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6020 19892 6076
rect 19940 6020 19996 6076
rect 20044 6020 20100 6076
rect 50556 6020 50612 6076
rect 50660 6020 50716 6076
rect 50764 6020 50820 6076
rect 4476 5012 4532 5068
rect 4580 5012 4636 5068
rect 4684 5012 4740 5068
rect 35196 5012 35252 5068
rect 35300 5012 35356 5068
rect 35404 5012 35460 5068
rect 19836 4004 19892 4060
rect 19940 4004 19996 4060
rect 20044 4004 20100 4060
rect 50556 4004 50612 4060
rect 50660 4004 50716 4060
rect 50764 4004 50820 4060
<< metal4 >>
rect 4448 55468 4768 56508
rect 4448 55412 4476 55468
rect 4532 55412 4580 55468
rect 4636 55412 4684 55468
rect 4740 55412 4768 55468
rect 4448 53452 4768 55412
rect 4448 53396 4476 53452
rect 4532 53396 4580 53452
rect 4636 53396 4684 53452
rect 4740 53396 4768 53452
rect 4448 51436 4768 53396
rect 4448 51380 4476 51436
rect 4532 51380 4580 51436
rect 4636 51380 4684 51436
rect 4740 51380 4768 51436
rect 4448 49420 4768 51380
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47404 4768 49364
rect 4448 47348 4476 47404
rect 4532 47348 4580 47404
rect 4636 47348 4684 47404
rect 4740 47348 4768 47404
rect 4448 45388 4768 47348
rect 4448 45332 4476 45388
rect 4532 45332 4580 45388
rect 4636 45332 4684 45388
rect 4740 45332 4768 45388
rect 4448 43372 4768 45332
rect 4448 43316 4476 43372
rect 4532 43316 4580 43372
rect 4636 43316 4684 43372
rect 4740 43316 4768 43372
rect 4448 41356 4768 43316
rect 4448 41300 4476 41356
rect 4532 41300 4580 41356
rect 4636 41300 4684 41356
rect 4740 41300 4768 41356
rect 4448 39340 4768 41300
rect 4448 39284 4476 39340
rect 4532 39284 4580 39340
rect 4636 39284 4684 39340
rect 4740 39284 4768 39340
rect 4448 37324 4768 39284
rect 4448 37268 4476 37324
rect 4532 37268 4580 37324
rect 4636 37268 4684 37324
rect 4740 37268 4768 37324
rect 4448 35308 4768 37268
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33292 4768 35252
rect 4448 33236 4476 33292
rect 4532 33236 4580 33292
rect 4636 33236 4684 33292
rect 4740 33236 4768 33292
rect 4448 31276 4768 33236
rect 4448 31220 4476 31276
rect 4532 31220 4580 31276
rect 4636 31220 4684 31276
rect 4740 31220 4768 31276
rect 4448 29260 4768 31220
rect 4448 29204 4476 29260
rect 4532 29204 4580 29260
rect 4636 29204 4684 29260
rect 4740 29204 4768 29260
rect 4448 27244 4768 29204
rect 4448 27188 4476 27244
rect 4532 27188 4580 27244
rect 4636 27188 4684 27244
rect 4740 27188 4768 27244
rect 4448 25228 4768 27188
rect 4448 25172 4476 25228
rect 4532 25172 4580 25228
rect 4636 25172 4684 25228
rect 4740 25172 4768 25228
rect 4448 23212 4768 25172
rect 4448 23156 4476 23212
rect 4532 23156 4580 23212
rect 4636 23156 4684 23212
rect 4740 23156 4768 23212
rect 4448 21196 4768 23156
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19180 4768 21140
rect 4448 19124 4476 19180
rect 4532 19124 4580 19180
rect 4636 19124 4684 19180
rect 4740 19124 4768 19180
rect 4448 17164 4768 19124
rect 4448 17108 4476 17164
rect 4532 17108 4580 17164
rect 4636 17108 4684 17164
rect 4740 17108 4768 17164
rect 4448 15148 4768 17108
rect 4448 15092 4476 15148
rect 4532 15092 4580 15148
rect 4636 15092 4684 15148
rect 4740 15092 4768 15148
rect 4448 13132 4768 15092
rect 4448 13076 4476 13132
rect 4532 13076 4580 13132
rect 4636 13076 4684 13132
rect 4740 13076 4768 13132
rect 4448 11116 4768 13076
rect 4448 11060 4476 11116
rect 4532 11060 4580 11116
rect 4636 11060 4684 11116
rect 4740 11060 4768 11116
rect 4448 9100 4768 11060
rect 4448 9044 4476 9100
rect 4532 9044 4580 9100
rect 4636 9044 4684 9100
rect 4740 9044 4768 9100
rect 4448 7084 4768 9044
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5068 4768 7028
rect 4448 5012 4476 5068
rect 4532 5012 4580 5068
rect 4636 5012 4684 5068
rect 4740 5012 4768 5068
rect 4448 3972 4768 5012
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54460 20128 56420
rect 19808 54404 19836 54460
rect 19892 54404 19940 54460
rect 19996 54404 20044 54460
rect 20100 54404 20128 54460
rect 19808 52444 20128 54404
rect 19808 52388 19836 52444
rect 19892 52388 19940 52444
rect 19996 52388 20044 52444
rect 20100 52388 20128 52444
rect 19808 50428 20128 52388
rect 19808 50372 19836 50428
rect 19892 50372 19940 50428
rect 19996 50372 20044 50428
rect 20100 50372 20128 50428
rect 19808 48412 20128 50372
rect 19808 48356 19836 48412
rect 19892 48356 19940 48412
rect 19996 48356 20044 48412
rect 20100 48356 20128 48412
rect 19808 46396 20128 48356
rect 19808 46340 19836 46396
rect 19892 46340 19940 46396
rect 19996 46340 20044 46396
rect 20100 46340 20128 46396
rect 19808 44380 20128 46340
rect 19808 44324 19836 44380
rect 19892 44324 19940 44380
rect 19996 44324 20044 44380
rect 20100 44324 20128 44380
rect 19808 42364 20128 44324
rect 35168 55468 35488 56508
rect 35168 55412 35196 55468
rect 35252 55412 35300 55468
rect 35356 55412 35404 55468
rect 35460 55412 35488 55468
rect 35168 53452 35488 55412
rect 35168 53396 35196 53452
rect 35252 53396 35300 53452
rect 35356 53396 35404 53452
rect 35460 53396 35488 53452
rect 35168 51436 35488 53396
rect 35168 51380 35196 51436
rect 35252 51380 35300 51436
rect 35356 51380 35404 51436
rect 35460 51380 35488 51436
rect 35168 49420 35488 51380
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47404 35488 49364
rect 35168 47348 35196 47404
rect 35252 47348 35300 47404
rect 35356 47348 35404 47404
rect 35460 47348 35488 47404
rect 35168 45388 35488 47348
rect 35168 45332 35196 45388
rect 35252 45332 35300 45388
rect 35356 45332 35404 45388
rect 35460 45332 35488 45388
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40348 20128 42308
rect 23548 43876 23604 43886
rect 23548 41972 23604 43820
rect 23548 41906 23604 41916
rect 35168 43372 35488 45332
rect 35168 43316 35196 43372
rect 35252 43316 35300 43372
rect 35356 43316 35404 43372
rect 35460 43316 35488 43372
rect 19808 40292 19836 40348
rect 19892 40292 19940 40348
rect 19996 40292 20044 40348
rect 20100 40292 20128 40348
rect 19808 38332 20128 40292
rect 19808 38276 19836 38332
rect 19892 38276 19940 38332
rect 19996 38276 20044 38332
rect 20100 38276 20128 38332
rect 19808 36316 20128 38276
rect 19808 36260 19836 36316
rect 19892 36260 19940 36316
rect 19996 36260 20044 36316
rect 20100 36260 20128 36316
rect 19808 34300 20128 36260
rect 19808 34244 19836 34300
rect 19892 34244 19940 34300
rect 19996 34244 20044 34300
rect 20100 34244 20128 34300
rect 19808 32284 20128 34244
rect 35168 41356 35488 43316
rect 35168 41300 35196 41356
rect 35252 41300 35300 41356
rect 35356 41300 35404 41356
rect 35460 41300 35488 41356
rect 35168 39340 35488 41300
rect 35168 39284 35196 39340
rect 35252 39284 35300 39340
rect 35356 39284 35404 39340
rect 35460 39284 35488 39340
rect 35168 37324 35488 39284
rect 35168 37268 35196 37324
rect 35252 37268 35300 37324
rect 35356 37268 35404 37324
rect 35460 37268 35488 37324
rect 35168 35308 35488 37268
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 19808 32228 19836 32284
rect 19892 32228 19940 32284
rect 19996 32228 20044 32284
rect 20100 32228 20128 32284
rect 19808 30268 20128 32228
rect 25788 33348 25844 33358
rect 25788 31668 25844 33292
rect 35168 33292 35488 35252
rect 35168 33236 35196 33292
rect 35252 33236 35300 33292
rect 35356 33236 35404 33292
rect 35460 33236 35488 33292
rect 25788 31602 25844 31612
rect 26460 31892 26516 31902
rect 19808 30212 19836 30268
rect 19892 30212 19940 30268
rect 19996 30212 20044 30268
rect 20100 30212 20128 30268
rect 19808 28252 20128 30212
rect 26460 28420 26516 31836
rect 26460 28354 26516 28364
rect 35168 31276 35488 33236
rect 35168 31220 35196 31276
rect 35252 31220 35300 31276
rect 35356 31220 35404 31276
rect 35460 31220 35488 31276
rect 35168 29260 35488 31220
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54460 50848 56420
rect 50528 54404 50556 54460
rect 50612 54404 50660 54460
rect 50716 54404 50764 54460
rect 50820 54404 50848 54460
rect 50528 52444 50848 54404
rect 50528 52388 50556 52444
rect 50612 52388 50660 52444
rect 50716 52388 50764 52444
rect 50820 52388 50848 52444
rect 50528 50428 50848 52388
rect 50528 50372 50556 50428
rect 50612 50372 50660 50428
rect 50716 50372 50764 50428
rect 50820 50372 50848 50428
rect 50528 48412 50848 50372
rect 50528 48356 50556 48412
rect 50612 48356 50660 48412
rect 50716 48356 50764 48412
rect 50820 48356 50848 48412
rect 50528 46396 50848 48356
rect 50528 46340 50556 46396
rect 50612 46340 50660 46396
rect 50716 46340 50764 46396
rect 50820 46340 50848 46396
rect 50528 44380 50848 46340
rect 50528 44324 50556 44380
rect 50612 44324 50660 44380
rect 50716 44324 50764 44380
rect 50820 44324 50848 44380
rect 50528 42364 50848 44324
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40348 50848 42308
rect 50528 40292 50556 40348
rect 50612 40292 50660 40348
rect 50716 40292 50764 40348
rect 50820 40292 50848 40348
rect 50528 38332 50848 40292
rect 50528 38276 50556 38332
rect 50612 38276 50660 38332
rect 50716 38276 50764 38332
rect 50820 38276 50848 38332
rect 50528 36316 50848 38276
rect 50528 36260 50556 36316
rect 50612 36260 50660 36316
rect 50716 36260 50764 36316
rect 50820 36260 50848 36316
rect 50528 34300 50848 36260
rect 50528 34244 50556 34300
rect 50612 34244 50660 34300
rect 50716 34244 50764 34300
rect 50820 34244 50848 34300
rect 50528 32284 50848 34244
rect 50528 32228 50556 32284
rect 50612 32228 50660 32284
rect 50716 32228 50764 32284
rect 50820 32228 50848 32284
rect 38220 30660 38276 30670
rect 38220 30324 38276 30604
rect 38220 30258 38276 30268
rect 50528 30268 50848 32228
rect 35168 29204 35196 29260
rect 35252 29204 35300 29260
rect 35356 29204 35404 29260
rect 35460 29204 35488 29260
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26236 20128 28196
rect 35168 27244 35488 29204
rect 19808 26180 19836 26236
rect 19892 26180 19940 26236
rect 19996 26180 20044 26236
rect 20100 26180 20128 26236
rect 19808 24220 20128 26180
rect 33628 27188 33684 27198
rect 33628 24388 33684 27132
rect 33628 24322 33684 24332
rect 35168 27188 35196 27244
rect 35252 27188 35300 27244
rect 35356 27188 35404 27244
rect 35460 27188 35488 27244
rect 35168 25228 35488 27188
rect 35168 25172 35196 25228
rect 35252 25172 35300 25228
rect 35356 25172 35404 25228
rect 35460 25172 35488 25228
rect 19808 24164 19836 24220
rect 19892 24164 19940 24220
rect 19996 24164 20044 24220
rect 20100 24164 20128 24220
rect 19808 22204 20128 24164
rect 19808 22148 19836 22204
rect 19892 22148 19940 22204
rect 19996 22148 20044 22204
rect 20100 22148 20128 22204
rect 19808 20188 20128 22148
rect 35168 23212 35488 25172
rect 35168 23156 35196 23212
rect 35252 23156 35300 23212
rect 35356 23156 35404 23212
rect 35460 23156 35488 23212
rect 35168 21196 35488 23156
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 19808 20132 19836 20188
rect 19892 20132 19940 20188
rect 19996 20132 20044 20188
rect 20100 20132 20128 20188
rect 19808 18172 20128 20132
rect 19808 18116 19836 18172
rect 19892 18116 19940 18172
rect 19996 18116 20044 18172
rect 20100 18116 20128 18172
rect 19808 16156 20128 18116
rect 19808 16100 19836 16156
rect 19892 16100 19940 16156
rect 19996 16100 20044 16156
rect 20100 16100 20128 16156
rect 19808 14140 20128 16100
rect 27468 20244 27524 20254
rect 27468 15204 27524 20188
rect 27468 15138 27524 15148
rect 35168 19180 35488 21140
rect 35168 19124 35196 19180
rect 35252 19124 35300 19180
rect 35356 19124 35404 19180
rect 35460 19124 35488 19180
rect 35168 17164 35488 19124
rect 35168 17108 35196 17164
rect 35252 17108 35300 17164
rect 35356 17108 35404 17164
rect 35460 17108 35488 17164
rect 35168 15148 35488 17108
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12124 20128 14084
rect 19808 12068 19836 12124
rect 19892 12068 19940 12124
rect 19996 12068 20044 12124
rect 20100 12068 20128 12124
rect 19808 10108 20128 12068
rect 19808 10052 19836 10108
rect 19892 10052 19940 10108
rect 19996 10052 20044 10108
rect 20100 10052 20128 10108
rect 19808 8092 20128 10052
rect 19808 8036 19836 8092
rect 19892 8036 19940 8092
rect 19996 8036 20044 8092
rect 20100 8036 20128 8092
rect 19808 6076 20128 8036
rect 19808 6020 19836 6076
rect 19892 6020 19940 6076
rect 19996 6020 20044 6076
rect 20100 6020 20128 6076
rect 19808 4060 20128 6020
rect 19808 4004 19836 4060
rect 19892 4004 19940 4060
rect 19996 4004 20044 4060
rect 20100 4004 20128 4060
rect 19808 3972 20128 4004
rect 35168 15092 35196 15148
rect 35252 15092 35300 15148
rect 35356 15092 35404 15148
rect 35460 15092 35488 15148
rect 35168 13132 35488 15092
rect 35168 13076 35196 13132
rect 35252 13076 35300 13132
rect 35356 13076 35404 13132
rect 35460 13076 35488 13132
rect 35168 11116 35488 13076
rect 35168 11060 35196 11116
rect 35252 11060 35300 11116
rect 35356 11060 35404 11116
rect 35460 11060 35488 11116
rect 35168 9100 35488 11060
rect 35168 9044 35196 9100
rect 35252 9044 35300 9100
rect 35356 9044 35404 9100
rect 35460 9044 35488 9100
rect 35168 7084 35488 9044
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5068 35488 7028
rect 35168 5012 35196 5068
rect 35252 5012 35300 5068
rect 35356 5012 35404 5068
rect 35460 5012 35488 5068
rect 35168 3972 35488 5012
rect 50528 30212 50556 30268
rect 50612 30212 50660 30268
rect 50716 30212 50764 30268
rect 50820 30212 50848 30268
rect 50528 28252 50848 30212
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26236 50848 28196
rect 50528 26180 50556 26236
rect 50612 26180 50660 26236
rect 50716 26180 50764 26236
rect 50820 26180 50848 26236
rect 50528 24220 50848 26180
rect 50528 24164 50556 24220
rect 50612 24164 50660 24220
rect 50716 24164 50764 24220
rect 50820 24164 50848 24220
rect 50528 22204 50848 24164
rect 50528 22148 50556 22204
rect 50612 22148 50660 22204
rect 50716 22148 50764 22204
rect 50820 22148 50848 22204
rect 50528 20188 50848 22148
rect 50528 20132 50556 20188
rect 50612 20132 50660 20188
rect 50716 20132 50764 20188
rect 50820 20132 50848 20188
rect 50528 18172 50848 20132
rect 50528 18116 50556 18172
rect 50612 18116 50660 18172
rect 50716 18116 50764 18172
rect 50820 18116 50848 18172
rect 50528 16156 50848 18116
rect 50528 16100 50556 16156
rect 50612 16100 50660 16156
rect 50716 16100 50764 16156
rect 50820 16100 50848 16156
rect 50528 14140 50848 16100
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12124 50848 14084
rect 50528 12068 50556 12124
rect 50612 12068 50660 12124
rect 50716 12068 50764 12124
rect 50820 12068 50848 12124
rect 50528 10108 50848 12068
rect 50528 10052 50556 10108
rect 50612 10052 50660 10108
rect 50716 10052 50764 10108
rect 50820 10052 50848 10108
rect 50528 8092 50848 10052
rect 50528 8036 50556 8092
rect 50612 8036 50660 8092
rect 50716 8036 50764 8092
rect 50820 8036 50848 8092
rect 50528 6076 50848 8036
rect 50528 6020 50556 6076
rect 50612 6020 50660 6076
rect 50716 6020 50764 6076
rect 50820 6020 50848 6076
rect 50528 4060 50848 6020
rect 50528 4004 50556 4060
rect 50612 4004 50660 4060
rect 50716 4004 50764 4060
rect 50820 4004 50848 4060
rect 50528 3972 50848 4004
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _244_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 14560 0 -1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _245_
timestamp 1698431365
transform 1 0 27328 0 -1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _246_
timestamp 1698431365
transform -1 0 27328 0 1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _247_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 35168 0 -1 36288
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _248_
timestamp 1698431365
transform 1 0 35728 0 -1 22176
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _249_
timestamp 1698431365
transform -1 0 34944 0 -1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _250_
timestamp 1698431365
transform 1 0 34720 0 -1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _251_
timestamp 1698431365
transform -1 0 28784 0 1 16128
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _252_
timestamp 1698431365
transform -1 0 27776 0 1 16128
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _253_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 31024 0 -1 18144
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _254_
timestamp 1698431365
transform -1 0 34608 0 -1 22176
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _255_
timestamp 1698431365
transform -1 0 27104 0 1 14112
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _256_
timestamp 1698431365
transform -1 0 22512 0 -1 14112
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _257_
timestamp 1698431365
transform 1 0 23296 0 1 16128
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _258_
timestamp 1698431365
transform 1 0 19600 0 -1 18144
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _259_
timestamp 1698431365
transform 1 0 18816 0 -1 16128
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _260_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _261_
timestamp 1698431365
transform -1 0 33600 0 -1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _262_
timestamp 1698431365
transform 1 0 26208 0 1 18144
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _263_
timestamp 1698431365
transform 1 0 30576 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _264_
timestamp 1698431365
transform 1 0 34272 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _265_
timestamp 1698431365
transform -1 0 34720 0 -1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _266_
timestamp 1698431365
transform 1 0 22736 0 1 18144
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _267_
timestamp 1698431365
transform -1 0 32704 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _268_
timestamp 1698431365
transform -1 0 32368 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _269_
timestamp 1698431365
transform -1 0 28000 0 1 22176
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _270_
timestamp 1698431365
transform -1 0 25760 0 -1 26208
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  _271_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 24640 0 1 26208
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _272_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 22624 0 1 20160
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _273_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 1 24192
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _274_
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _275_
timestamp 1698431365
transform -1 0 30688 0 -1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _276_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 31136 0 1 28224
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _277_
timestamp 1698431365
transform 1 0 22624 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _278_
timestamp 1698431365
transform 1 0 21392 0 -1 6048
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _279_
timestamp 1698431365
transform 1 0 21168 0 1 10080
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _280_
timestamp 1698431365
transform 1 0 23072 0 -1 12096
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _281_
timestamp 1698431365
transform 1 0 23408 0 1 26208
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _282_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 24864 0 -1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _283_
timestamp 1698431365
transform 1 0 22624 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _284_
timestamp 1698431365
transform -1 0 24416 0 1 30240
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _285_
timestamp 1698431365
transform 1 0 14000 0 -1 34272
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _286_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 16576 0 -1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _287_
timestamp 1698431365
transform 1 0 25088 0 -1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _288_
timestamp 1698431365
transform 1 0 27440 0 -1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _289_
timestamp 1698431365
transform -1 0 36848 0 -1 38304
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _290_
timestamp 1698431365
transform 1 0 43904 0 -1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _291_
timestamp 1698431365
transform 1 0 40768 0 -1 38304
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _292_
timestamp 1698431365
transform 1 0 37520 0 1 36288
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _293_
timestamp 1698431365
transform 1 0 47040 0 -1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _294_
timestamp 1698431365
transform 1 0 50064 0 -1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _295_
timestamp 1698431365
transform 1 0 52640 0 -1 42336
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _296_
timestamp 1698431365
transform 1 0 46144 0 -1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _297_
timestamp 1698431365
transform 1 0 46256 0 1 38304
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _298_
timestamp 1698431365
transform 1 0 44912 0 -1 40320
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _299_
timestamp 1698431365
transform 1 0 49392 0 -1 40320
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _300_
timestamp 1698431365
transform 1 0 46368 0 -1 38304
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _301_
timestamp 1698431365
transform 1 0 45024 0 1 36288
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  _302_
timestamp 1698431365
transform -1 0 28000 0 1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _303_
timestamp 1698431365
transform -1 0 32256 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _304_
timestamp 1698431365
transform -1 0 27216 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _305_
timestamp 1698431365
transform 1 0 25760 0 -1 10080
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _306_
timestamp 1698431365
transform 1 0 33040 0 1 14112
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _307_
timestamp 1698431365
transform 1 0 34608 0 1 18144
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _308_
timestamp 1698431365
transform 1 0 32928 0 -1 8064
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _309_
timestamp 1698431365
transform -1 0 27888 0 1 10080
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _310_
timestamp 1698431365
transform -1 0 34272 0 -1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _311_
timestamp 1698431365
transform 1 0 36064 0 -1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _312_
timestamp 1698431365
transform 1 0 37520 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _313_
timestamp 1698431365
transform -1 0 36176 0 1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _314_
timestamp 1698431365
transform -1 0 32816 0 1 22176
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__nand3_1  _315_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29232 0 1 24192
box -86 -90 870 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _316_
timestamp 1698431365
transform 1 0 40768 0 -1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _317_
timestamp 1698431365
transform 1 0 42224 0 1 26208
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _318_
timestamp 1698431365
transform -1 0 31024 0 -1 26208
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_1  _319_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 30464 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _320_
timestamp 1698431365
transform 1 0 25088 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _321_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 26432 0 1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__nor3_1  _322_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 24416 0 1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _323_
timestamp 1698431365
transform 1 0 14896 0 -1 32256
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _324_
timestamp 1698431365
transform 1 0 32928 0 -1 12096
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _325_
timestamp 1698431365
transform -1 0 43232 0 -1 22176
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _326_
timestamp 1698431365
transform 1 0 40768 0 -1 10080
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _327_
timestamp 1698431365
transform 1 0 31920 0 1 12096
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _328_
timestamp 1698431365
transform 1 0 31248 0 -1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  _329_
timestamp 1698431365
transform -1 0 26544 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _330_
timestamp 1698431365
transform -1 0 26656 0 -1 22176
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _331_
timestamp 1698431365
transform -1 0 23296 0 -1 26208
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _332_
timestamp 1698431365
transform 1 0 15904 0 1 26208
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _333_
timestamp 1698431365
transform 1 0 24640 0 1 26208
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  _334_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 32480 0 -1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _335_
timestamp 1698431365
transform 1 0 34048 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _336_
timestamp 1698431365
transform -1 0 31136 0 1 24192
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _337_
timestamp 1698431365
transform -1 0 27328 0 -1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _338_
timestamp 1698431365
transform 1 0 23408 0 -1 26208
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _339_
timestamp 1698431365
transform 1 0 26656 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _340_
timestamp 1698431365
transform 1 0 32368 0 1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _341_
timestamp 1698431365
transform -1 0 32704 0 -1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _342_
timestamp 1698431365
transform 1 0 36848 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _343_
timestamp 1698431365
transform 1 0 38192 0 1 36288
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _344_
timestamp 1698431365
transform -1 0 32368 0 1 32256
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _345_
timestamp 1698431365
transform 1 0 29792 0 1 26208
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  _346_
timestamp 1698431365
transform 1 0 35840 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _347_
timestamp 1698431365
transform 1 0 33488 0 1 26208
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _348_
timestamp 1698431365
transform -1 0 36624 0 -1 40320
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _349_
timestamp 1698431365
transform 1 0 33040 0 1 32256
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _350_
timestamp 1698431365
transform -1 0 32704 0 -1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _351_
timestamp 1698431365
transform 1 0 33376 0 1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _352_
timestamp 1698431365
transform -1 0 49056 0 1 26208
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _353_
timestamp 1698431365
transform 1 0 37072 0 -1 24192
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _354_
timestamp 1698431365
transform -1 0 36064 0 -1 28224
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _355_
timestamp 1698431365
transform 1 0 33824 0 1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_1  _356_
timestamp 1698431365
transform -1 0 31136 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _357_
timestamp 1698431365
transform 1 0 22400 0 -1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _358_
timestamp 1698431365
transform 1 0 26208 0 -1 30240
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _359_
timestamp 1698431365
transform 1 0 15008 0 1 30240
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _360_
timestamp 1698431365
transform 1 0 36624 0 -1 16128
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _361_
timestamp 1698431365
transform 1 0 38752 0 1 38304
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _362_
timestamp 1698431365
transform 1 0 40432 0 1 18144
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _363_
timestamp 1698431365
transform 1 0 38640 0 1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _364_
timestamp 1698431365
transform 1 0 35168 0 1 20160
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _365_
timestamp 1698431365
transform -1 0 18704 0 -1 26208
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _366_
timestamp 1698431365
transform 1 0 25648 0 1 26208
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _367_
timestamp 1698431365
transform 1 0 48608 0 -1 36288
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _368_
timestamp 1698431365
transform 1 0 49728 0 -1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _369_
timestamp 1698431365
transform 1 0 49280 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _370_
timestamp 1698431365
transform 1 0 52752 0 1 32256
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _371_
timestamp 1698431365
transform -1 0 50848 0 1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _372_
timestamp 1698431365
transform 1 0 52864 0 1 36288
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _373_
timestamp 1698431365
transform 1 0 52080 0 -1 34272
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _374_
timestamp 1698431365
transform 1 0 50848 0 1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _375_
timestamp 1698431365
transform 1 0 48608 0 -1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  _376_
timestamp 1698431365
transform -1 0 27440 0 -1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _377_
timestamp 1698431365
transform -1 0 26208 0 -1 30240
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _378_
timestamp 1698431365
transform 1 0 14000 0 1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _379_
timestamp 1698431365
transform 1 0 13552 0 1 30240
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _380_
timestamp 1698431365
transform 1 0 41552 0 -1 14112
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _381_
timestamp 1698431365
transform -1 0 38080 0 -1 40320
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _382_
timestamp 1698431365
transform -1 0 43120 0 1 40320
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _383_
timestamp 1698431365
transform 1 0 40768 0 -1 44352
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _384_
timestamp 1698431365
transform 1 0 40096 0 1 28224
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _385_
timestamp 1698431365
transform -1 0 22624 0 1 26208
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  _386_
timestamp 1698431365
transform -1 0 25760 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _387_
timestamp 1698431365
transform 1 0 24304 0 1 28224
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  _388_
timestamp 1698431365
transform -1 0 33264 0 1 20160
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _389_
timestamp 1698431365
transform 1 0 31136 0 1 24192
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _390_
timestamp 1698431365
transform 1 0 25872 0 1 22176
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _391_
timestamp 1698431365
transform 1 0 26320 0 1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _392_
timestamp 1698431365
transform 1 0 42672 0 -1 34272
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _393_
timestamp 1698431365
transform -1 0 32032 0 -1 32256
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _394_
timestamp 1698431365
transform 1 0 30576 0 -1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  _395_
timestamp 1698431365
transform 1 0 33040 0 -1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _396_
timestamp 1698431365
transform -1 0 35728 0 1 26208
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _397_
timestamp 1698431365
transform 1 0 33040 0 -1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _398_
timestamp 1698431365
transform -1 0 33376 0 1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _399_
timestamp 1698431365
transform 1 0 38304 0 1 26208
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _400_
timestamp 1698431365
transform -1 0 35504 0 -1 28224
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _401_
timestamp 1698431365
transform 1 0 32704 0 1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_1  _402_
timestamp 1698431365
transform -1 0 30240 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _403_
timestamp 1698431365
transform -1 0 24864 0 -1 30240
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _404_
timestamp 1698431365
transform 1 0 14000 0 1 28224
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _405_
timestamp 1698431365
transform -1 0 28672 0 -1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _406_
timestamp 1698431365
transform 1 0 40768 0 -1 40320
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _407_
timestamp 1698431365
transform 1 0 31584 0 1 42336
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _408_
timestamp 1698431365
transform 1 0 34496 0 -1 40320
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _409_
timestamp 1698431365
transform 1 0 26096 0 1 38304
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _410_
timestamp 1698431365
transform 1 0 25088 0 -1 38304
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _411_
timestamp 1698431365
transform 1 0 51184 0 -1 30240
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _412_
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _413_
timestamp 1698431365
transform 1 0 49952 0 1 26208
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _414_
timestamp 1698431365
transform 1 0 51968 0 -1 28224
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _415_
timestamp 1698431365
transform 1 0 46480 0 -1 28224
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _416_
timestamp 1698431365
transform 1 0 50848 0 1 28224
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _417_
timestamp 1698431365
transform 1 0 52976 0 1 24192
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _418_
timestamp 1698431365
transform 1 0 49280 0 -1 22176
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _419_
timestamp 1698431365
transform 1 0 50176 0 1 24192
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _420_
timestamp 1698431365
transform 1 0 48608 0 -1 30240
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  _421_
timestamp 1698431365
transform -1 0 28784 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _422_
timestamp 1698431365
transform 1 0 25536 0 -1 32256
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _423_
timestamp 1698431365
transform 1 0 14224 0 -1 30240
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _424_
timestamp 1698431365
transform 1 0 41216 0 -1 16128
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _425_
timestamp 1698431365
transform 1 0 39536 0 1 42336
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _426_
timestamp 1698431365
transform 1 0 40768 0 -1 30240
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _427_
timestamp 1698431365
transform -1 0 22736 0 -1 28224
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _428_
timestamp 1698431365
transform 1 0 26432 0 1 30240
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  _429_
timestamp 1698431365
transform -1 0 31024 0 1 20160
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _430_
timestamp 1698431365
transform -1 0 30576 0 1 22176
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _431_
timestamp 1698431365
transform 1 0 24864 0 1 24192
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _432_
timestamp 1698431365
transform 1 0 25760 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _433_
timestamp 1698431365
transform 1 0 42224 0 -1 30240
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _434_
timestamp 1698431365
transform -1 0 31584 0 1 30240
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _435_
timestamp 1698431365
transform 1 0 29456 0 -1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  _436_
timestamp 1698431365
transform 1 0 31808 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _437_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _438_
timestamp 1698431365
transform 1 0 32704 0 1 38304
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _439_
timestamp 1698431365
transform 1 0 32928 0 -1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _440_
timestamp 1698431365
transform 1 0 36176 0 -1 32256
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  _441_
timestamp 1698431365
transform -1 0 35952 0 -1 30240
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  _442_
timestamp 1698431365
transform 1 0 32928 0 -1 30240
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_1  _443_
timestamp 1698431365
transform -1 0 30016 0 -1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _444_
timestamp 1698431365
transform -1 0 26432 0 1 30240
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _445_
timestamp 1698431365
transform 1 0 14672 0 1 32256
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _446_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _447_
timestamp 1698431365
transform 1 0 26320 0 -1 42336
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _448_
timestamp 1698431365
transform 1 0 28784 0 -1 40320
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _449_
timestamp 1698431365
transform -1 0 27552 0 -1 38304
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _450_
timestamp 1698431365
transform 1 0 27552 0 1 38304
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _451_
timestamp 1698431365
transform 1 0 46480 0 1 22176
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _452_
timestamp 1698431365
transform 1 0 49392 0 -1 18144
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _453_
timestamp 1698431365
transform 1 0 47376 0 1 24192
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _454_
timestamp 1698431365
transform 1 0 53536 0 1 22176
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _455_
timestamp 1698431365
transform 1 0 51744 0 -1 20160
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _456_
timestamp 1698431365
transform 1 0 50848 0 1 22176
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _457_
timestamp 1698431365
transform 1 0 45808 0 -1 26208
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  _458_
timestamp 1698431365
transform -1 0 28112 0 1 30240
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  _459_
timestamp 1698431365
transform -1 0 27328 0 1 32256
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _460_
timestamp 1698431365
transform 1 0 12544 0 -1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _461_
timestamp 1698431365
transform -1 0 20944 0 1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _462_
timestamp 1698431365
transform 1 0 21616 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__or4_1  _463_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 24528 0 -1 32256
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _464_
timestamp 1698431365
transform 1 0 20720 0 -1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _465_
timestamp 1698431365
transform 1 0 18704 0 1 30240
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _466_
timestamp 1698431365
transform 1 0 17248 0 1 30240
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _467_
timestamp 1698431365
transform 1 0 17920 0 -1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  _468_
timestamp 1698431365
transform 1 0 16800 0 1 32256
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _469_
timestamp 1698431365
transform -1 0 12992 0 1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _470_
timestamp 1698431365
transform -1 0 22848 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _471_
timestamp 1698431365
transform 1 0 21952 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  _472_
timestamp 1698431365
transform 1 0 21840 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__oai31_1  _473_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 21840 0 1 36288
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _474_
timestamp 1698431365
transform 1 0 22736 0 -1 36288
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _475_
timestamp 1698431365
transform -1 0 24864 0 -1 36288
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _476_
timestamp 1698431365
transform -1 0 28112 0 1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _477_
timestamp 1698431365
transform -1 0 30464 0 1 36288
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _478_
timestamp 1698431365
transform 1 0 20272 0 1 36288
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _479_
timestamp 1698431365
transform 1 0 21168 0 1 36288
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _480_
timestamp 1698431365
transform -1 0 26096 0 -1 36288
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _481_
timestamp 1698431365
transform -1 0 24528 0 1 34272
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  _482_
timestamp 1698431365
transform -1 0 23520 0 1 34272
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _483_
timestamp 1698431365
transform 1 0 23072 0 1 36288
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _484_
timestamp 1698431365
transform 1 0 21168 0 1 38304
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _485_
timestamp 1698431365
transform 1 0 17360 0 -1 40320
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _486_
timestamp 1698431365
transform 1 0 18032 0 1 38304
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _487_
timestamp 1698431365
transform 1 0 21952 0 -1 40320
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _488_
timestamp 1698431365
transform 1 0 19488 0 -1 38304
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _489_
timestamp 1698431365
transform 1 0 19488 0 1 38304
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  _490_
timestamp 1698431365
transform 1 0 19376 0 -1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  _491_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 14784 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__nand4_1  _492_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 21952 0 -1 38304
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _493_
timestamp 1698431365
transform 1 0 19376 0 1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _494_
timestamp 1698431365
transform 1 0 17920 0 -1 36288
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  _495_
timestamp 1698431365
transform 1 0 18032 0 1 36288
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _496_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29232 0 -1 36288
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _497_
timestamp 1698431365
transform 1 0 28560 0 -1 34272
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _498_
timestamp 1698431365
transform 1 0 29120 0 1 34272
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _499_
timestamp 1698431365
transform 1 0 26096 0 -1 36288
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _500_
timestamp 1698431365
transform 1 0 23072 0 1 32256
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _501_
timestamp 1698431365
transform 1 0 21728 0 -1 34272
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _502_
timestamp 1698431365
transform 1 0 22512 0 1 38304
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _503_
timestamp 1698431365
transform 1 0 16912 0 1 42336
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _504_
timestamp 1698431365
transform 1 0 17248 0 -1 44352
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _505_
timestamp 1698431365
transform -1 0 21504 0 -1 42336
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _506_
timestamp 1698431365
transform 1 0 17808 0 1 40320
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _507_
timestamp 1698431365
transform 1 0 18816 0 -1 40320
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _508_
timestamp 1698431365
transform 1 0 11200 0 -1 36288
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _509_
timestamp 1698431365
transform -1 0 20720 0 -1 32256
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _510_
timestamp 1698431365
transform 1 0 15680 0 1 34272
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  _511_
timestamp 1698431365
transform 1 0 14896 0 1 36288
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__tiel  _512_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 8736 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__tiel  _513_
timestamp 1698431365
transform -1 0 4480 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__tiel  _514_
timestamp 1698431365
transform 1 0 54992 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__tiel  _515_
timestamp 1698431365
transform -1 0 6160 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__tiel  _516_
timestamp 1698431365
transform -1 0 4928 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__248__I test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 35728 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__249__I
timestamp 1698431365
transform 1 0 34944 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__250__I
timestamp 1698431365
transform 1 0 36624 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__251__I
timestamp 1698431365
transform -1 0 29456 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__254__I
timestamp 1698431365
transform -1 0 35056 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__261__I
timestamp 1698431365
transform 1 0 33936 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__262__I
timestamp 1698431365
transform 1 0 26880 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__265__I
timestamp 1698431365
transform 1 0 37072 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__266__S1
timestamp 1698431365
transform -1 0 26432 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__267__I
timestamp 1698431365
transform 1 0 32032 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__274__I
timestamp 1698431365
transform 1 0 45136 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__280__S
timestamp 1698431365
transform 1 0 25312 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__281__A1
timestamp 1698431365
transform -1 0 23408 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__289__I
timestamp 1698431365
transform 1 0 35952 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__290__I
timestamp 1698431365
transform 1 0 43680 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__291__S1
timestamp 1698431365
transform 1 0 45248 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__292__I
timestamp 1698431365
transform 1 0 36400 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__293__I
timestamp 1698431365
transform 1 0 47936 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__295__S0
timestamp 1698431365
transform -1 0 50960 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__296__I
timestamp 1698431365
transform 1 0 47040 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__298__S0
timestamp 1698431365
transform 1 0 44464 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__298__S1
timestamp 1698431365
transform 1 0 44912 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__299__S0
timestamp 1698431365
transform 1 0 49168 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__301__S
timestamp 1698431365
transform -1 0 45024 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__302__A2
timestamp 1698431365
transform -1 0 28448 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__304__I
timestamp 1698431365
transform 1 0 27440 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__307__I
timestamp 1698431365
transform 1 0 35280 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__309__S
timestamp 1698431365
transform 1 0 27776 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__312__I
timestamp 1698431365
transform 1 0 37968 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__316__I
timestamp 1698431365
transform 1 0 40320 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__321__A2
timestamp 1698431365
transform 1 0 27552 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__325__I
timestamp 1698431365
transform -1 0 43680 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__327__S
timestamp 1698431365
transform 1 0 34496 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__328__I
timestamp 1698431365
transform 1 0 31024 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__329__A1
timestamp 1698431365
transform -1 0 27104 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__333__A2
timestamp 1698431365
transform 1 0 27328 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__337__I
timestamp 1698431365
transform 1 0 26432 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__342__I
timestamp 1698431365
transform 1 0 37520 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__349__S
timestamp 1698431365
transform -1 0 35840 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__353__S1
timestamp 1698431365
transform 1 0 42784 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__355__B
timestamp 1698431365
transform 1 0 36064 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__362__S0
timestamp 1698431365
transform -1 0 38640 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__364__S
timestamp 1698431365
transform -1 0 37296 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__367__S0
timestamp 1698431365
transform -1 0 48384 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__368__I
timestamp 1698431365
transform 1 0 49504 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__375__S
timestamp 1698431365
transform 1 0 48160 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__376__A2
timestamp 1698431365
transform 1 0 28336 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__380__S0
timestamp 1698431365
transform 1 0 42336 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__382__I
timestamp 1698431365
transform -1 0 43568 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__384__S
timestamp 1698431365
transform 1 0 39872 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__397__S
timestamp 1698431365
transform 1 0 34720 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__399__S1
timestamp 1698431365
transform 1 0 43904 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__401__B
timestamp 1698431365
transform 1 0 37072 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__405__I
timestamp 1698431365
transform 1 0 28896 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__406__S0
timestamp 1698431365
transform -1 0 40544 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__407__S1
timestamp 1698431365
transform 1 0 35280 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__408__S
timestamp 1698431365
transform -1 0 37072 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__412__I
timestamp 1698431365
transform -1 0 48384 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__418__S0
timestamp 1698431365
transform 1 0 50512 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__418__S1
timestamp 1698431365
transform 1 0 48832 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__420__S
timestamp 1698431365
transform 1 0 48160 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__421__A2
timestamp 1698431365
transform 1 0 29232 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__424__S0
timestamp 1698431365
transform 1 0 40992 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__426__S
timestamp 1698431365
transform 1 0 39424 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__438__S
timestamp 1698431365
transform 1 0 34384 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__442__B
timestamp 1698431365
transform 1 0 36176 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__447__S0
timestamp 1698431365
transform 1 0 30464 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__447__S1
timestamp 1698431365
transform 1 0 29792 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__452__S0
timestamp 1698431365
transform -1 0 49392 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__455__S0
timestamp 1698431365
transform 1 0 53088 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__455__S1
timestamp 1698431365
transform 1 0 53648 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__457__S
timestamp 1698431365
transform -1 0 45808 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__458__A2
timestamp 1698431365
transform 1 0 29680 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__470__I
timestamp 1698431365
transform 1 0 22176 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__471__I
timestamp 1698431365
transform 1 0 23520 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__472__I
timestamp 1698431365
transform -1 0 21840 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__473__B
timestamp 1698431365
transform -1 0 21392 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__475__I0
timestamp 1698431365
transform 1 0 22512 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__476__I0
timestamp 1698431365
transform 1 0 28112 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__477__I0
timestamp 1698431365
transform 1 0 30688 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__478__I
timestamp 1698431365
transform 1 0 20048 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__483__I0
timestamp 1698431365
transform -1 0 23296 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__483__I1
timestamp 1698431365
transform 1 0 24752 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__485__I0
timestamp 1698431365
transform -1 0 16576 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__485__I1
timestamp 1698431365
transform 1 0 16800 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__486__I0
timestamp 1698431365
transform -1 0 17136 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__486__I1
timestamp 1698431365
transform 1 0 17808 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__487__I0
timestamp 1698431365
transform -1 0 21952 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__487__I1
timestamp 1698431365
transform 1 0 21840 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__488__I0
timestamp 1698431365
transform 1 0 17360 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__488__I1
timestamp 1698431365
transform -1 0 19488 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__489__I0
timestamp 1698431365
transform -1 0 16688 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__489__I1
timestamp 1698431365
transform 1 0 21392 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__492__A1
timestamp 1698431365
transform 1 0 18368 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__492__A2
timestamp 1698431365
transform 1 0 17472 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__492__A3
timestamp 1698431365
transform 1 0 16800 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__492__A4
timestamp 1698431365
transform 1 0 18816 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__493__I0
timestamp 1698431365
transform 1 0 19152 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__494__I0
timestamp 1698431365
transform 1 0 20496 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__495__I0
timestamp 1698431365
transform 1 0 17920 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__496__CLK
timestamp 1698431365
transform 1 0 28560 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__497__CLK
timestamp 1698431365
transform 1 0 27664 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__498__CLK
timestamp 1698431365
transform 1 0 28560 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__499__CLK
timestamp 1698431365
transform 1 0 25872 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__500__CLK
timestamp 1698431365
transform 1 0 22400 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__501__CLK
timestamp 1698431365
transform 1 0 21504 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__502__CLK
timestamp 1698431365
transform 1 0 22288 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__503__CLK
timestamp 1698431365
transform 1 0 16688 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__504__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__505__CLK
timestamp 1698431365
transform 1 0 18144 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__506__CLK
timestamp 1698431365
transform 1 0 17136 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__507__CLK
timestamp 1698431365
transform 1 0 17584 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__508__CLK
timestamp 1698431365
transform 1 0 10976 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__509__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__510__CLK
timestamp 1698431365
transform 1 0 15456 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__511__CLK
timestamp 1698431365
transform 1 0 14672 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_1_inst_A
timestamp 1698431365
transform 1 0 41888 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_1_inst_B
timestamp 1698431365
transform 1 0 40320 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_1_inst_CI
timestamp 1698431365
transform 1 0 40320 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_2_inst_A
timestamp 1698431365
transform 1 0 45584 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_2_inst_B
timestamp 1698431365
transform 1 0 47488 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_2_inst_CI
timestamp 1698431365
transform 1 0 45136 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_4_inst_A
timestamp 1698431365
transform 1 0 45472 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_4_inst_B
timestamp 1698431365
transform 1 0 46032 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addf_4_inst_CI
timestamp 1698431365
transform 1 0 45584 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addh_1_inst_A
timestamp 1698431365
transform 1 0 45584 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addh_1_inst_B
timestamp 1698431365
transform 1 0 46032 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addh_2_inst_A
timestamp 1698431365
transform 1 0 37296 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addh_2_inst_B
timestamp 1698431365
transform 1 0 37296 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addh_4_inst_A
timestamp 1698431365
transform 1 0 44800 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.addh_4_inst_B
timestamp 1698431365
transform 1 0 44240 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and2_1_inst_A1
timestamp 1698431365
transform 1 0 31136 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and2_1_inst_A2
timestamp 1698431365
transform 1 0 28560 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and2_2_inst_A1
timestamp 1698431365
transform 1 0 51072 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and2_2_inst_A2
timestamp 1698431365
transform 1 0 50624 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and2_4_inst_A1
timestamp 1698431365
transform 1 0 34160 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and2_4_inst_A2
timestamp 1698431365
transform 1 0 33040 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_1_inst_A1
timestamp 1698431365
transform 1 0 50400 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_1_inst_A2
timestamp 1698431365
transform 1 0 49056 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_1_inst_A3
timestamp 1698431365
transform 1 0 49952 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_2_inst_A1
timestamp 1698431365
transform 1 0 36400 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_2_inst_A2
timestamp 1698431365
transform 1 0 29344 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_2_inst_A3
timestamp 1698431365
transform 1 0 29568 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_4_inst_A1
timestamp 1698431365
transform 1 0 53200 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_4_inst_A2
timestamp 1698431365
transform 1 0 50176 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_4_inst_A3
timestamp 1698431365
transform 1 0 49728 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_1_inst_A1
timestamp 1698431365
transform 1 0 20160 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_1_inst_A2
timestamp 1698431365
transform 1 0 22288 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_1_inst_A3
timestamp 1698431365
transform 1 0 21840 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_1_inst_A4
timestamp 1698431365
transform 1 0 21392 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_2_inst_A1
timestamp 1698431365
transform 1 0 50848 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_2_inst_A2
timestamp 1698431365
transform 1 0 49504 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_2_inst_A3
timestamp 1698431365
transform 1 0 49056 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_2_inst_A4
timestamp 1698431365
transform 1 0 48832 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_4_inst_A1
timestamp 1698431365
transform 1 0 35504 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_4_inst_A2
timestamp 1698431365
transform 1 0 33488 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_4_inst_A3
timestamp 1698431365
transform 1 0 28560 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_4_inst_A4
timestamp 1698431365
transform 1 0 31920 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_1_inst_A1
timestamp 1698431365
transform 1 0 25424 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_1_inst_A2
timestamp 1698431365
transform 1 0 24192 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_1_inst_B
timestamp 1698431365
transform 1 0 23744 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_2_inst_A1
timestamp 1698431365
transform 1 0 57680 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_2_inst_A2
timestamp 1698431365
transform 1 0 56672 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_2_inst_B
timestamp 1698431365
transform 1 0 58128 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_4_inst_A1
timestamp 1698431365
transform 1 0 25872 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_4_inst_A2
timestamp 1698431365
transform 1 0 22848 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi21_4_inst_B
timestamp 1698431365
transform 1 0 19376 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_1_inst_A1
timestamp 1698431365
transform 1 0 56672 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_1_inst_A2
timestamp 1698431365
transform 1 0 58128 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_1_inst_B1
timestamp 1698431365
transform 1 0 55776 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_1_inst_B2
timestamp 1698431365
transform 1 0 57680 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_2_inst_A1
timestamp 1698431365
transform 1 0 26880 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_2_inst_A2
timestamp 1698431365
transform 1 0 22960 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_2_inst_B1
timestamp 1698431365
transform 1 0 24640 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_2_inst_B2
timestamp 1698431365
transform 1 0 22512 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_4_inst_A1
timestamp 1698431365
transform 1 0 51184 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_4_inst_A2
timestamp 1698431365
transform 1 0 50064 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_4_inst_B1
timestamp 1698431365
transform 1 0 50960 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_4_inst_B2
timestamp 1698431365
transform 1 0 50512 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_1_inst_A1
timestamp 1698431365
transform 1 0 25872 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_1_inst_A2
timestamp 1698431365
transform 1 0 22624 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_1_inst_B
timestamp 1698431365
transform 1 0 24192 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_1_inst_C
timestamp 1698431365
transform 1 0 24192 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_2_inst_A1
timestamp 1698431365
transform 1 0 54208 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_2_inst_A2
timestamp 1698431365
transform 1 0 57120 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_2_inst_B
timestamp 1698431365
transform 1 0 53760 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_2_inst_C
timestamp 1698431365
transform 1 0 53312 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_4_inst_A1
timestamp 1698431365
transform 1 0 24080 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_4_inst_A2
timestamp 1698431365
transform 1 0 19824 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_4_inst_B
timestamp 1698431365
transform 1 0 23296 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi211_4_inst_C
timestamp 1698431365
transform 1 0 24528 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_1_inst_A1
timestamp 1698431365
transform 1 0 58128 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_1_inst_A2
timestamp 1698431365
transform 1 0 57120 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_1_inst_B1
timestamp 1698431365
transform 1 0 56000 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_1_inst_B2
timestamp 1698431365
transform 1 0 55552 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_1_inst_C
timestamp 1698431365
transform 1 0 55104 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_2_inst_A1
timestamp 1698431365
transform 1 0 24640 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_2_inst_A2
timestamp 1698431365
transform 1 0 20272 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_2_inst_B1
timestamp 1698431365
transform 1 0 19824 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_2_inst_B2
timestamp 1698431365
transform 1 0 19824 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_2_inst_C
timestamp 1698431365
transform 1 0 20496 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_4_inst_A1
timestamp 1698431365
transform 1 0 56000 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_4_inst_A2
timestamp 1698431365
transform 1 0 55664 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_4_inst_B1
timestamp 1698431365
transform 1 0 52080 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_4_inst_B2
timestamp 1698431365
transform 1 0 52752 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_4_inst_C
timestamp 1698431365
transform 1 0 52080 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_1_inst_A1
timestamp 1698431365
transform 1 0 22064 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_1_inst_A2
timestamp 1698431365
transform 1 0 21616 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_1_inst_B1
timestamp 1698431365
transform 1 0 22400 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_1_inst_B2
timestamp 1698431365
transform 1 0 20720 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_1_inst_C1
timestamp 1698431365
transform 1 0 20272 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_1_inst_C2
timestamp 1698431365
transform 1 0 22064 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_2_inst_A1
timestamp 1698431365
transform 1 0 55552 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_2_inst_A2
timestamp 1698431365
transform 1 0 52752 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_2_inst_B1
timestamp 1698431365
transform 1 0 52080 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_2_inst_B2
timestamp 1698431365
transform 1 0 51632 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_2_inst_C1
timestamp 1698431365
transform 1 0 50736 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_2_inst_C2
timestamp 1698431365
transform 1 0 51184 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_4_inst_A1
timestamp 1698431365
transform 1 0 27328 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_4_inst_A2
timestamp 1698431365
transform 1 0 20944 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_4_inst_B1
timestamp 1698431365
transform 1 0 21392 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_4_inst_B2
timestamp 1698431365
transform 1 0 28112 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_4_inst_C1
timestamp 1698431365
transform 1 0 20496 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi222_4_inst_C2
timestamp 1698431365
transform 1 0 27664 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_1_inst_I
timestamp 1698431365
transform 1 0 35168 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_2_inst_I
timestamp 1698431365
transform 1 0 55552 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_3_inst_I
timestamp 1698431365
transform 1 0 32704 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_4_inst_I
timestamp 1698431365
transform 1 0 52976 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_8_inst_I
timestamp 1698431365
transform 1 0 32480 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_12_inst_I
timestamp 1698431365
transform 1 0 55440 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_16_inst_I
timestamp 1698431365
transform 1 0 18144 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.buf_20_inst_I
timestamp 1698431365
transform 1 0 48160 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_1_inst_EN
timestamp 1698431365
transform 1 0 38976 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_1_inst_I
timestamp 1698431365
transform 1 0 38528 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_2_inst_EN
timestamp 1698431365
transform 1 0 37072 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_2_inst_I
timestamp 1698431365
transform 1 0 36400 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_3_inst_EN
timestamp 1698431365
transform 1 0 32256 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_3_inst_I
timestamp 1698431365
transform 1 0 34048 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_4_inst_EN
timestamp 1698431365
transform 1 0 47600 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_4_inst_I
timestamp 1698431365
transform 1 0 45584 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_8_inst_EN
timestamp 1698431365
transform 1 0 43568 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_8_inst_I
timestamp 1698431365
transform 1 0 44016 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_12_inst_EN
timestamp 1698431365
transform 1 0 44464 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_12_inst_I
timestamp 1698431365
transform 1 0 44912 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_16_inst_EN
timestamp 1698431365
transform 1 0 41104 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_16_inst_I
timestamp 1698431365
transform 1 0 41552 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_1_inst_I
timestamp 1698431365
transform 1 0 40320 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_2_inst_I
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_3_inst_I
timestamp 1698431365
transform 1 0 42896 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_4_inst_I
timestamp 1698431365
transform 1 0 32480 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_8_inst_I
timestamp 1698431365
transform 1 0 20720 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_12_inst_I
timestamp 1698431365
transform 1 0 40320 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_16_inst_I
timestamp 1698431365
transform 1 0 19152 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkbuf_20_inst_I
timestamp 1698431365
transform 1 0 17472 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_1_inst_I
timestamp 1698431365
transform 1 0 23408 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_2_inst_I
timestamp 1698431365
transform 1 0 28560 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_3_inst_I
timestamp 1698431365
transform 1 0 22288 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_4_inst_I
timestamp 1698431365
transform 1 0 26096 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_8_inst_I
timestamp 1698431365
transform 1 0 20272 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_12_inst_I
timestamp 1698431365
transform 1 0 41776 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_16_inst_I
timestamp 1698431365
transform 1 0 17584 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.clkinv_20_inst_I
timestamp 1698431365
transform 1 0 18928 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnq_1_inst_CLKN
timestamp 1698431365
transform 1 0 25536 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnq_1_inst_D
timestamp 1698431365
transform 1 0 24640 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnq_2_inst_CLKN
timestamp 1698431365
transform 1 0 21840 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnq_2_inst_D
timestamp 1698431365
transform 1 0 21392 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnq_4_inst_CLKN
timestamp 1698431365
transform 1 0 33712 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnq_4_inst_D
timestamp 1698431365
transform 1 0 32368 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_CLKN
timestamp 1698431365
transform 1 0 38304 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_D
timestamp 1698431365
transform 1 0 39200 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_RN
timestamp 1698431365
transform 1 0 38752 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_CLKN
timestamp 1698431365
transform 1 0 38864 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_D
timestamp 1698431365
transform 1 0 39312 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_RN
timestamp 1698431365
transform 1 0 39760 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_CLKN
timestamp 1698431365
transform 1 0 38976 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_D
timestamp 1698431365
transform 1 0 39872 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_RN
timestamp 1698431365
transform 1 0 39424 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_CLKN
timestamp 1698431365
transform 1 0 29456 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_D
timestamp 1698431365
transform 1 0 28560 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_RN
timestamp 1698431365
transform 1 0 29232 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 27776 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_CLKN
timestamp 1698431365
transform 1 0 37856 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_D
timestamp 1698431365
transform 1 0 36400 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_RN
timestamp 1698431365
transform 1 0 37632 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 37184 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_CLKN
timestamp 1698431365
transform 1 0 27328 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_D
timestamp 1698431365
transform 1 0 23072 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_RN
timestamp 1698431365
transform 1 0 22624 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 22176 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_CLKN
timestamp 1698431365
transform 1 0 18480 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_D
timestamp 1698431365
transform 1 0 18928 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 20608 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_CLKN
timestamp 1698431365
transform 1 0 28336 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_D
timestamp 1698431365
transform 1 0 27888 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 27440 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_CLKN
timestamp 1698431365
transform 1 0 34720 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_D
timestamp 1698431365
transform 1 0 35616 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 35168 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffq_1_inst_CLK
timestamp 1698431365
transform 1 0 37520 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffq_1_inst_D
timestamp 1698431365
transform 1 0 37072 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffq_2_inst_CLK
timestamp 1698431365
transform 1 0 36960 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffq_2_inst_D
timestamp 1698431365
transform 1 0 36400 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffq_4_inst_CLK
timestamp 1698431365
transform 1 0 27664 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffq_4_inst_D
timestamp 1698431365
transform 1 0 27216 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_1_inst_CLK
timestamp 1698431365
transform 1 0 35840 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_1_inst_D
timestamp 1698431365
transform 1 0 35616 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_1_inst_RN
timestamp 1698431365
transform 1 0 35616 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_2_inst_CLK
timestamp 1698431365
transform 1 0 26320 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_2_inst_D
timestamp 1698431365
transform 1 0 22064 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_2_inst_RN
timestamp 1698431365
transform 1 0 21616 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_4_inst_CLK
timestamp 1698431365
transform 1 0 22848 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_4_inst_D
timestamp 1698431365
transform 1 0 22400 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrnq_4_inst_RN
timestamp 1698431365
transform 1 0 21952 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_CLK
timestamp 1698431365
transform 1 0 28448 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_D
timestamp 1698431365
transform 1 0 26992 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_RN
timestamp 1698431365
transform 1 0 28896 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 27664 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_CLK
timestamp 1698431365
transform 1 0 37520 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_D
timestamp 1698431365
transform 1 0 37072 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_RN
timestamp 1698431365
transform 1 0 36624 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 36176 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_CLK
timestamp 1698431365
transform 1 0 36400 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_D
timestamp 1698431365
transform 1 0 35952 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_RN
timestamp 1698431365
transform 1 0 35504 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 35168 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_1_inst_CLK
timestamp 1698431365
transform 1 0 35392 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_1_inst_D
timestamp 1698431365
transform 1 0 36288 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 35840 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_2_inst_CLK
timestamp 1698431365
transform 1 0 26880 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_2_inst_D
timestamp 1698431365
transform 1 0 27552 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 26432 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_4_inst_CLK
timestamp 1698431365
transform 1 0 34608 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_4_inst_D
timestamp 1698431365
transform 1 0 35504 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 35056 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlya_1_inst_I
timestamp 1698431365
transform 1 0 18928 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlya_2_inst_I
timestamp 1698431365
transform 1 0 26320 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlya_4_inst_I
timestamp 1698431365
transform 1 0 30576 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyb_1_inst_I
timestamp 1698431365
transform 1 0 33488 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyb_2_inst_I
timestamp 1698431365
transform 1 0 40208 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyb_4_inst_I
timestamp 1698431365
transform 1 0 37184 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyc_1_inst_I
timestamp 1698431365
transform 1 0 38080 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyc_2_inst_I
timestamp 1698431365
transform 1 0 30016 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyc_4_inst_I
timestamp 1698431365
transform 1 0 20944 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyd_1_inst_I
timestamp 1698431365
transform 1 0 25424 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyd_2_inst_I
timestamp 1698431365
transform 1 0 29232 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.dlyd_4_inst_I
timestamp 1698431365
transform 1 0 32704 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_1_inst_CLKN
timestamp 1698431365
transform 1 0 20944 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_1_inst_E
timestamp 1698431365
transform 1 0 21840 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_1_inst_TE
timestamp 1698431365
transform 1 0 21392 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_2_inst_CLKN
timestamp 1698431365
transform 1 0 27328 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_2_inst_E
timestamp 1698431365
transform 1 0 23520 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_2_inst_TE
timestamp 1698431365
transform 1 0 23072 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_4_inst_CLKN
timestamp 1698431365
transform 1 0 20272 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_4_inst_E
timestamp 1698431365
transform 1 0 20720 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_4_inst_TE
timestamp 1698431365
transform 1 0 22736 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_1_inst_CLK
timestamp 1698431365
transform 1 0 28112 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_1_inst_E
timestamp 1698431365
transform 1 0 24640 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_1_inst_TE
timestamp 1698431365
transform 1 0 24192 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_2_inst_CLK
timestamp 1698431365
transform 1 0 18816 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_2_inst_E
timestamp 1698431365
transform 1 0 20720 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_2_inst_TE
timestamp 1698431365
transform 1 0 21616 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_4_inst_CLK
timestamp 1698431365
transform 1 0 27440 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_4_inst_E
timestamp 1698431365
transform 1 0 27888 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_4_inst_TE
timestamp 1698431365
transform 1 0 27328 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_1_inst_I
timestamp 1698431365
transform 1 0 32032 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_2_inst_I
timestamp 1698431365
transform 1 0 55776 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_3_inst_I
timestamp 1698431365
transform 1 0 34720 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_4_inst_I
timestamp 1698431365
transform 1 0 52752 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_8_inst_I
timestamp 1698431365
transform 1 0 32144 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_12_inst_I
timestamp 1698431365
transform 1 0 53200 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_16_inst_I
timestamp 1698431365
transform 1 0 19376 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.inv_20_inst_I
timestamp 1698431365
transform 1 0 47152 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_1_inst_EN
timestamp 1698431365
transform 1 0 45360 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_1_inst_I
timestamp 1698431365
transform 1 0 45136 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_2_inst_EN
timestamp 1698431365
transform 1 0 44912 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_2_inst_I
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_3_inst_EN
timestamp 1698431365
transform 1 0 45360 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_3_inst_I
timestamp 1698431365
transform 1 0 43792 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_4_inst_EN
timestamp 1698431365
transform 1 0 43456 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_4_inst_I
timestamp 1698431365
transform 1 0 43904 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_8_inst_EN
timestamp 1698431365
transform 1 0 30800 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_8_inst_I
timestamp 1698431365
transform 1 0 31248 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_12_inst_EN
timestamp 1698431365
transform 1 0 30128 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.invz_12_inst_I
timestamp 1698431365
transform 1 0 29680 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latq_1_inst_D
timestamp 1698431365
transform 1 0 46704 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latq_1_inst_E
timestamp 1698431365
transform 1 0 46704 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latq_2_inst_D
timestamp 1698431365
transform 1 0 41440 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latq_2_inst_E
timestamp 1698431365
transform 1 0 40992 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latq_4_inst_D
timestamp 1698431365
transform 1 0 48272 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latq_4_inst_E
timestamp 1698431365
transform 1 0 48720 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_1_inst_D
timestamp 1698431365
transform 1 0 39872 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_1_inst_E
timestamp 1698431365
transform 1 0 40320 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_1_inst_RN
timestamp 1698431365
transform 1 0 40544 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_2_inst_D
timestamp 1698431365
transform 1 0 44912 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_2_inst_E
timestamp 1698431365
transform 1 0 44576 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_2_inst_RN
timestamp 1698431365
transform 1 0 44128 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_4_inst_D
timestamp 1698431365
transform 1 0 22736 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_4_inst_E
timestamp 1698431365
transform 1 0 23632 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrnq_4_inst_RN
timestamp 1698431365
transform 1 0 23184 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_1_inst_D
timestamp 1698431365
transform 1 0 33264 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_1_inst_E
timestamp 1698431365
transform 1 0 32816 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_1_inst_RN
timestamp 1698431365
transform 1 0 31920 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 32368 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_2_inst_D
timestamp 1698431365
transform 1 0 40320 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_2_inst_E
timestamp 1698431365
transform 1 0 41888 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_2_inst_RN
timestamp 1698431365
transform 1 0 41440 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 40992 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_4_inst_D
timestamp 1698431365
transform 1 0 40208 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_4_inst_E
timestamp 1698431365
transform 1 0 42336 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_4_inst_RN
timestamp 1698431365
transform 1 0 41888 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latrsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 40768 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_1_inst_D
timestamp 1698431365
transform 1 0 42224 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_1_inst_E
timestamp 1698431365
transform 1 0 41776 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 41328 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_2_inst_D
timestamp 1698431365
transform 1 0 33152 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_2_inst_E
timestamp 1698431365
transform 1 0 32480 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 32256 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_4_inst_D
timestamp 1698431365
transform 1 0 41664 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_4_inst_E
timestamp 1698431365
transform 1 0 41216 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.latsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 40768 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_1_inst_I0
timestamp 1698431365
transform 1 0 54656 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_1_inst_I1
timestamp 1698431365
transform 1 0 50960 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_1_inst_S
timestamp 1698431365
transform 1 0 51072 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_2_inst_I0
timestamp 1698431365
transform 1 0 43232 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_2_inst_I1
timestamp 1698431365
transform 1 0 39872 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_2_inst_S
timestamp 1698431365
transform 1 0 41664 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_4_inst_I0
timestamp 1698431365
transform 1 0 44800 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_4_inst_I1
timestamp 1698431365
transform 1 0 45696 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux2_4_inst_S
timestamp 1698431365
transform 1 0 45248 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_1_inst_I0
timestamp 1698431365
transform 1 0 29680 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_1_inst_I1
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_1_inst_I2
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_1_inst_I3
timestamp 1698431365
transform 1 0 26768 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_1_inst_S0
timestamp 1698431365
transform 1 0 27664 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_1_inst_S1
timestamp 1698431365
transform 1 0 25760 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_2_inst_I0
timestamp 1698431365
transform 1 0 39648 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_2_inst_I1
timestamp 1698431365
transform 1 0 39200 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_2_inst_I2
timestamp 1698431365
transform 1 0 38752 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_2_inst_I3
timestamp 1698431365
transform 1 0 37632 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_2_inst_S0
timestamp 1698431365
transform 1 0 38528 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_2_inst_S1
timestamp 1698431365
transform 1 0 38080 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_4_inst_I0
timestamp 1698431365
transform 1 0 36960 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_4_inst_I1
timestamp 1698431365
transform 1 0 36736 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_4_inst_I2
timestamp 1698431365
transform 1 0 36288 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_4_inst_I3
timestamp 1698431365
transform 1 0 35168 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_4_inst_S0
timestamp 1698431365
transform 1 0 36064 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.mux4_4_inst_S1
timestamp 1698431365
transform 1 0 35616 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand2_1_inst_A1
timestamp 1698431365
transform 1 0 53424 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand2_1_inst_A2
timestamp 1698431365
transform 1 0 52304 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand2_2_inst_A1
timestamp 1698431365
transform 1 0 35952 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand2_2_inst_A2
timestamp 1698431365
transform 1 0 34608 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand2_4_inst_A1
timestamp 1698431365
transform 1 0 47936 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand2_4_inst_A2
timestamp 1698431365
transform 1 0 48384 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_1_inst_A1
timestamp 1698431365
transform 1 0 28896 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_1_inst_A2
timestamp 1698431365
transform 1 0 28448 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_1_inst_A3
timestamp 1698431365
transform 1 0 28000 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_2_inst_A1
timestamp 1698431365
transform 1 0 49280 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_2_inst_A2
timestamp 1698431365
transform 1 0 48832 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_2_inst_A3
timestamp 1698431365
transform 1 0 47936 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_4_inst_A1
timestamp 1698431365
transform 1 0 25312 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_4_inst_A2
timestamp 1698431365
transform 1 0 20608 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_4_inst_A3
timestamp 1698431365
transform 1 0 20384 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_1_inst_A1
timestamp 1698431365
transform 1 0 48608 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_1_inst_A2
timestamp 1698431365
transform 1 0 47376 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_1_inst_A3
timestamp 1698431365
transform 1 0 46928 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_1_inst_A4
timestamp 1698431365
transform 1 0 46704 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_2_inst_A1
timestamp 1698431365
transform 1 0 42224 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_2_inst_A2
timestamp 1698431365
transform 1 0 41776 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_2_inst_A3
timestamp 1698431365
transform 1 0 41328 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_2_inst_A4
timestamp 1698431365
transform 1 0 39984 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_4_inst_A1
timestamp 1698431365
transform 1 0 54208 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_4_inst_A2
timestamp 1698431365
transform 1 0 57120 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_4_inst_A3
timestamp 1698431365
transform 1 0 58016 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand4_4_inst_A4
timestamp 1698431365
transform 1 0 56672 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor2_1_inst_A1
timestamp 1698431365
transform 1 0 42000 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor2_1_inst_A2
timestamp 1698431365
transform 1 0 40992 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor2_2_inst_A1
timestamp 1698431365
transform 1 0 57568 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor2_2_inst_A2
timestamp 1698431365
transform 1 0 57792 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor2_4_inst_A1
timestamp 1698431365
transform 1 0 38864 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor2_4_inst_A2
timestamp 1698431365
transform 1 0 38416 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_1_inst_A1
timestamp 1698431365
transform 1 0 58128 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_1_inst_A2
timestamp 1698431365
transform 1 0 57120 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_1_inst_A3
timestamp 1698431365
transform 1 0 56672 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_2_inst_A1
timestamp 1698431365
transform 1 0 22960 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_2_inst_A2
timestamp 1698431365
transform 1 0 20272 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_2_inst_A3
timestamp 1698431365
transform 1 0 19824 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_4_inst_A1
timestamp 1698431365
transform 1 0 46256 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_4_inst_A2
timestamp 1698431365
transform 1 0 45808 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor3_4_inst_A3
timestamp 1698431365
transform 1 0 45360 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_1_inst_A1
timestamp 1698431365
transform 1 0 42672 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_1_inst_A2
timestamp 1698431365
transform 1 0 41440 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_1_inst_A3
timestamp 1698431365
transform 1 0 40992 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_1_inst_A4
timestamp 1698431365
transform 1 0 38192 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_2_inst_A1
timestamp 1698431365
transform 1 0 57568 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_2_inst_A2
timestamp 1698431365
transform 1 0 57568 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_2_inst_A3
timestamp 1698431365
transform 1 0 57120 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_2_inst_A4
timestamp 1698431365
transform 1 0 56000 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_4_inst_A1
timestamp 1698431365
transform 1 0 39536 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_4_inst_A2
timestamp 1698431365
transform 1 0 39424 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_4_inst_A3
timestamp 1698431365
transform 1 0 39088 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.nor4_4_inst_A4
timestamp 1698431365
transform 1 0 38640 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_1_inst_A1
timestamp 1698431365
transform 1 0 51520 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_1_inst_A2
timestamp 1698431365
transform 1 0 51968 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_1_inst_B
timestamp 1698431365
transform 1 0 53984 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_2_inst_A1
timestamp 1698431365
transform 1 0 29232 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_2_inst_A2
timestamp 1698431365
transform 1 0 28560 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_2_inst_B
timestamp 1698431365
transform 1 0 27216 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_4_inst_A1
timestamp 1698431365
transform 1 0 51520 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_4_inst_A2
timestamp 1698431365
transform 1 0 52416 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai21_4_inst_B
timestamp 1698431365
transform 1 0 51968 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_1_inst_A1
timestamp 1698431365
transform 1 0 29904 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_1_inst_A2
timestamp 1698431365
transform 1 0 29456 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_1_inst_B1
timestamp 1698431365
transform 1 0 33936 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_1_inst_B2
timestamp 1698431365
transform 1 0 28560 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_2_inst_A1
timestamp 1698431365
transform 1 0 50624 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_2_inst_A2
timestamp 1698431365
transform 1 0 47712 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_2_inst_B1
timestamp 1698431365
transform 1 0 49728 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_2_inst_B2
timestamp 1698431365
transform 1 0 49280 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_4_inst_A1
timestamp 1698431365
transform 1 0 27216 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_4_inst_A2
timestamp 1698431365
transform 1 0 26768 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_4_inst_B1
timestamp 1698431365
transform 1 0 26320 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_4_inst_B2
timestamp 1698431365
transform 1 0 26880 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_1_inst_A1
timestamp 1698431365
transform 1 0 47488 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_1_inst_A2
timestamp 1698431365
transform 1 0 48832 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_1_inst_A3
timestamp 1698431365
transform 1 0 47488 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_1_inst_B
timestamp 1698431365
transform 1 0 46368 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_2_inst_A1
timestamp 1698431365
transform 1 0 24640 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_2_inst_A2
timestamp 1698431365
transform 1 0 22736 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_2_inst_A3
timestamp 1698431365
transform 1 0 23184 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_2_inst_B
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_4_inst_A1
timestamp 1698431365
transform 1 0 51184 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_4_inst_A2
timestamp 1698431365
transform 1 0 52752 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_4_inst_A3
timestamp 1698431365
transform 1 0 52080 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_4_inst_B
timestamp 1698431365
transform 1 0 51632 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_1_inst_A1
timestamp 1698431365
transform 1 0 32256 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_1_inst_A2
timestamp 1698431365
transform 1 0 33488 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_1_inst_A3
timestamp 1698431365
transform 1 0 28112 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_1_inst_B1
timestamp 1698431365
transform 1 0 28896 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_1_inst_B2
timestamp 1698431365
transform 1 0 27664 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_2_inst_A1
timestamp 1698431365
transform 1 0 53200 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_2_inst_A2
timestamp 1698431365
transform 1 0 52752 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_2_inst_A3
timestamp 1698431365
transform 1 0 52080 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_2_inst_B1
timestamp 1698431365
transform 1 0 53872 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_2_inst_B2
timestamp 1698431365
transform 1 0 51520 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_4_inst_A1
timestamp 1698431365
transform 1 0 29568 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_4_inst_A2
timestamp 1698431365
transform 1 0 28560 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_4_inst_A3
timestamp 1698431365
transform 1 0 27664 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_4_inst_B1
timestamp 1698431365
transform 1 0 27216 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai32_4_inst_B2
timestamp 1698431365
transform 1 0 27328 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_A1
timestamp 1698431365
transform 1 0 51520 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_A2
timestamp 1698431365
transform 1 0 51072 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_A3
timestamp 1698431365
transform 1 0 50624 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_B1
timestamp 1698431365
transform 1 0 50176 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_B2
timestamp 1698431365
transform 1 0 49728 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_B3
timestamp 1698431365
transform 1 0 49280 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_2_inst_A1
timestamp 1698431365
transform 1 0 28448 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_2_inst_A2
timestamp 1698431365
transform 1 0 28000 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_2_inst_A3
timestamp 1698431365
transform 1 0 27552 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_2_inst_B1
timestamp 1698431365
transform 1 0 28112 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_2_inst_B2
timestamp 1698431365
transform 1 0 26432 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_2_inst_B3
timestamp 1698431365
transform 1 0 25984 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_4_inst_A1
timestamp 1698431365
transform 1 0 47152 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_4_inst_A2
timestamp 1698431365
transform 1 0 46704 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_4_inst_A3
timestamp 1698431365
transform 1 0 46256 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_4_inst_B1
timestamp 1698431365
transform 1 0 45808 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_4_inst_B2
timestamp 1698431365
transform 1 0 45696 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_4_inst_B3
timestamp 1698431365
transform 1 0 45248 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_1_inst_A1
timestamp 1698431365
transform 1 0 29680 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_1_inst_A2
timestamp 1698431365
transform 1 0 30128 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_1_inst_B
timestamp 1698431365
transform 1 0 29232 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_1_inst_C
timestamp 1698431365
transform 1 0 28784 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_2_inst_A1
timestamp 1698431365
transform 1 0 44352 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_2_inst_A2
timestamp 1698431365
transform 1 0 42336 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_2_inst_B
timestamp 1698431365
transform 1 0 41888 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_2_inst_C
timestamp 1698431365
transform 1 0 40320 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_4_inst_A1
timestamp 1698431365
transform 1 0 39648 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_4_inst_A2
timestamp 1698431365
transform 1 0 39200 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_4_inst_B
timestamp 1698431365
transform 1 0 38752 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai211_4_inst_C
timestamp 1698431365
transform 1 0 39088 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_1_inst_A1
timestamp 1698431365
transform 1 0 50176 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_1_inst_A2
timestamp 1698431365
transform 1 0 48160 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_1_inst_B1
timestamp 1698431365
transform 1 0 49728 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_1_inst_B2
timestamp 1698431365
transform 1 0 49280 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_1_inst_C
timestamp 1698431365
transform 1 0 48832 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_2_inst_A1
timestamp 1698431365
transform 1 0 46592 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_2_inst_A2
timestamp 1698431365
transform 1 0 45584 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_2_inst_B1
timestamp 1698431365
transform 1 0 44128 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_2_inst_B2
timestamp 1698431365
transform 1 0 44016 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_2_inst_C
timestamp 1698431365
transform 1 0 43568 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_4_inst_A1
timestamp 1698431365
transform 1 0 54880 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_4_inst_A2
timestamp 1698431365
transform 1 0 52528 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_4_inst_B1
timestamp 1698431365
transform 1 0 50512 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_4_inst_B2
timestamp 1698431365
transform 1 0 52752 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai221_4_inst_C
timestamp 1698431365
transform 1 0 52752 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_1_inst_A1
timestamp 1698431365
transform 1 0 46368 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_1_inst_A2
timestamp 1698431365
transform 1 0 47040 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_1_inst_B1
timestamp 1698431365
transform 1 0 45920 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_1_inst_B2
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_1_inst_C1
timestamp 1698431365
transform 1 0 43792 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_1_inst_C2
timestamp 1698431365
transform 1 0 43344 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_2_inst_A1
timestamp 1698431365
transform 1 0 47040 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_2_inst_A2
timestamp 1698431365
transform 1 0 47824 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_2_inst_B1
timestamp 1698431365
transform 1 0 45472 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_2_inst_B2
timestamp 1698431365
transform 1 0 46816 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_2_inst_C1
timestamp 1698431365
transform 1 0 46368 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_2_inst_C2
timestamp 1698431365
transform 1 0 45920 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_4_inst_A1
timestamp 1698431365
transform 1 0 26768 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_4_inst_A2
timestamp 1698431365
transform 1 0 27216 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_4_inst_B1
timestamp 1698431365
transform 1 0 26320 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_4_inst_B2
timestamp 1698431365
transform 1 0 25424 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_4_inst_C1
timestamp 1698431365
transform 1 0 25312 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai222_4_inst_C2
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or2_1_inst_A1
timestamp 1698431365
transform 1 0 57568 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or2_1_inst_A2
timestamp 1698431365
transform 1 0 57120 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or2_2_inst_A1
timestamp 1698431365
transform 1 0 37520 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or2_2_inst_A2
timestamp 1698431365
transform 1 0 37296 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or2_4_inst_A1
timestamp 1698431365
transform 1 0 57120 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or2_4_inst_A2
timestamp 1698431365
transform 1 0 56672 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_1_inst_A1
timestamp 1698431365
transform 1 0 16576 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_1_inst_A2
timestamp 1698431365
transform 1 0 17024 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_1_inst_A3
timestamp 1698431365
transform 1 0 17472 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_2_inst_A1
timestamp 1698431365
transform 1 0 43904 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_2_inst_A2
timestamp 1698431365
transform 1 0 43008 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_2_inst_A3
timestamp 1698431365
transform 1 0 43456 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_4_inst_A1
timestamp 1698431365
transform 1 0 36848 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_4_inst_A2
timestamp 1698431365
transform 1 0 36400 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or3_4_inst_A3
timestamp 1698431365
transform 1 0 36400 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_1_inst_A1
timestamp 1698431365
transform 1 0 50848 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_1_inst_A2
timestamp 1698431365
transform 1 0 50400 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_1_inst_A3
timestamp 1698431365
transform 1 0 51072 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_1_inst_A4
timestamp 1698431365
transform 1 0 50624 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_2_inst_A1
timestamp 1698431365
transform 1 0 37968 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_2_inst_A2
timestamp 1698431365
transform 1 0 37520 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_2_inst_A3
timestamp 1698431365
transform 1 0 37072 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_2_inst_A4
timestamp 1698431365
transform 1 0 36960 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_4_inst_A1
timestamp 1698431365
transform 1 0 49504 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_4_inst_A2
timestamp 1698431365
transform 1 0 49952 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_4_inst_A3
timestamp 1698431365
transform 1 0 50624 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.or4_4_inst_A4
timestamp 1698431365
transform 1 0 50176 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_1_inst_CLK
timestamp 1698431365
transform 1 0 27776 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_1_inst_D
timestamp 1698431365
transform 1 0 22288 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_1_inst_SE
timestamp 1698431365
transform 1 0 21840 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_1_inst_SI
timestamp 1698431365
transform 1 0 21392 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_2_inst_CLK
timestamp 1698431365
transform 1 0 26320 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_2_inst_D
timestamp 1698431365
transform 1 0 20496 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_2_inst_SE
timestamp 1698431365
transform 1 0 20048 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_2_inst_SI
timestamp 1698431365
transform 1 0 25872 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_4_inst_CLK
timestamp 1698431365
transform 1 0 30688 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_4_inst_D
timestamp 1698431365
transform 1 0 25312 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_4_inst_SE
timestamp 1698431365
transform 1 0 24640 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffq_4_inst_SI
timestamp 1698431365
transform 1 0 24192 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_CLK
timestamp 1698431365
transform 1 0 31136 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_D
timestamp 1698431365
transform 1 0 30688 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_RN
timestamp 1698431365
transform 1 0 30240 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_SE
timestamp 1698431365
transform 1 0 29792 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_SI
timestamp 1698431365
transform 1 0 30240 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_CLK
timestamp 1698431365
transform 1 0 34048 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_D
timestamp 1698431365
transform 1 0 33600 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_RN
timestamp 1698431365
transform 1 0 32032 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_SE
timestamp 1698431365
transform 1 0 33152 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_SI
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_CLK
timestamp 1698431365
transform 1 0 39200 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_D
timestamp 1698431365
transform 1 0 38752 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_RN
timestamp 1698431365
transform 1 0 38976 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_SE
timestamp 1698431365
transform 1 0 38528 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_SI
timestamp 1698431365
transform 1 0 38080 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_CLK
timestamp 1698431365
transform 1 0 37072 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_D
timestamp 1698431365
transform 1 0 37968 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_RN
timestamp 1698431365
transform 1 0 37520 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SE
timestamp 1698431365
transform 1 0 37072 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SETN
timestamp 1698431365
transform -1 0 36848 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SI
timestamp 1698431365
transform 1 0 37072 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_CLK
timestamp 1698431365
transform 1 0 40320 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_D
timestamp 1698431365
transform 1 0 37632 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_RN
timestamp 1698431365
transform 1 0 37296 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 38192 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SE
timestamp 1698431365
transform 1 0 38640 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SI
timestamp 1698431365
transform 1 0 37744 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_CLK
timestamp 1698431365
transform 1 0 30240 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_D
timestamp 1698431365
transform 1 0 29792 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_RN
timestamp 1698431365
transform 1 0 29344 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SE
timestamp 1698431365
transform 1 0 30016 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 29344 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SI
timestamp 1698431365
transform -1 0 29456 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_CLK
timestamp 1698431365
transform 1 0 23968 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_D
timestamp 1698431365
transform 1 0 24640 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SETN
timestamp 1698431365
transform 1 0 25312 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SE
timestamp 1698431365
transform 1 0 23296 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SI
timestamp 1698431365
transform 1 0 24640 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_CLK
timestamp 1698431365
transform 1 0 31136 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_D
timestamp 1698431365
transform 1 0 20720 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SE
timestamp 1698431365
transform 1 0 20272 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 19824 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SI
timestamp 1698431365
transform 1 0 19376 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_CLK
timestamp 1698431365
transform 1 0 28560 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_D
timestamp 1698431365
transform 1 0 28112 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 29120 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SE
timestamp 1698431365
transform 1 0 28672 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SI
timestamp 1698431365
transform 1 0 28224 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor2_1_inst_A1
timestamp 1698431365
transform 1 0 35616 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor2_1_inst_A2
timestamp 1698431365
transform 1 0 35168 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor2_2_inst_A1
timestamp 1698431365
transform 1 0 56224 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor2_2_inst_A2
timestamp 1698431365
transform 1 0 55776 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor2_4_inst_A1
timestamp 1698431365
transform 1 0 18592 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor2_4_inst_A2
timestamp 1698431365
transform 1 0 16800 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_1_inst_A1
timestamp 1698431365
transform 1 0 44912 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_1_inst_A2
timestamp 1698431365
transform 1 0 43904 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_1_inst_A3
timestamp 1698431365
transform 1 0 44016 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_2_inst_A1
timestamp 1698431365
transform 1 0 36624 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_2_inst_A2
timestamp 1698431365
transform 1 0 35728 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_2_inst_A3
timestamp 1698431365
transform 1 0 36176 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_4_inst_A1
timestamp 1698431365
transform 1 0 53648 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_4_inst_A2
timestamp 1698431365
transform 1 0 51744 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xnor3_4_inst_A3
timestamp 1698431365
transform 1 0 51296 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor2_1_inst_A1
timestamp 1698431365
transform 1 0 38976 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor2_1_inst_A2
timestamp 1698431365
transform 1 0 38528 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor2_2_inst_A1
timestamp 1698431365
transform 1 0 53200 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor2_2_inst_A2
timestamp 1698431365
transform 1 0 52752 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor2_4_inst_A1
timestamp 1698431365
transform 1 0 30800 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor2_4_inst_A2
timestamp 1698431365
transform 1 0 31248 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_1_inst_A1
timestamp 1698431365
transform 1 0 55328 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_1_inst_A2
timestamp 1698431365
transform 1 0 56000 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_1_inst_A3
timestamp 1698431365
transform 1 0 54880 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_2_inst_A1
timestamp 1698431365
transform 1 0 27776 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_2_inst_A2
timestamp 1698431365
transform 1 0 23744 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_2_inst_A3
timestamp 1698431365
transform 1 0 23296 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_4_inst_A1
timestamp 1698431365
transform 1 0 56672 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_4_inst_A2
timestamp 1698431365
transform 1 0 56672 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_cm_inst.cc_inst.xor3_4_inst_A3
timestamp 1698431365
transform 1 0 49952 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[1\].div_flop_RN
timestamp 1698431365
transform 1 0 10416 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[2\].div_flop_RN
timestamp 1698431365
transform 1 0 8512 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[3\].div_flop_RN
timestamp 1698431365
transform 1 0 9296 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[4\].div_flop_RN
timestamp 1698431365
transform 1 0 9296 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[5\].div_flop_RN
timestamp 1698431365
transform 1 0 8960 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[6\].div_flop_RN
timestamp 1698431365
transform 1 0 2912 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[7\].div_flop_RN
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[8\].div_flop_RN
timestamp 1698431365
transform 1 0 5712 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[9\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[10\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[11\].div_flop_RN
timestamp 1698431365
transform 1 0 2352 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[12\].div_flop_RN
timestamp 1698431365
transform 1 0 2352 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[13\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[14\].div_flop_RN
timestamp 1698431365
transform 1 0 2688 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[15\].div_flop_RN
timestamp 1698431365
transform 1 0 3136 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[16\].div_flop_RN
timestamp 1698431365
transform 1 0 3808 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[17\].div_flop_RN
timestamp 1698431365
transform 1 0 4032 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[18\].div_flop_RN
timestamp 1698431365
transform 1 0 4592 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[19\].div_flop_RN
timestamp 1698431365
transform 1 0 3024 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[20\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[21\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[22\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[23\].div_flop_RN
timestamp 1698431365
transform 1 0 1792 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[24\].div_flop_RN
timestamp 1698431365
transform 1 0 3024 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[25\].div_flop_RN
timestamp 1698431365
transform 1 0 4144 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[26\].div_flop_RN
timestamp 1698431365
transform 1 0 6608 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[27\].div_flop_RN
timestamp 1698431365
transform 1 0 6160 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[28\].div_flop_RN
timestamp 1698431365
transform 1 0 9632 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[29\].div_flop_RN
timestamp 1698431365
transform 1 0 9296 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[30\].div_flop_RN
timestamp 1698431365
transform 1 0 9856 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[31\].div_flop_RN
timestamp 1698431365
transform 1 0 10416 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[32\].div_flop_RN
timestamp 1698431365
transform 1 0 9296 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[33\].div_flop_RN
timestamp 1698431365
transform 1 0 10416 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.gcount\[34\].div_flop_RN
timestamp 1698431365
transform 1 0 11312 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA_ro_inst.slow_clock_inv_I
timestamp 1698431365
transform 1 0 8512 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__addf_1  cm_inst.cc_inst.addf_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 36288
box -86 -90 3446 1098
use gf180mcu_fd_sc_mcu9t5v0__addf_2  cm_inst.cc_inst.addf_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 45808 0 1 32256
box -86 -90 3894 1098
use gf180mcu_fd_sc_mcu9t5v0__addf_4  cm_inst.cc_inst.addf_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 45696 0 1 28224
box -86 -90 4790 1098
use gf180mcu_fd_sc_mcu9t5v0__addh_1  cm_inst.cc_inst.addh_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 48384 0 -1 20160
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__addh_2  cm_inst.cc_inst.addh_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 40096 0 -1 36288
box -86 -90 2438 1098
use gf180mcu_fd_sc_mcu9t5v0__addh_4  cm_inst.cc_inst.addh_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 48944 0 1 34272
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_1  cm_inst.cc_inst.and2_1_inst
timestamp 1698431365
transform 1 0 31360 0 1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_2  cm_inst.cc_inst.and2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 51072 0 -1 34272
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__and2_4  cm_inst.cc_inst.and2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 26208
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__and3_1  cm_inst.cc_inst.and3_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 48608 0 -1 24192
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__and3_2  cm_inst.cc_inst.and3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 32256 0 1 26208
box -86 -90 1318 1098
use gf180mcu_fd_sc_mcu9t5v0__and3_4  cm_inst.cc_inst.and3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 50064 0 1 18144
box -86 -90 2326 1098
use gf180mcu_fd_sc_mcu9t5v0__and4_1  cm_inst.cc_inst.and4_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 18928 0 1 18144
box -86 -90 1318 1098
use gf180mcu_fd_sc_mcu9t5v0__and4_2  cm_inst.cc_inst.and4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 49168 0 -1 42336
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__and4_4  cm_inst.cc_inst.and4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 32592 0 1 24192
box -86 -90 2774 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_1  cm_inst.cc_inst.aoi21_1_inst
timestamp 1698431365
transform 1 0 25088 0 -1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_2  cm_inst.cc_inst.aoi21_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 57904 0 -1 34272
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi21_4  cm_inst.cc_inst.aoi21_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 23184 0 1 22176
box -86 -90 2774 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_1  cm_inst.cc_inst.aoi22_1_inst
timestamp 1698431365
transform -1 0 57456 0 -1 28224
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_2  cm_inst.cc_inst.aoi22_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 26880 0 -1 24192
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi22_4  cm_inst.cc_inst.aoi22_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 54880 0 -1 16128
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_1  cm_inst.cc_inst.aoi211_1_inst
timestamp 1698431365
transform -1 0 26208 0 -1 16128
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_2  cm_inst.cc_inst.aoi211_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 54208 0 -1 40320
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi211_4  cm_inst.cc_inst.aoi211_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 24080 0 -1 22176
box -86 -90 4118 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi221_1  cm_inst.cc_inst.aoi221_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 57456 0 1 32256
box -86 -90 1318 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi221_2  cm_inst.cc_inst.aoi221_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 22512 0 -1 24192
box -86 -90 2438 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi221_4  cm_inst.cc_inst.aoi221_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 57680 0 1 26208
box -86 -90 4566 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi222_1  cm_inst.cc_inst.aoi222_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 23296 0 1 24192
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi222_2  cm_inst.cc_inst.aoi222_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 52528 0 1 16128
box -86 -90 2886 1098
use gf180mcu_fd_sc_mcu9t5v0__aoi222_4  cm_inst.cc_inst.aoi222_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 26432 0 1 14112
box -86 -90 5350 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  cm_inst.cc_inst.buf_1_inst
timestamp 1698431365
transform -1 0 36064 0 -1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_2  cm_inst.cc_inst.buf_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 56112 0 -1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_3  cm_inst.cc_inst.buf_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 33376 0 1 34272
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_4  cm_inst.cc_inst.buf_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 50736 0 1 20160
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_8  cm_inst.cc_inst.buf_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 35840 0 -1 38304
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_12  cm_inst.cc_inst.buf_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 58128 0 1 18144
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_16  cm_inst.cc_inst.buf_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 14000 0 1 16128
box -86 -90 5686 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_20  cm_inst.cc_inst.buf_20_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 55552 0 -1 44352
box -86 -90 7030 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_1  cm_inst.cc_inst.bufz_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 39984 0 1 14112
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_2  cm_inst.cc_inst.bufz_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -90 1766 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_3  cm_inst.cc_inst.bufz_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 34496 0 1 14112
box -86 -90 2214 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_4  cm_inst.cc_inst.bufz_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 46032 0 -1 14112
box -86 -90 2438 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_8  cm_inst.cc_inst.bufz_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 48384 0 -1 12096
box -86 -90 3782 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_12  cm_inst.cc_inst.bufz_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 50288 0 1 12096
box -86 -90 5126 1098
use gf180mcu_fd_sc_mcu9t5v0__bufz_16  cm_inst.cc_inst.bufz_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 48384 0 -1 46368
box -86 -90 6470 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_1  cm_inst.cc_inst.clkbuf_1_inst
timestamp 1698431365
transform 1 0 40880 0 -1 14112
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_2  cm_inst.cc_inst.clkbuf_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_3  cm_inst.cc_inst.clkbuf_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 41104 0 -1 18144
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_4  cm_inst.cc_inst.clkbuf_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 40320
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_8  cm_inst.cc_inst.clkbuf_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 20160
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_12  cm_inst.cc_inst.clkbuf_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 45808 0 -1 26208
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_16  cm_inst.cc_inst.clkbuf_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 24192
box -86 -90 5686 1098
use gf180mcu_fd_sc_mcu9t5v0__clkbuf_20  cm_inst.cc_inst.clkbuf_20_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 10080 0 -1 24192
box -86 -90 7030 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_1  cm_inst.cc_inst.clkinv_1_inst
timestamp 1698431365
transform -1 0 23184 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_2  cm_inst.cc_inst.clkinv_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 -1 40320
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_3  cm_inst.cc_inst.clkinv_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_4  cm_inst.cc_inst.clkinv_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 27328 0 1 40320
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_8  cm_inst.cc_inst.clkinv_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 20048 0 1 20160
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_12  cm_inst.cc_inst.clkinv_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 42000 0 -1 28224
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_16  cm_inst.cc_inst.clkinv_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 17360 0 1 22176
box -86 -90 3894 1098
use gf180mcu_fd_sc_mcu9t5v0__clkinv_20  cm_inst.cc_inst.clkinv_20_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 26208
box -86 -90 4790 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnq_1  cm_inst.cc_inst.dffnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 25760 0 -1 48384
box -86 -90 3446 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnq_2  cm_inst.cc_inst.dffnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17472 0 1 12096
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnq_4  cm_inst.cc_inst.dffnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 6048
box -86 -90 4006 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1  cm_inst.cc_inst.dffnrnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 39424 0 1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2  cm_inst.cc_inst.dffnrnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 20160
box -86 -90 4006 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4  cm_inst.cc_inst.dffnrnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 40096 0 1 46368
box -86 -90 4454 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1  cm_inst.cc_inst.dffnrsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29680 0 1 44352
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2  cm_inst.cc_inst.dffnrsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 38080 0 1 44352
box -86 -90 4566 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4  cm_inst.cc_inst.dffnrsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 23296 0 1 44352
box -86 -90 5014 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1  cm_inst.cc_inst.dffnsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 1 10080
box -86 -90 4118 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2  cm_inst.cc_inst.dffnsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 6048
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4  cm_inst.cc_inst.dffnsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 35840 0 -1 10080
box -86 -90 4790 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_1  cm_inst.cc_inst.dffq_1_inst
timestamp 1698431365
transform 1 0 37408 0 1 20160
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_2  cm_inst.cc_inst.dffq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 37184 0 1 48384
box -86 -90 3446 1098
use gf180mcu_fd_sc_mcu9t5v0__dffq_4  cm_inst.cc_inst.dffq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 27888 0 -1 44352
box -86 -90 4006 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  cm_inst.cc_inst.dffrnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 36064 0 -1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_2  cm_inst.cc_inst.dffrnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 1 46368
box -86 -90 3894 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_4  cm_inst.cc_inst.dffrnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 12096
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1  cm_inst.cc_inst.dffrsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 28560 0 -1 6048
box -86 -90 4230 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2  cm_inst.cc_inst.dffrsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 37072 0 1 8064
box -86 -90 4454 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4  cm_inst.cc_inst.dffrsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 35728 0 -1 20160
box -86 -90 4902 1098
use gf180mcu_fd_sc_mcu9t5v0__dffsnq_1  cm_inst.cc_inst.dffsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 36512 0 -1 48384
box -86 -90 4118 1098
use gf180mcu_fd_sc_mcu9t5v0__dffsnq_2  cm_inst.cc_inst.dffsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 28000 0 -1 46368
box -86 -90 4230 1098
use gf180mcu_fd_sc_mcu9t5v0__dffsnq_4  cm_inst.cc_inst.dffsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 35728 0 -1 46368
box -86 -90 4790 1098
use gf180mcu_fd_sc_mcu9t5v0__dlya_1  cm_inst.cc_inst.dlya_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 22400 0 1 8064
box -86 -90 1318 1098
use gf180mcu_fd_sc_mcu9t5v0__dlya_2  cm_inst.cc_inst.dlya_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 24864 0 1 10080
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__dlya_4  cm_inst.cc_inst.dlya_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 30800 0 -1 12096
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyb_1  cm_inst.cc_inst.dlyb_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 33712 0 1 16128
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyb_2  cm_inst.cc_inst.dlyb_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 40432 0 1 14112
box -86 -90 1766 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyb_4  cm_inst.cc_inst.dlyb_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 38192 0 -1 40320
box -86 -90 2214 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyc_1  cm_inst.cc_inst.dlyc_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 38304 0 -1 18144
box -86 -90 2326 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyc_2  cm_inst.cc_inst.dlyc_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 30240 0 -1 40320
box -86 -90 2550 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyc_4  cm_inst.cc_inst.dlyc_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 18032 0 1 6048
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyd_1  cm_inst.cc_inst.dlyd_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 28672 0 1 6048
box -86 -90 3110 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyd_2  cm_inst.cc_inst.dlyd_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29456 0 -1 10080
box -86 -90 3334 1098
use gf180mcu_fd_sc_mcu9t5v0__dlyd_4  cm_inst.cc_inst.dlyd_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 16128
box -86 -90 3782 1098
use gf180mcu_fd_sc_mcu9t5v0__hold  cm_inst.cc_inst.hold_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 45696 0 -1 44352
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__icgtn_1  cm_inst.cc_inst.icgtn_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 1 26208
box -86 -90 3446 1098
use gf180mcu_fd_sc_mcu9t5v0__icgtn_2  cm_inst.cc_inst.icgtn_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 23744 0 1 40320
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__icgtn_4  cm_inst.cc_inst.icgtn_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -90 4118 1098
use gf180mcu_fd_sc_mcu9t5v0__icgtp_1  cm_inst.cc_inst.icgtp_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 40320
box -86 -90 3110 1098
use gf180mcu_fd_sc_mcu9t5v0__icgtp_2  cm_inst.cc_inst.icgtp_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 19040 0 -1 24192
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__icgtp_4  cm_inst.cc_inst.icgtp_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 27440 0 -1 24192
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  cm_inst.cc_inst.inv_1_inst
timestamp 1698431365
transform 1 0 32256 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_2  cm_inst.cc_inst.inv_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 56224 0 -1 34272
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_3  cm_inst.cc_inst.inv_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 35392 0 -1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_4  cm_inst.cc_inst.inv_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 51744 0 -1 20160
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_8  cm_inst.cc_inst.inv_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 32368 0 1 36288
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_12  cm_inst.cc_inst.inv_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 53312 0 -1 18144
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_16  cm_inst.cc_inst.inv_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 19376 0 1 14112
box -86 -90 3894 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_20  cm_inst.cc_inst.inv_20_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 47376 0 1 40320
box -86 -90 4790 1098
use gf180mcu_fd_sc_mcu9t5v0__invz_1  cm_inst.cc_inst.invz_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 45584 0 1 44352
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__invz_2  cm_inst.cc_inst.invz_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 16128
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__invz_3  cm_inst.cc_inst.invz_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 47264 0 -1 16128
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__invz_4  cm_inst.cc_inst.invz_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 47040 0 -1 18144
box -86 -90 2774 1098
use gf180mcu_fd_sc_mcu9t5v0__invz_8  cm_inst.cc_inst.invz_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 31696 0 1 48384
box -86 -90 4230 1098
use gf180mcu_fd_sc_mcu9t5v0__invz_12  cm_inst.cc_inst.invz_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 30352 0 1 46368
box -86 -90 5910 1098
use gf180mcu_fd_sc_mcu9t5v0__latq_1  cm_inst.cc_inst.latq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 46928 0 1 36288
box -86 -90 2326 1098
use gf180mcu_fd_sc_mcu9t5v0__latq_2  cm_inst.cc_inst.latq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 41440 0 1 34272
box -86 -90 2550 1098
use gf180mcu_fd_sc_mcu9t5v0__latq_4  cm_inst.cc_inst.latq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 49168 0 1 30240
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__latrnq_1  cm_inst.cc_inst.latrnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 1 30240
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__latrnq_2  cm_inst.cc_inst.latrnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 44800 0 -1 22176
box -86 -90 2886 1098
use gf180mcu_fd_sc_mcu9t5v0__latrnq_4  cm_inst.cc_inst.latrnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 19152 0 -1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__latrsnq_1  cm_inst.cc_inst.latrsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 33264 0 1 6048
box -86 -90 2774 1098
use gf180mcu_fd_sc_mcu9t5v0__latrsnq_2  cm_inst.cc_inst.latrsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 41440 0 1 8064
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__latrsnq_4  cm_inst.cc_inst.latrsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 40992 0 1 20160
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__latsnq_1  cm_inst.cc_inst.latsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 42000 0 1 48384
box -86 -90 2438 1098
use gf180mcu_fd_sc_mcu9t5v0__latsnq_2  cm_inst.cc_inst.latsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 44352
box -86 -90 2550 1098
use gf180mcu_fd_sc_mcu9t5v0__latsnq_4  cm_inst.cc_inst.latsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 44240 0 -1 48384
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_1  cm_inst.cc_inst.mux2_1_inst
timestamp 1698431365
transform 1 0 52528 0 1 30240
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_2  cm_inst.cc_inst.mux2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 42224 0 -1 32256
box -86 -90 1766 1098
use gf180mcu_fd_sc_mcu9t5v0__mux2_4  cm_inst.cc_inst.mux2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 45920 0 -1 24192
box -86 -90 2214 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_1  cm_inst.cc_inst.mux4_1_inst
timestamp 1698431365
transform 1 0 29008 0 1 16128
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_2  cm_inst.cc_inst.mux4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 43232 0 1 38304
box -86 -90 3894 1098
use gf180mcu_fd_sc_mcu9t5v0__mux4_4  cm_inst.cc_inst.mux4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 36960 0 1 34272
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  cm_inst.cc_inst.nand2_1_inst
timestamp 1698431365
transform 1 0 52640 0 1 34272
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_2  cm_inst.cc_inst.nand2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 35840 0 -1 26208
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_4  cm_inst.cc_inst.nand2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 48832 0 -1 20160
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__nand3_1  cm_inst.cc_inst.nand3_1_inst
timestamp 1698431365
transform 1 0 31024 0 -1 26208
box -86 -90 870 1098
use gf180mcu_fd_sc_mcu9t5v0__nand3_2  cm_inst.cc_inst.nand3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 50064 0 1 18144
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__nand3_4  cm_inst.cc_inst.nand3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 -1 20160
box -86 -90 2886 1098
use gf180mcu_fd_sc_mcu9t5v0__nand4_1  cm_inst.cc_inst.nand4_1_inst
timestamp 1698431365
transform 1 0 47376 0 1 42336
box -86 -90 1094 1098
use gf180mcu_fd_sc_mcu9t5v0__nand4_2  cm_inst.cc_inst.nand4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 24192
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__nand4_4  cm_inst.cc_inst.nand4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 57792 0 1 34272
box -86 -90 3558 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_1  cm_inst.cc_inst.nor2_1_inst
timestamp 1698431365
transform 1 0 40880 0 -1 26208
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_2  cm_inst.cc_inst.nor2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 57568 0 1 24192
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__nor2_4  cm_inst.cc_inst.nor2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 38304 0 1 30240
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__nor3_1  cm_inst.cc_inst.nor3_1_inst
timestamp 1698431365
transform -1 0 57904 0 1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__nor3_2  cm_inst.cc_inst.nor3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 16128
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__nor3_4  cm_inst.cc_inst.nor3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 45472 0 -1 42336
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__nor4_1  cm_inst.cc_inst.nor4_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 41104 0 1 22176
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__nor4_2  cm_inst.cc_inst.nor4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 58352 0 1 36288
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__nor4_4  cm_inst.cc_inst.nor4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 43792 0 1 24192
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_1  cm_inst.cc_inst.oai21_1_inst
timestamp 1698431365
transform 1 0 52864 0 -1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_2  cm_inst.cc_inst.oai21_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 32592 0 -1 24192
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__oai21_4  cm_inst.cc_inst.oai21_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 52640 0 -1 32256
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__oai22_1  cm_inst.cc_inst.oai22_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 30576 0 1 22176
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__oai22_2  cm_inst.cc_inst.oai22_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 49952 0 -1 28224
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__oai22_4  cm_inst.cc_inst.oai22_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 27776 0 -1 22176
box -86 -90 3894 1098
use gf180mcu_fd_sc_mcu9t5v0__oai31_1  cm_inst.cc_inst.oai31_1_inst
timestamp 1698431365
transform 1 0 47264 0 -1 18144
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__oai31_2  cm_inst.cc_inst.oai31_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 22848 0 -1 16128
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__oai31_4  cm_inst.cc_inst.oai31_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 56448 0 1 40320
box -86 -90 4006 1098
use gf180mcu_fd_sc_mcu9t5v0__oai32_1  cm_inst.cc_inst.oai32_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 31024 0 1 20160
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__oai32_2  cm_inst.cc_inst.oai32_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 55216 0 -1 36288
box -86 -90 2550 1098
use gf180mcu_fd_sc_mcu9t5v0__oai32_4  cm_inst.cc_inst.oai32_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29792 0 1 18144
box -86 -90 4902 1098
use gf180mcu_fd_sc_mcu9t5v0__oai33_1  cm_inst.cc_inst.oai33_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 50624 0 1 26208
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__oai33_2  cm_inst.cc_inst.oai33_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29120 0 -1 20160
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__oai33_4  cm_inst.cc_inst.oai33_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 46592 0 1 16128
box -86 -90 5798 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_1  cm_inst.cc_inst.oai211_1_inst
timestamp 1698431365
transform -1 0 31024 0 1 14112
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_2  cm_inst.cc_inst.oai211_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 44352 0 1 36288
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__oai211_4  cm_inst.cc_inst.oai211_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 39424 0 1 32256
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__oai221_1  cm_inst.cc_inst.oai221_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 49504 0 1 36288
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__oai221_2  cm_inst.cc_inst.oai221_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 47040 0 -1 32256
box -86 -90 2550 1098
use gf180mcu_fd_sc_mcu9t5v0__oai221_4  cm_inst.cc_inst.oai221_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 57792 0 1 28224
box -86 -90 4902 1098
use gf180mcu_fd_sc_mcu9t5v0__oai222_1  cm_inst.cc_inst.oai222_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 46368 0 1 30240
box -86 -90 1766 1098
use gf180mcu_fd_sc_mcu9t5v0__oai222_2  cm_inst.cc_inst.oai222_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 47264 0 1 20160
box -86 -90 3110 1098
use gf180mcu_fd_sc_mcu9t5v0__oai222_4  cm_inst.cc_inst.oai222_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 -1 16128
box -86 -90 5798 1098
use gf180mcu_fd_sc_mcu9t5v0__or2_1  cm_inst.cc_inst.or2_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 55776 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__or2_2  cm_inst.cc_inst.or2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 37744 0 1 32256
box -86 -90 1206 1098
use gf180mcu_fd_sc_mcu9t5v0__or2_4  cm_inst.cc_inst.or2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 54208 0 -1 24192
box -86 -90 2102 1098
use gf180mcu_fd_sc_mcu9t5v0__or3_1  cm_inst.cc_inst.or3_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17696 0 1 18144
box -86 -90 1318 1098
use gf180mcu_fd_sc_mcu9t5v0__or3_2  cm_inst.cc_inst.or3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 44128 0 -1 42336
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__or3_4  cm_inst.cc_inst.or3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 39312 0 1 24192
box -86 -90 2550 1098
use gf180mcu_fd_sc_mcu9t5v0__or4_1  cm_inst.cc_inst.or4_1_inst
timestamp 1698431365
transform 1 0 50848 0 1 36288
box -86 -90 1542 1098
use gf180mcu_fd_sc_mcu9t5v0__or4_2  cm_inst.cc_inst.or4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 37408 0 -1 26208
box -86 -90 1654 1098
use gf180mcu_fd_sc_mcu9t5v0__or4_4  cm_inst.cc_inst.or4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 50960 0 -1 24192
box -86 -90 2998 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffq_1  cm_inst.cc_inst.sdffq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 22512 0 1 42336
box -86 -90 4342 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffq_2  cm_inst.cc_inst.sdffq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 6048
box -86 -90 4566 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffq_4  cm_inst.cc_inst.sdffq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 8064
box -86 -90 5014 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1  cm_inst.cc_inst.sdffrnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 31360 0 1 8064
box -86 -90 4678 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2  cm_inst.cc_inst.sdffrnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 33600 0 -1 14112
box -86 -90 4790 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4  cm_inst.cc_inst.sdffrnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 39200 0 1 12096
box -86 -90 5350 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1  cm_inst.cc_inst.sdffrsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 37296 0 1 40320
box -86 -90 5238 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2  cm_inst.cc_inst.sdffrsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 39088 0 1 16128
box -86 -90 5462 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4  cm_inst.cc_inst.sdffrsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 30464 0 1 40320
box -86 -90 5910 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1  cm_inst.cc_inst.sdffsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 19264 0 -1 8064
box -86 -90 5014 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2  cm_inst.cc_inst.sdffsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 23520 0 1 8064
box -86 -90 5126 1098
use gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4  cm_inst.cc_inst.sdffsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 29344 0 1 10080
box -86 -90 5574 1098
use gf180mcu_fd_sc_mcu9t5v0__tieh  cm_inst.cc_inst.tieh_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 20496 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__tiel  cm_inst.cc_inst.tiel_inst
timestamp 1698431365
transform -1 0 52640 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor2_1  cm_inst.cc_inst.xnor2_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 35280 0 1 30240
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor2_2  cm_inst.cc_inst.xnor2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 52752 0 1 20160
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor2_4  cm_inst.cc_inst.xnor2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 18144
box -86 -90 2438 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor3_1  cm_inst.cc_inst.xnor3_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 47264 0 1 40320
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor3_2  cm_inst.cc_inst.xnor3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 39984 0 1 22176
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor3_4  cm_inst.cc_inst.xnor3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 51744 0 -1 38304
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__xor2_1  cm_inst.cc_inst.xor2_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 40320 0 -1 26208
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__xor2_2  cm_inst.cc_inst.xor2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 54880 0 -1 26208
box -86 -90 1990 1098
use gf180mcu_fd_sc_mcu9t5v0__xor2_4  cm_inst.cc_inst.xor2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 33824 0 -1 32256
box -86 -90 2438 1098
use gf180mcu_fd_sc_mcu9t5v0__xor3_1  cm_inst.cc_inst.xor3_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 55776 0 -1 22176
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__xor3_2  cm_inst.cc_inst.xor3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 23968 0 1 12096
box -86 -90 3222 1098
use gf180mcu_fd_sc_mcu9t5v0__xor3_4  cm_inst.cc_inst.xor3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 57456 0 1 38304
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_0_172 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 20608 0 1 4032
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_0_188 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 22400 0 1 4032
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_0_196 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 23296 0 1 4032
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_0_200 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 23744 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_0_210
timestamp 1698431365
transform 1 0 24864 0 1 4032
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_0_214 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 25312 0 1 4032
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_0_217
timestamp 1698431365
transform 1 0 25648 0 1 4032
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_0_233
timestamp 1698431365
transform 1 0 27440 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 4032
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_0_244
timestamp 1698431365
transform 1 0 28672 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_0_248
timestamp 1698431365
transform 1 0 29120 0 1 4032
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_0_264
timestamp 1698431365
transform 1 0 30912 0 1 4032
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_0_276
timestamp 1698431365
transform 1 0 32256 0 1 4032
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_0_279
timestamp 1698431365
transform 1 0 32592 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_0_283
timestamp 1698431365
transform 1 0 33040 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_0_287
timestamp 1698431365
transform 1 0 33488 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_0_291
timestamp 1698431365
transform 1 0 33936 0 1 4032
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_0_299
timestamp 1698431365
transform 1 0 34832 0 1 4032
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_0_303
timestamp 1698431365
transform 1 0 35280 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 4032
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 4032
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_0_494
timestamp 1698431365
transform 1 0 56672 0 1 4032
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_0_502
timestamp 1698431365
transform 1 0 57568 0 1 4032
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_0_506
timestamp 1698431365
transform 1 0 58016 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_0_508
timestamp 1698431365
transform 1 0 58240 0 1 4032
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 6048
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_1_158
timestamp 1698431365
transform 1 0 19040 0 -1 6048
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_1_166
timestamp 1698431365
transform 1 0 19936 0 -1 6048
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_1_169
timestamp 1698431365
transform 1 0 20272 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_1_173
timestamp 1698431365
transform 1 0 20720 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_1_177
timestamp 1698431365
transform 1 0 21168 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_1_216
timestamp 1698431365
transform 1 0 25536 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_1_218
timestamp 1698431365
transform 1 0 25760 0 -1 6048
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_1_221
timestamp 1698431365
transform 1 0 26096 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_225
timestamp 1698431365
transform 1 0 26544 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_1_231
timestamp 1698431365
transform 1 0 27216 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_1_235
timestamp 1698431365
transform 1 0 27664 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_1_239
timestamp 1698431365
transform 1 0 28112 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_1_317
timestamp 1698431365
transform 1 0 36848 0 -1 6048
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 6048
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698431365
transform 1 0 47936 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698431365
transform 1 0 55776 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 6048
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_1_508
timestamp 1698431365
transform 1 0 58240 0 -1 6048
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 6048
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_18
timestamp 1698431365
transform 1 0 3360 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_2_22
timestamp 1698431365
transform 1 0 3808 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_2_32
timestamp 1698431365
transform 1 0 4928 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 6048
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 6048
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_2_139
timestamp 1698431365
transform 1 0 16912 0 1 6048
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_2_147
timestamp 1698431365
transform 1 0 17808 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 6048
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_309
timestamp 1698431365
transform 1 0 35952 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_2_313
timestamp 1698431365
transform 1 0 36400 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_451
timestamp 1698431365
transform 1 0 51856 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 6048
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698431365
transform 1 0 56112 0 1 6048
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_505
timestamp 1698431365
transform 1 0 57904 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 8064
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_158
timestamp 1698431365
transform 1 0 19040 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_204
timestamp 1698431365
transform 1 0 24192 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_256
timestamp 1698431365
transform 1 0 30016 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_260
timestamp 1698431365
transform 1 0 30464 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_264
timestamp 1698431365
transform 1 0 30912 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_268
timestamp 1698431365
transform 1 0 31360 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_3_272
timestamp 1698431365
transform 1 0 31808 0 -1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_275
timestamp 1698431365
transform 1 0 32144 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_313
timestamp 1698431365
transform 1 0 36400 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_317
timestamp 1698431365
transform 1 0 36848 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_321
timestamp 1698431365
transform 1 0 37296 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_3_325
timestamp 1698431365
transform 1 0 37744 0 -1 8064
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_341
timestamp 1698431365
transform 1 0 39536 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_345
timestamp 1698431365
transform 1 0 39984 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_3_347
timestamp 1698431365
transform 1 0 40208 0 -1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_356
timestamp 1698431365
transform 1 0 41216 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_3_360
timestamp 1698431365
transform 1 0 41664 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_3_364
timestamp 1698431365
transform 1 0 42112 0 -1 8064
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_3_396
timestamp 1698431365
transform 1 0 45696 0 -1 8064
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_3_412
timestamp 1698431365
transform 1 0 47488 0 -1 8064
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698431365
transform 1 0 55776 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 8064
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_3_508
timestamp 1698431365
transform 1 0 58240 0 -1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 8064
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 8064
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_4_139
timestamp 1698431365
transform 1 0 16912 0 1 8064
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_155
timestamp 1698431365
transform 1 0 18704 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_159
timestamp 1698431365
transform 1 0 19152 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_163
timestamp 1698431365
transform 1 0 19600 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_167
timestamp 1698431365
transform 1 0 20048 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_188
timestamp 1698431365
transform 1 0 22400 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_4_190
timestamp 1698431365
transform 1 0 22624 0 1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_193
timestamp 1698431365
transform 1 0 22960 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_4_195
timestamp 1698431365
transform 1 0 23184 0 1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_243
timestamp 1698431365
transform 1 0 28560 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_251
timestamp 1698431365
transform 1 0 29456 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_4_253
timestamp 1698431365
transform 1 0 29680 0 1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_256
timestamp 1698431365
transform 1 0 30016 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_260
timestamp 1698431365
transform 1 0 30464 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_264
timestamp 1698431365
transform 1 0 30912 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_309
timestamp 1698431365
transform 1 0 35952 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_313
timestamp 1698431365
transform 1 0 36400 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_4_384
timestamp 1698431365
transform 1 0 44352 0 1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698431365
transform 1 0 51856 0 1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 8064
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_4_489
timestamp 1698431365
transform 1 0 56112 0 1 8064
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_4_505
timestamp 1698431365
transform 1 0 57904 0 1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 10080
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_150
timestamp 1698431365
transform 1 0 18144 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_5_152
timestamp 1698431365
transform 1 0 18368 0 -1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_155
timestamp 1698431365
transform 1 0 18704 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_191
timestamp 1698431365
transform 1 0 22736 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_197
timestamp 1698431365
transform 1 0 23408 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_201
timestamp 1698431365
transform 1 0 23856 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_5_203
timestamp 1698431365
transform 1 0 24080 0 -1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_249
timestamp 1698431365
transform 1 0 29232 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 10080
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_300
timestamp 1698431365
transform 1 0 34944 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_5_304
timestamp 1698431365
transform 1 0 35392 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_5_383
timestamp 1698431365
transform 1 0 44240 0 -1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_415
timestamp 1698431365
transform 1 0 47824 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_5_419
timestamp 1698431365
transform 1 0 48272 0 -1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 10080
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_5_508
timestamp 1698431365
transform 1 0 58240 0 -1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 10080
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_6_123
timestamp 1698431365
transform 1 0 15120 0 1 10080
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_6_131
timestamp 1698431365
transform 1 0 16016 0 1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_168
timestamp 1698431365
transform 1 0 20160 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_208
timestamp 1698431365
transform 1 0 24640 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_6_223
timestamp 1698431365
transform 1 0 26320 0 1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_237
timestamp 1698431365
transform 1 0 27888 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_6_249
timestamp 1698431365
transform 1 0 29232 0 1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_6_299
timestamp 1698431365
transform 1 0 34832 0 1 10080
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 10080
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_325
timestamp 1698431365
transform 1 0 37744 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_6_329
timestamp 1698431365
transform 1 0 38192 0 1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_332
timestamp 1698431365
transform 1 0 38528 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_336
timestamp 1698431365
transform 1 0 38976 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_6_372
timestamp 1698431365
transform 1 0 43008 0 1 10080
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_380
timestamp 1698431365
transform 1 0 43904 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_6_384
timestamp 1698431365
transform 1 0 44352 0 1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698431365
transform 1 0 51856 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_6_489
timestamp 1698431365
transform 1 0 56112 0 1 10080
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_505
timestamp 1698431365
transform 1 0 57904 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_180
timestamp 1698431365
transform 1 0 21504 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_186
timestamp 1698431365
transform 1 0 22176 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_190
timestamp 1698431365
transform 1 0 22624 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_207
timestamp 1698431365
transform 1 0 24528 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_216
timestamp 1698431365
transform 1 0 25536 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_220
timestamp 1698431365
transform 1 0 25984 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_222
timestamp 1698431365
transform 1 0 26208 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_7_225
timestamp 1698431365
transform 1 0 26544 0 -1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_233
timestamp 1698431365
transform 1 0 27440 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_235
timestamp 1698431365
transform 1 0 27664 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_238
timestamp 1698431365
transform 1 0 28000 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_242
timestamp 1698431365
transform 1 0 28448 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_246
timestamp 1698431365
transform 1 0 28896 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_7_250
timestamp 1698431365
transform 1 0 29344 0 -1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_258
timestamp 1698431365
transform 1 0 30240 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_260
timestamp 1698431365
transform 1 0 30464 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_7_313
timestamp 1698431365
transform 1 0 36400 0 -1 12096
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_329
timestamp 1698431365
transform 1 0 38192 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_333
timestamp 1698431365
transform 1 0 38640 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_336
timestamp 1698431365
transform 1 0 38976 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_7_340
timestamp 1698431365
transform 1 0 39424 0 -1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_348
timestamp 1698431365
transform 1 0 40320 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 12096
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_7_368
timestamp 1698431365
transform 1 0 42560 0 -1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_376
timestamp 1698431365
transform 1 0 43456 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_379
timestamp 1698431365
transform 1 0 43792 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_7_383
timestamp 1698431365
transform 1 0 44240 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698431365
transform 1 0 55776 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 12096
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_508
timestamp 1698431365
transform 1 0 58240 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 12096
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 12096
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_139
timestamp 1698431365
transform 1 0 16912 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_143
timestamp 1698431365
transform 1 0 17360 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_181
timestamp 1698431365
transform 1 0 21616 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_8_185
timestamp 1698431365
transform 1 0 22064 0 1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_193
timestamp 1698431365
transform 1 0 22960 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_195
timestamp 1698431365
transform 1 0 23184 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_198
timestamp 1698431365
transform 1 0 23520 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_230
timestamp 1698431365
transform 1 0 27104 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_234
timestamp 1698431365
transform 1 0 27552 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_238
timestamp 1698431365
transform 1 0 28000 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_242
timestamp 1698431365
transform 1 0 28448 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 12096
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_8_263
timestamp 1698431365
transform 1 0 30800 0 1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_271
timestamp 1698431365
transform 1 0 31696 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_286
timestamp 1698431365
transform 1 0 33376 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_290
timestamp 1698431365
transform 1 0 33824 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_294
timestamp 1698431365
transform 1 0 34272 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_8_298
timestamp 1698431365
transform 1 0 34720 0 1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_306
timestamp 1698431365
transform 1 0 35616 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_310
timestamp 1698431365
transform 1 0 36064 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_312
timestamp 1698431365
transform 1 0 36288 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_321
timestamp 1698431365
transform 1 0 37296 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_327
timestamp 1698431365
transform 1 0 37968 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_330
timestamp 1698431365
transform 1 0 38304 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_334
timestamp 1698431365
transform 1 0 38752 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_391
timestamp 1698431365
transform 1 0 45136 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_8_437
timestamp 1698431365
transform 1 0 50288 0 1 12096
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_453
timestamp 1698431365
transform 1 0 52080 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 12096
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_8_489
timestamp 1698431365
transform 1 0 56112 0 1 12096
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_505
timestamp 1698431365
transform 1 0 57904 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_158
timestamp 1698431365
transform 1 0 19040 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_160
timestamp 1698431365
transform 1 0 19264 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_9_163
timestamp 1698431365
transform 1 0 19600 0 -1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_173
timestamp 1698431365
transform 1 0 20720 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_177
timestamp 1698431365
transform 1 0 21168 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_181
timestamp 1698431365
transform 1 0 21616 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_189
timestamp 1698431365
transform 1 0 22512 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_193
timestamp 1698431365
transform 1 0 22960 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_197
timestamp 1698431365
transform 1 0 23408 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_201
timestamp 1698431365
transform 1 0 23856 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_203
timestamp 1698431365
transform 1 0 24080 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_214
timestamp 1698431365
transform 1 0 25312 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_217
timestamp 1698431365
transform 1 0 25648 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_221
timestamp 1698431365
transform 1 0 26096 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_225
timestamp 1698431365
transform 1 0 26544 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_229
timestamp 1698431365
transform 1 0 26992 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_233
timestamp 1698431365
transform 1 0 27440 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_237
timestamp 1698431365
transform 1 0 27888 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_241
timestamp 1698431365
transform 1 0 28336 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_247
timestamp 1698431365
transform 1 0 29008 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_251
timestamp 1698431365
transform 1 0 29456 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_255
timestamp 1698431365
transform 1 0 29904 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_9_259
timestamp 1698431365
transform 1 0 30352 0 -1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_267
timestamp 1698431365
transform 1 0 31248 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_271
timestamp 1698431365
transform 1 0 31696 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_273
timestamp 1698431365
transform 1 0 31920 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_286
timestamp 1698431365
transform 1 0 33376 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_330
timestamp 1698431365
transform 1 0 38304 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_334
timestamp 1698431365
transform 1 0 38752 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_9_338
timestamp 1698431365
transform 1 0 39200 0 -1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_390
timestamp 1698431365
transform 1 0 45024 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_394
timestamp 1698431365
transform 1 0 45472 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_397
timestamp 1698431365
transform 1 0 45808 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_438
timestamp 1698431365
transform 1 0 50400 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_442
timestamp 1698431365
transform 1 0 50848 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_444
timestamp 1698431365
transform 1 0 51072 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_9_447
timestamp 1698431365
transform 1 0 51408 0 -1 14112
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_9_479
timestamp 1698431365
transform 1 0 54992 0 -1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_9_487
timestamp 1698431365
transform 1 0 55888 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_489
timestamp 1698431365
transform 1 0 56112 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_123
timestamp 1698431365
transform 1 0 15120 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_161
timestamp 1698431365
transform 1 0 19376 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_167
timestamp 1698431365
transform 1 0 20048 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_230
timestamp 1698431365
transform 1 0 27104 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_10_234
timestamp 1698431365
transform 1 0 27552 0 1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_237
timestamp 1698431365
transform 1 0 27888 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_251
timestamp 1698431365
transform 1 0 29456 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_10_265
timestamp 1698431365
transform 1 0 31024 0 1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_273
timestamp 1698431365
transform 1 0 31920 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_10_275
timestamp 1698431365
transform 1 0 32144 0 1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_278
timestamp 1698431365
transform 1 0 32480 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_10_282
timestamp 1698431365
transform 1 0 32928 0 1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_289
timestamp 1698431365
transform 1 0 33712 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_10_291
timestamp 1698431365
transform 1 0 33936 0 1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_294
timestamp 1698431365
transform 1 0 34272 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_345
timestamp 1698431365
transform 1 0 39984 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_364
timestamp 1698431365
transform 1 0 42112 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_10_368
timestamp 1698431365
transform 1 0 42560 0 1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_376
timestamp 1698431365
transform 1 0 43456 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_10_378
timestamp 1698431365
transform 1 0 43680 0 1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_391
timestamp 1698431365
transform 1 0 45136 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_395
timestamp 1698431365
transform 1 0 45584 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_399
timestamp 1698431365
transform 1 0 46032 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_403
timestamp 1698431365
transform 1 0 46480 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_407
timestamp 1698431365
transform 1 0 46928 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_411
timestamp 1698431365
transform 1 0 47376 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_10_415
timestamp 1698431365
transform 1 0 47824 0 1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_423
timestamp 1698431365
transform 1 0 48720 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_429
timestamp 1698431365
transform 1 0 49392 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_433
timestamp 1698431365
transform 1 0 49840 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_437
timestamp 1698431365
transform 1 0 50288 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_441
timestamp 1698431365
transform 1 0 50736 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_445
timestamp 1698431365
transform 1 0 51184 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_451
timestamp 1698431365
transform 1 0 51856 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_461
timestamp 1698431365
transform 1 0 52976 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_10_465
timestamp 1698431365
transform 1 0 53424 0 1 14112
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_10_497
timestamp 1698431365
transform 1 0 57008 0 1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_505
timestamp 1698431365
transform 1 0 57904 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 16128
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_152
timestamp 1698431365
transform 1 0 18368 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_187
timestamp 1698431365
transform 1 0 22288 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_11_189
timestamp 1698431365
transform 1 0 22512 0 -1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_222
timestamp 1698431365
transform 1 0 26208 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_11_226
timestamp 1698431365
transform 1 0 26656 0 -1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_346
timestamp 1698431365
transform 1 0 40096 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_410
timestamp 1698431365
transform 1 0 47264 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_414
timestamp 1698431365
transform 1 0 47712 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_418
timestamp 1698431365
transform 1 0 48160 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_426
timestamp 1698431365
transform 1 0 49056 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_430
timestamp 1698431365
transform 1 0 49504 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_434
timestamp 1698431365
transform 1 0 49952 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_438
timestamp 1698431365
transform 1 0 50400 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_11_440
timestamp 1698431365
transform 1 0 50624 0 -1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_11_443
timestamp 1698431365
transform 1 0 50960 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_11_478
timestamp 1698431365
transform 1 0 54880 0 -1 16128
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698431365
transform 1 0 55776 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 16128
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_11_508
timestamp 1698431365
transform 1 0 58240 0 -1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 16128
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_111
timestamp 1698431365
transform 1 0 13776 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_163
timestamp 1698431365
transform 1 0 19600 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_167
timestamp 1698431365
transform 1 0 20048 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_170
timestamp 1698431365
transform 1 0 20384 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_191
timestamp 1698431365
transform 1 0 22736 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_195
timestamp 1698431365
transform 1 0 23184 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_227
timestamp 1698431365
transform 1 0 26768 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_229
timestamp 1698431365
transform 1 0 26992 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_236
timestamp 1698431365
transform 1 0 27776 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_238
timestamp 1698431365
transform 1 0 28000 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_12_278
timestamp 1698431365
transform 1 0 32480 0 1 16128
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_286
timestamp 1698431365
transform 1 0 33376 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_12_302
timestamp 1698431365
transform 1 0 35168 0 1 16128
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_310
timestamp 1698431365
transform 1 0 36064 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_323
timestamp 1698431365
transform 1 0 37520 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_327
timestamp 1698431365
transform 1 0 37968 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_331
timestamp 1698431365
transform 1 0 38416 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_335
timestamp 1698431365
transform 1 0 38864 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_482
timestamp 1698431365
transform 1 0 55328 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_12_486
timestamp 1698431365
transform 1 0 55776 0 1 16128
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_502
timestamp 1698431365
transform 1 0 57568 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_506
timestamp 1698431365
transform 1 0 58016 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_508
timestamp 1698431365
transform 1 0 58240 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 18144
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 18144
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_13_194
timestamp 1698431365
transform 1 0 23072 0 -1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_202
timestamp 1698431365
transform 1 0 23968 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_216
timestamp 1698431365
transform 1 0 25536 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_13_224
timestamp 1698431365
transform 1 0 26432 0 -1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_230
timestamp 1698431365
transform 1 0 27104 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_13_265
timestamp 1698431365
transform 1 0 31024 0 -1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_13_273
timestamp 1698431365
transform 1 0 31920 0 -1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_277
timestamp 1698431365
transform 1 0 32368 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 18144
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_13_298
timestamp 1698431365
transform 1 0 34720 0 -1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_302
timestamp 1698431365
transform 1 0 35168 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_13_305
timestamp 1698431365
transform 1 0 35504 0 -1 18144
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_321
timestamp 1698431365
transform 1 0 37296 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_323
timestamp 1698431365
transform 1 0 37520 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_326
timestamp 1698431365
transform 1 0 37856 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_354
timestamp 1698431365
transform 1 0 40992 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_369
timestamp 1698431365
transform 1 0 42672 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_373
timestamp 1698431365
transform 1 0 43120 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_375
timestamp 1698431365
transform 1 0 43344 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_378
timestamp 1698431365
transform 1 0 43680 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_382
timestamp 1698431365
transform 1 0 44128 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_408
timestamp 1698431365
transform 1 0 47040 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_426
timestamp 1698431365
transform 1 0 49056 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_428
timestamp 1698431365
transform 1 0 49280 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_460
timestamp 1698431365
transform 1 0 52864 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 18144
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 18144
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 18144
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 18144
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698431365
transform 1 0 15120 0 1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_131
timestamp 1698431365
transform 1 0 16016 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_135
timestamp 1698431365
transform 1 0 16464 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_138
timestamp 1698431365
transform 1 0 16800 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_142
timestamp 1698431365
transform 1 0 17248 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_168
timestamp 1698431365
transform 1 0 20160 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_172
timestamp 1698431365
transform 1 0 20608 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_181
timestamp 1698431365
transform 1 0 21616 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_185
timestamp 1698431365
transform 1 0 22064 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_189
timestamp 1698431365
transform 1 0 22512 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_228
timestamp 1698431365
transform 1 0 26880 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_230
timestamp 1698431365
transform 1 0 27104 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_233
timestamp 1698431365
transform 1 0 27440 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_237
timestamp 1698431365
transform 1 0 27888 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_241
timestamp 1698431365
transform 1 0 28336 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_251
timestamp 1698431365
transform 1 0 29456 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_303
timestamp 1698431365
transform 1 0 35280 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_307
timestamp 1698431365
transform 1 0 35728 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_325
timestamp 1698431365
transform 1 0 37744 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_329
timestamp 1698431365
transform 1 0 38192 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_333
timestamp 1698431365
transform 1 0 38640 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_337
timestamp 1698431365
transform 1 0 39088 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_341
timestamp 1698431365
transform 1 0 39536 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_345
timestamp 1698431365
transform 1 0 39984 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_380
timestamp 1698431365
transform 1 0 43904 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_384
timestamp 1698431365
transform 1 0 44352 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_391
timestamp 1698431365
transform 1 0 45136 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_394
timestamp 1698431365
transform 1 0 45472 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_398
timestamp 1698431365
transform 1 0 45920 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_404
timestamp 1698431365
transform 1 0 46592 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_410
timestamp 1698431365
transform 1 0 47264 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_414
timestamp 1698431365
transform 1 0 47712 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_418
timestamp 1698431365
transform 1 0 48160 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_461
timestamp 1698431365
transform 1 0 52976 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_465
timestamp 1698431365
transform 1 0 53424 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_507
timestamp 1698431365
transform 1 0 58128 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 20160
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 20160
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_168
timestamp 1698431365
transform 1 0 20160 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_199
timestamp 1698431365
transform 1 0 23632 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_205
timestamp 1698431365
transform 1 0 24304 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_222
timestamp 1698431365
transform 1 0 26208 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_226
timestamp 1698431365
transform 1 0 26656 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_230
timestamp 1698431365
transform 1 0 27104 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_236
timestamp 1698431365
transform 1 0 27776 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_240
timestamp 1698431365
transform 1 0 28224 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_244
timestamp 1698431365
transform 1 0 28672 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_274
timestamp 1698431365
transform 1 0 32032 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_278
timestamp 1698431365
transform 1 0 32480 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_300
timestamp 1698431365
transform 1 0 34944 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_304
timestamp 1698431365
transform 1 0 35392 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_306
timestamp 1698431365
transform 1 0 35616 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_15_387
timestamp 1698431365
transform 1 0 44688 0 -1 20160
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_397
timestamp 1698431365
transform 1 0 45808 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_401
timestamp 1698431365
transform 1 0 46256 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_481
timestamp 1698431365
transform 1 0 55216 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_485
timestamp 1698431365
transform 1 0 55664 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_489
timestamp 1698431365
transform 1 0 56112 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 20160
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_508
timestamp 1698431365
transform 1 0 58240 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 20160
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 20160
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 20160
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_16_139
timestamp 1698431365
transform 1 0 16912 0 1 20160
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_147
timestamp 1698431365
transform 1 0 17808 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_167
timestamp 1698431365
transform 1 0 20048 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_190
timestamp 1698431365
transform 1 0 22624 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_194
timestamp 1698431365
transform 1 0 23072 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_198
timestamp 1698431365
transform 1 0 23520 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_202
timestamp 1698431365
transform 1 0 23968 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_206
timestamp 1698431365
transform 1 0 24416 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_210
timestamp 1698431365
transform 1 0 24864 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_214
timestamp 1698431365
transform 1 0 25312 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_217
timestamp 1698431365
transform 1 0 25648 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_221
timestamp 1698431365
transform 1 0 26096 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_225
timestamp 1698431365
transform 1 0 26544 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_229
timestamp 1698431365
transform 1 0 26992 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_233
timestamp 1698431365
transform 1 0 27440 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_237
timestamp 1698431365
transform 1 0 27888 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_241
timestamp 1698431365
transform 1 0 28336 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_253
timestamp 1698431365
transform 1 0 29680 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_285
timestamp 1698431365
transform 1 0 33264 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_289
timestamp 1698431365
transform 1 0 33712 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_293
timestamp 1698431365
transform 1 0 34160 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_297
timestamp 1698431365
transform 1 0 34608 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_299
timestamp 1698431365
transform 1 0 34832 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_321
timestamp 1698431365
transform 1 0 37296 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_350
timestamp 1698431365
transform 1 0 40544 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_391
timestamp 1698431365
transform 1 0 45136 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_393
timestamp 1698431365
transform 1 0 45360 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_396
timestamp 1698431365
transform 1 0 45696 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_400
timestamp 1698431365
transform 1 0 46144 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_404
timestamp 1698431365
transform 1 0 46592 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_408
timestamp 1698431365
transform 1 0 47040 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_437
timestamp 1698431365
transform 1 0 50288 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_476
timestamp 1698431365
transform 1 0 54656 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_480
timestamp 1698431365
transform 1 0 55104 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_484
timestamp 1698431365
transform 1 0 55552 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_488
timestamp 1698431365
transform 1 0 56000 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_16_492
timestamp 1698431365
transform 1 0 56448 0 1 20160
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_508
timestamp 1698431365
transform 1 0 58240 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 22176
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 22176
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 22176
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_158
timestamp 1698431365
transform 1 0 19040 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_162
timestamp 1698431365
transform 1 0 19488 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_17_164
timestamp 1698431365
transform 1 0 19712 0 -1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_203
timestamp 1698431365
transform 1 0 24080 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_17_207
timestamp 1698431365
transform 1 0 24528 0 -1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_226
timestamp 1698431365
transform 1 0 26656 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_230
timestamp 1698431365
transform 1 0 27104 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_234
timestamp 1698431365
transform 1 0 27552 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_278
timestamp 1698431365
transform 1 0 32480 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_17_290
timestamp 1698431365
transform 1 0 33824 0 -1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_297
timestamp 1698431365
transform 1 0 34608 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_301
timestamp 1698431365
transform 1 0 35056 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_313
timestamp 1698431365
transform 1 0 36400 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_317
timestamp 1698431365
transform 1 0 36848 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_321
timestamp 1698431365
transform 1 0 37296 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_325
timestamp 1698431365
transform 1 0 37744 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_331
timestamp 1698431365
transform 1 0 38416 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_335
timestamp 1698431365
transform 1 0 38864 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_339
timestamp 1698431365
transform 1 0 39312 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_343
timestamp 1698431365
transform 1 0 39760 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_347
timestamp 1698431365
transform 1 0 40208 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_356
timestamp 1698431365
transform 1 0 41216 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_360
timestamp 1698431365
transform 1 0 41664 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_364
timestamp 1698431365
transform 1 0 42112 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_374
timestamp 1698431365
transform 1 0 43232 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_378
timestamp 1698431365
transform 1 0 43680 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_384
timestamp 1698431365
transform 1 0 44352 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_413
timestamp 1698431365
transform 1 0 47600 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_417
timestamp 1698431365
transform 1 0 48048 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_17_419
timestamp 1698431365
transform 1 0 48272 0 -1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_426
timestamp 1698431365
transform 1 0 49056 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_459
timestamp 1698431365
transform 1 0 52752 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_486
timestamp 1698431365
transform 1 0 55776 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_17_496
timestamp 1698431365
transform 1 0 56896 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_17_500
timestamp 1698431365
transform 1 0 57344 0 -1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_17_508
timestamp 1698431365
transform 1 0 58240 0 -1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 22176
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 22176
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_143
timestamp 1698431365
transform 1 0 17360 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_18_147
timestamp 1698431365
transform 1 0 17808 0 1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_155
timestamp 1698431365
transform 1 0 18704 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_159
timestamp 1698431365
transform 1 0 19152 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_163
timestamp 1698431365
transform 1 0 19600 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_167
timestamp 1698431365
transform 1 0 20048 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_183
timestamp 1698431365
transform 1 0 21840 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_187
timestamp 1698431365
transform 1 0 22288 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_191
timestamp 1698431365
transform 1 0 22736 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_238
timestamp 1698431365
transform 1 0 28000 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_18_242
timestamp 1698431365
transform 1 0 28448 0 1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_271
timestamp 1698431365
transform 1 0 31696 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_281
timestamp 1698431365
transform 1 0 32816 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_285
timestamp 1698431365
transform 1 0 33264 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_289
timestamp 1698431365
transform 1 0 33712 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_18_293
timestamp 1698431365
transform 1 0 34160 0 1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_301
timestamp 1698431365
transform 1 0 35056 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_305
timestamp 1698431365
transform 1 0 35504 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_309
timestamp 1698431365
transform 1 0 35952 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_313
timestamp 1698431365
transform 1 0 36400 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_355
timestamp 1698431365
transform 1 0 41104 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_359
timestamp 1698431365
transform 1 0 41552 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_363
timestamp 1698431365
transform 1 0 42000 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_367
timestamp 1698431365
transform 1 0 42448 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_18_371
timestamp 1698431365
transform 1 0 42896 0 1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_379
timestamp 1698431365
transform 1 0 43792 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_383
timestamp 1698431365
transform 1 0 44240 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 22176
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_434
timestamp 1698431365
transform 1 0 49952 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_438
timestamp 1698431365
transform 1 0 50400 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_461
timestamp 1698431365
transform 1 0 52976 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_18_465
timestamp 1698431365
transform 1 0 53424 0 1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_505
timestamp 1698431365
transform 1 0 57904 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 24192
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_76
timestamp 1698431365
transform 1 0 9856 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_19_146
timestamp 1698431365
transform 1 0 17696 0 -1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_154
timestamp 1698431365
transform 1 0 18592 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_186
timestamp 1698431365
transform 1 0 22176 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_188
timestamp 1698431365
transform 1 0 22400 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_228
timestamp 1698431365
transform 1 0 26880 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_230
timestamp 1698431365
transform 1 0 27104 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_291
timestamp 1698431365
transform 1 0 33936 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_295
timestamp 1698431365
transform 1 0 34384 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_19_299
timestamp 1698431365
transform 1 0 34832 0 -1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_19_307
timestamp 1698431365
transform 1 0 35728 0 -1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_311
timestamp 1698431365
transform 1 0 36176 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_315
timestamp 1698431365
transform 1 0 36624 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_368
timestamp 1698431365
transform 1 0 42560 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_19_372
timestamp 1698431365
transform 1 0 43008 0 -1 24192
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_390
timestamp 1698431365
transform 1 0 45024 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_394
timestamp 1698431365
transform 1 0 45472 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_417
timestamp 1698431365
transform 1 0 48048 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_419
timestamp 1698431365
transform 1 0 48272 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_432
timestamp 1698431365
transform 1 0 49728 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_436
timestamp 1698431365
transform 1 0 50176 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_440
timestamp 1698431365
transform 1 0 50624 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_442
timestamp 1698431365
transform 1 0 50848 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_469
timestamp 1698431365
transform 1 0 53872 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_471
timestamp 1698431365
transform 1 0 54096 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_496
timestamp 1698431365
transform 1 0 56896 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_19_500
timestamp 1698431365
transform 1 0 57344 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_19_504
timestamp 1698431365
transform 1 0 57792 0 -1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 24192
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 24192
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_157
timestamp 1698431365
transform 1 0 18928 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_161
timestamp 1698431365
transform 1 0 19376 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_167
timestamp 1698431365
transform 1 0 20048 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_183
timestamp 1698431365
transform 1 0 21840 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_231
timestamp 1698431365
transform 1 0 27216 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_235
timestamp 1698431365
transform 1 0 27664 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_239
timestamp 1698431365
transform 1 0 28112 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_276
timestamp 1698431365
transform 1 0 32256 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_20_278
timestamp 1698431365
transform 1 0 32480 0 1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_303
timestamp 1698431365
transform 1 0 35280 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_307
timestamp 1698431365
transform 1 0 35728 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_311
timestamp 1698431365
transform 1 0 36176 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_339
timestamp 1698431365
transform 1 0 39312 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_379
timestamp 1698431365
transform 1 0 43792 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_383
timestamp 1698431365
transform 1 0 44240 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_20_397
timestamp 1698431365
transform 1 0 45808 0 1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_405
timestamp 1698431365
transform 1 0 46704 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_409
timestamp 1698431365
transform 1 0 47152 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_424
timestamp 1698431365
transform 1 0 48832 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_428
timestamp 1698431365
transform 1 0 49280 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_432
timestamp 1698431365
transform 1 0 49728 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_449
timestamp 1698431365
transform 1 0 51632 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_502
timestamp 1698431365
transform 1 0 57568 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_506
timestamp 1698431365
transform 1 0 58016 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_20_508
timestamp 1698431365
transform 1 0 58240 0 1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 26208
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 26208
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_21_88
timestamp 1698431365
transform 1 0 11200 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_96
timestamp 1698431365
transform 1 0 12096 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_155
timestamp 1698431365
transform 1 0 18704 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_21_159
timestamp 1698431365
transform 1 0 19152 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_21_167
timestamp 1698431365
transform 1 0 20048 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_173
timestamp 1698431365
transform 1 0 20720 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_177
timestamp 1698431365
transform 1 0 21168 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_181
timestamp 1698431365
transform 1 0 21616 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_185
timestamp 1698431365
transform 1 0 22064 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_187
timestamp 1698431365
transform 1 0 22288 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_196
timestamp 1698431365
transform 1 0 23296 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_21_234
timestamp 1698431365
transform 1 0 27552 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_240
timestamp 1698431365
transform 1 0 28224 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_244
timestamp 1698431365
transform 1 0 28672 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_248
timestamp 1698431365
transform 1 0 29120 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_316
timestamp 1698431365
transform 1 0 36736 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_320
timestamp 1698431365
transform 1 0 37184 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_348
timestamp 1698431365
transform 1 0 40320 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_21_410
timestamp 1698431365
transform 1 0 47264 0 -1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_418
timestamp 1698431365
transform 1 0 48160 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_426
timestamp 1698431365
transform 1 0 49056 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_430
timestamp 1698431365
transform 1 0 49504 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_434
timestamp 1698431365
transform 1 0 49952 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_438
timestamp 1698431365
transform 1 0 50400 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_442
timestamp 1698431365
transform 1 0 50848 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_446
timestamp 1698431365
transform 1 0 51296 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_450
timestamp 1698431365
transform 1 0 51744 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_452
timestamp 1698431365
transform 1 0 51968 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_455
timestamp 1698431365
transform 1 0 52304 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_459
timestamp 1698431365
transform 1 0 52752 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_496
timestamp 1698431365
transform 1 0 56896 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_21_500
timestamp 1698431365
transform 1 0 57344 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_21_504
timestamp 1698431365
transform 1 0 57792 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_508
timestamp 1698431365
transform 1 0 58240 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 26208
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_22_41
timestamp 1698431365
transform 1 0 5936 0 1 26208
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 26208
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_22_123
timestamp 1698431365
transform 1 0 15120 0 1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_127
timestamp 1698431365
transform 1 0 15568 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_129
timestamp 1698431365
transform 1 0 15792 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_143
timestamp 1698431365
transform 1 0 17360 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_22_190
timestamp 1698431365
transform 1 0 22624 0 1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_194
timestamp 1698431365
transform 1 0 23072 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_226
timestamp 1698431365
transform 1 0 26656 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_230
timestamp 1698431365
transform 1 0 27104 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_22_234
timestamp 1698431365
transform 1 0 27552 0 1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_242
timestamp 1698431365
transform 1 0 28448 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_251
timestamp 1698431365
transform 1 0 29456 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_264
timestamp 1698431365
transform 1 0 30912 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_321
timestamp 1698431365
transform 1 0 37296 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_325
timestamp 1698431365
transform 1 0 37744 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_329
timestamp 1698431365
transform 1 0 38192 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_361
timestamp 1698431365
transform 1 0 41776 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_378
timestamp 1698431365
transform 1 0 43680 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_382
timestamp 1698431365
transform 1 0 44128 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_384
timestamp 1698431365
transform 1 0 44352 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_391
timestamp 1698431365
transform 1 0 45136 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_393
timestamp 1698431365
transform 1 0 45360 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_22_396
timestamp 1698431365
transform 1 0 45696 0 1 26208
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_22_412
timestamp 1698431365
transform 1 0 47488 0 1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_426
timestamp 1698431365
transform 1 0 49056 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_430
timestamp 1698431365
transform 1 0 49504 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_454
timestamp 1698431365
transform 1 0 52192 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_461
timestamp 1698431365
transform 1 0 52976 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_22_503
timestamp 1698431365
transform 1 0 57680 0 1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_507
timestamp 1698431365
transform 1 0 58128 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_23_6
timestamp 1698431365
transform 1 0 2016 0 -1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_14
timestamp 1698431365
transform 1 0 2912 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_23_52
timestamp 1698431365
transform 1 0 7168 0 -1 28224
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_23_105
timestamp 1698431365
transform 1 0 13104 0 -1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_137
timestamp 1698431365
transform 1 0 16688 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_195
timestamp 1698431365
transform 1 0 23184 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_199
timestamp 1698431365
transform 1 0 23632 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_218
timestamp 1698431365
transform 1 0 25760 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_231
timestamp 1698431365
transform 1 0 27216 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_23_235
timestamp 1698431365
transform 1 0 27664 0 -1 28224
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_277
timestamp 1698431365
transform 1 0 32368 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_298
timestamp 1698431365
transform 1 0 34720 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_23_310
timestamp 1698431365
transform 1 0 36064 0 -1 28224
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_326
timestamp 1698431365
transform 1 0 37856 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_330
timestamp 1698431365
transform 1 0 38304 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_334
timestamp 1698431365
transform 1 0 38752 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_338
timestamp 1698431365
transform 1 0 39200 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_342
timestamp 1698431365
transform 1 0 39648 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_346
timestamp 1698431365
transform 1 0 40096 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_356
timestamp 1698431365
transform 1 0 41216 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_360
timestamp 1698431365
transform 1 0 41664 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_389
timestamp 1698431365
transform 1 0 44912 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_393
timestamp 1698431365
transform 1 0 45360 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_397
timestamp 1698431365
transform 1 0 45808 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_401
timestamp 1698431365
transform 1 0 46256 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_409
timestamp 1698431365
transform 1 0 47152 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_413
timestamp 1698431365
transform 1 0 47600 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_416
timestamp 1698431365
transform 1 0 47936 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_483
timestamp 1698431365
transform 1 0 55440 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_487
timestamp 1698431365
transform 1 0 55888 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_489
timestamp 1698431365
transform 1 0 56112 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_501
timestamp 1698431365
transform 1 0 57456 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_23_505
timestamp 1698431365
transform 1 0 57904 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_69
timestamp 1698431365
transform 1 0 9072 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_111
timestamp 1698431365
transform 1 0 13776 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_24_126
timestamp 1698431365
transform 1 0 15456 0 1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_24_158
timestamp 1698431365
transform 1 0 19040 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_166
timestamp 1698431365
transform 1 0 19936 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_168
timestamp 1698431365
transform 1 0 20160 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_189
timestamp 1698431365
transform 1 0 22512 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_24_193
timestamp 1698431365
transform 1 0 22960 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_24_201
timestamp 1698431365
transform 1 0 23856 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_224
timestamp 1698431365
transform 1 0 26432 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_232
timestamp 1698431365
transform 1 0 27328 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_24_236
timestamp 1698431365
transform 1 0 27776 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_249
timestamp 1698431365
transform 1 0 29232 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_271
timestamp 1698431365
transform 1 0 31696 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_273
timestamp 1698431365
transform 1 0 31920 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_300
timestamp 1698431365
transform 1 0 34944 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_304
timestamp 1698431365
transform 1 0 35392 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_308
timestamp 1698431365
transform 1 0 35840 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_312
timestamp 1698431365
transform 1 0 36288 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_24_321
timestamp 1698431365
transform 1 0 37296 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_24_329
timestamp 1698431365
transform 1 0 38192 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_24_339
timestamp 1698431365
transform 1 0 39312 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_343
timestamp 1698431365
transform 1 0 39760 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_24_359
timestamp 1698431365
transform 1 0 41552 0 1 28224
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_377
timestamp 1698431365
transform 1 0 43568 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_381
timestamp 1698431365
transform 1 0 44016 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_393
timestamp 1698431365
transform 1 0 45360 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_395
timestamp 1698431365
transform 1 0 45584 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_438
timestamp 1698431365
transform 1 0 50400 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_24_504
timestamp 1698431365
transform 1 0 57792 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_508
timestamp 1698431365
transform 1 0 58240 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_25_6
timestamp 1698431365
transform 1 0 2016 0 -1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_60
timestamp 1698431365
transform 1 0 8064 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_74
timestamp 1698431365
transform 1 0 9632 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_25_128
timestamp 1698431365
transform 1 0 15680 0 -1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 30240
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_25_174
timestamp 1698431365
transform 1 0 20832 0 -1 30240
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_25_190
timestamp 1698431365
transform 1 0 22624 0 -1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_198
timestamp 1698431365
transform 1 0 23520 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_244
timestamp 1698431365
transform 1 0 28672 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_262
timestamp 1698431365
transform 1 0 30688 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_264
timestamp 1698431365
transform 1 0 30912 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_273
timestamp 1698431365
transform 1 0 31920 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_309
timestamp 1698431365
transform 1 0 35952 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_313
timestamp 1698431365
transform 1 0 36400 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_317
timestamp 1698431365
transform 1 0 36848 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_321
timestamp 1698431365
transform 1 0 37296 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_325
timestamp 1698431365
transform 1 0 37744 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_329
timestamp 1698431365
transform 1 0 38192 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_333
timestamp 1698431365
transform 1 0 38640 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_337
timestamp 1698431365
transform 1 0 39088 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_339
timestamp 1698431365
transform 1 0 39312 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_342
timestamp 1698431365
transform 1 0 39648 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_346
timestamp 1698431365
transform 1 0 40096 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_396
timestamp 1698431365
transform 1 0 45696 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_400
timestamp 1698431365
transform 1 0 46144 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_25_404
timestamp 1698431365
transform 1 0 46592 0 -1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_412
timestamp 1698431365
transform 1 0 47488 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_416
timestamp 1698431365
transform 1 0 47936 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_435
timestamp 1698431365
transform 1 0 50064 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_441
timestamp 1698431365
transform 1 0 50736 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_476
timestamp 1698431365
transform 1 0 54656 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_480
timestamp 1698431365
transform 1 0 55104 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_484
timestamp 1698431365
transform 1 0 55552 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_25_488
timestamp 1698431365
transform 1 0 56000 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 30240
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_508
timestamp 1698431365
transform 1 0 58240 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_26_45
timestamp 1698431365
transform 1 0 6384 0 1 30240
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_26_61
timestamp 1698431365
transform 1 0 8176 0 1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_69
timestamp 1698431365
transform 1 0 9072 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_135
timestamp 1698431365
transform 1 0 16464 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_139
timestamp 1698431365
transform 1 0 16912 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_141
timestamp 1698431365
transform 1 0 17136 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_168
timestamp 1698431365
transform 1 0 20160 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_172
timestamp 1698431365
transform 1 0 20608 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_185
timestamp 1698431365
transform 1 0 22064 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_189
timestamp 1698431365
transform 1 0 22512 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_251
timestamp 1698431365
transform 1 0 29456 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_255
timestamp 1698431365
transform 1 0 29904 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_259
timestamp 1698431365
transform 1 0 30352 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_276
timestamp 1698431365
transform 1 0 32256 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_300
timestamp 1698431365
transform 1 0 34944 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_302
timestamp 1698431365
transform 1 0 35168 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_329
timestamp 1698431365
transform 1 0 38192 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_348
timestamp 1698431365
transform 1 0 40320 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_375
timestamp 1698431365
transform 1 0 43344 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_379
timestamp 1698431365
transform 1 0 43792 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_383
timestamp 1698431365
transform 1 0 44240 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_402
timestamp 1698431365
transform 1 0 46368 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_406
timestamp 1698431365
transform 1 0 46816 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_26_410
timestamp 1698431365
transform 1 0 47264 0 1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_418
timestamp 1698431365
transform 1 0 48160 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_421
timestamp 1698431365
transform 1 0 48496 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_425
timestamp 1698431365
transform 1 0 48944 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_470
timestamp 1698431365
transform 1 0 53984 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_474
timestamp 1698431365
transform 1 0 54432 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_478
timestamp 1698431365
transform 1 0 54880 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_482
timestamp 1698431365
transform 1 0 55328 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_486
timestamp 1698431365
transform 1 0 55776 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_26_490
timestamp 1698431365
transform 1 0 56224 0 1 30240
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_506
timestamp 1698431365
transform 1 0 58016 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_508
timestamp 1698431365
transform 1 0 58240 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_6
timestamp 1698431365
transform 1 0 2016 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_8
timestamp 1698431365
transform 1 0 2240 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_27_43
timestamp 1698431365
transform 1 0 6160 0 -1 32256
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_27_59
timestamp 1698431365
transform 1 0 7952 0 -1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_67
timestamp 1698431365
transform 1 0 8848 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_80
timestamp 1698431365
transform 1 0 10304 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_119
timestamp 1698431365
transform 1 0 14672 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_27_134
timestamp 1698431365
transform 1 0 16352 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_144
timestamp 1698431365
transform 1 0 17472 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_185
timestamp 1698431365
transform 1 0 22064 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_187
timestamp 1698431365
transform 1 0 22288 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_207
timestamp 1698431365
transform 1 0 24528 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_226
timestamp 1698431365
transform 1 0 26656 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_239
timestamp 1698431365
transform 1 0 28112 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_27_243
timestamp 1698431365
transform 1 0 28560 0 -1 32256
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_27_259
timestamp 1698431365
transform 1 0 30352 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_265
timestamp 1698431365
transform 1 0 31024 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_342
timestamp 1698431365
transform 1 0 39648 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_346
timestamp 1698431365
transform 1 0 40096 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_358
timestamp 1698431365
transform 1 0 41440 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_362
timestamp 1698431365
transform 1 0 41888 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_364
timestamp 1698431365
transform 1 0 42112 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_414
timestamp 1698431365
transform 1 0 47712 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_418
timestamp 1698431365
transform 1 0 48160 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_27_438
timestamp 1698431365
transform 1 0 50400 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_442
timestamp 1698431365
transform 1 0 50848 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_446
timestamp 1698431365
transform 1 0 51296 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_450
timestamp 1698431365
transform 1 0 51744 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_454
timestamp 1698431365
transform 1 0 52192 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_484
timestamp 1698431365
transform 1 0 55552 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_488
timestamp 1698431365
transform 1 0 56000 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_27_496
timestamp 1698431365
transform 1 0 56896 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_27_500
timestamp 1698431365
transform 1 0 57344 0 -1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_508
timestamp 1698431365
transform 1 0 58240 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 32256
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_28_18
timestamp 1698431365
transform 1 0 3360 0 1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 32256
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_28_69
timestamp 1698431365
transform 1 0 9072 0 1 32256
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_85
timestamp 1698431365
transform 1 0 10864 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_89
timestamp 1698431365
transform 1 0 11312 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_91
timestamp 1698431365
transform 1 0 11536 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_96
timestamp 1698431365
transform 1 0 12096 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_111
timestamp 1698431365
transform 1 0 13776 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_132
timestamp 1698431365
transform 1 0 16128 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_136
timestamp 1698431365
transform 1 0 16576 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_187
timestamp 1698431365
transform 1 0 22288 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_238
timestamp 1698431365
transform 1 0 28000 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_242
timestamp 1698431365
transform 1 0 28448 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 32256
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_28_263
timestamp 1698431365
transform 1 0 30800 0 1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_271
timestamp 1698431365
transform 1 0 31696 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_296
timestamp 1698431365
transform 1 0 34496 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_300
timestamp 1698431365
transform 1 0 34944 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_304
timestamp 1698431365
transform 1 0 35392 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_308
timestamp 1698431365
transform 1 0 35840 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_312
timestamp 1698431365
transform 1 0 36288 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_323
timestamp 1698431365
transform 1 0 37520 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_335
timestamp 1698431365
transform 1 0 38864 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_339
timestamp 1698431365
transform 1 0 39312 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_372
timestamp 1698431365
transform 1 0 43008 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_376
timestamp 1698431365
transform 1 0 43456 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_380
timestamp 1698431365
transform 1 0 43904 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_393
timestamp 1698431365
transform 1 0 45360 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_28_431
timestamp 1698431365
transform 1 0 49616 0 1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_439
timestamp 1698431365
transform 1 0 50512 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_442
timestamp 1698431365
transform 1 0 50848 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_446
timestamp 1698431365
transform 1 0 51296 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_450
timestamp 1698431365
transform 1 0 51744 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_452
timestamp 1698431365
transform 1 0 51968 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_501
timestamp 1698431365
transform 1 0 57456 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_505
timestamp 1698431365
transform 1 0 57904 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_6
timestamp 1698431365
transform 1 0 2016 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_8
timestamp 1698431365
transform 1 0 2240 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_29_43
timestamp 1698431365
transform 1 0 6160 0 -1 34272
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_29_59
timestamp 1698431365
transform 1 0 7952 0 -1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_67
timestamp 1698431365
transform 1 0 8848 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_76
timestamp 1698431365
transform 1 0 9856 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_78
timestamp 1698431365
transform 1 0 10080 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_99
timestamp 1698431365
transform 1 0 12432 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_124
timestamp 1698431365
transform 1 0 15232 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_146
timestamp 1698431365
transform 1 0 17696 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_29_161
timestamp 1698431365
transform 1 0 19376 0 -1 34272
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_177
timestamp 1698431365
transform 1 0 21168 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_179
timestamp 1698431365
transform 1 0 21392 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_218
timestamp 1698431365
transform 1 0 25760 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_222
timestamp 1698431365
transform 1 0 26208 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_232
timestamp 1698431365
transform 1 0 27328 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_234
timestamp 1698431365
transform 1 0 27552 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_237
timestamp 1698431365
transform 1 0 27888 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_241
timestamp 1698431365
transform 1 0 28336 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_271
timestamp 1698431365
transform 1 0 31696 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_273
timestamp 1698431365
transform 1 0 31920 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_316
timestamp 1698431365
transform 1 0 36736 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_320
timestamp 1698431365
transform 1 0 37184 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_322
timestamp 1698431365
transform 1 0 37408 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_29_325
timestamp 1698431365
transform 1 0 37744 0 -1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_333
timestamp 1698431365
transform 1 0 38640 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_336
timestamp 1698431365
transform 1 0 38976 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_340
timestamp 1698431365
transform 1 0 39424 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_344
timestamp 1698431365
transform 1 0 39872 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_356
timestamp 1698431365
transform 1 0 41216 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_360
timestamp 1698431365
transform 1 0 41664 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_364
timestamp 1698431365
transform 1 0 42112 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_368
timestamp 1698431365
transform 1 0 42560 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_406
timestamp 1698431365
transform 1 0 46816 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_410
timestamp 1698431365
transform 1 0 47264 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_414
timestamp 1698431365
transform 1 0 47712 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_441
timestamp 1698431365
transform 1 0 50736 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_443
timestamp 1698431365
transform 1 0 50960 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_29_505
timestamp 1698431365
transform 1 0 57904 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_30_41
timestamp 1698431365
transform 1 0 5936 0 1 34272
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_57
timestamp 1698431365
transform 1 0 7728 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_61
timestamp 1698431365
transform 1 0 8176 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_63
timestamp 1698431365
transform 1 0 8400 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_30_112
timestamp 1698431365
transform 1 0 13888 0 1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_120
timestamp 1698431365
transform 1 0 14784 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_124
timestamp 1698431365
transform 1 0 15232 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_156
timestamp 1698431365
transform 1 0 18816 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_158
timestamp 1698431365
transform 1 0 19040 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_185
timestamp 1698431365
transform 1 0 22064 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_30_207
timestamp 1698431365
transform 1 0 24528 0 1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_215
timestamp 1698431365
transform 1 0 25424 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_221
timestamp 1698431365
transform 1 0 26096 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_225
timestamp 1698431365
transform 1 0 26544 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_239
timestamp 1698431365
transform 1 0 28112 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_276
timestamp 1698431365
transform 1 0 32256 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_296
timestamp 1698431365
transform 1 0 34496 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_300
timestamp 1698431365
transform 1 0 34944 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_304
timestamp 1698431365
transform 1 0 35392 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_308
timestamp 1698431365
transform 1 0 35840 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_356
timestamp 1698431365
transform 1 0 41216 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_380
timestamp 1698431365
transform 1 0 43904 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_382
timestamp 1698431365
transform 1 0 44128 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_425
timestamp 1698431365
transform 1 0 48944 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_463
timestamp 1698431365
transform 1 0 53200 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_467
timestamp 1698431365
transform 1 0 53648 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_471
timestamp 1698431365
transform 1 0 54096 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_504
timestamp 1698431365
transform 1 0 57792 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_508
timestamp 1698431365
transform 1 0 58240 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_10
timestamp 1698431365
transform 1 0 2464 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_31_46
timestamp 1698431365
transform 1 0 6496 0 -1 36288
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_31_62
timestamp 1698431365
transform 1 0 8288 0 -1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_31_120
timestamp 1698431365
transform 1 0 14784 0 -1 36288
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_146
timestamp 1698431365
transform 1 0 17696 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_169
timestamp 1698431365
transform 1 0 20272 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_173
timestamp 1698431365
transform 1 0 20720 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_179
timestamp 1698431365
transform 1 0 21392 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_187
timestamp 1698431365
transform 1 0 22288 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_277
timestamp 1698431365
transform 1 0 32368 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_279
timestamp 1698431365
transform 1 0 32592 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_290
timestamp 1698431365
transform 1 0 33824 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_294
timestamp 1698431365
transform 1 0 34272 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_31_302
timestamp 1698431365
transform 1 0 35168 0 -1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_310
timestamp 1698431365
transform 1 0 36064 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_314
timestamp 1698431365
transform 1 0 36512 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_318
timestamp 1698431365
transform 1 0 36960 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_320
timestamp 1698431365
transform 1 0 37184 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_323
timestamp 1698431365
transform 1 0 37520 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_346
timestamp 1698431365
transform 1 0 40096 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_382
timestamp 1698431365
transform 1 0 44128 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_386
timestamp 1698431365
transform 1 0 44576 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_390
timestamp 1698431365
transform 1 0 45024 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_394
timestamp 1698431365
transform 1 0 45472 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_31_397
timestamp 1698431365
transform 1 0 45808 0 -1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_31_407
timestamp 1698431365
transform 1 0 46928 0 -1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_415
timestamp 1698431365
transform 1 0 47824 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_417
timestamp 1698431365
transform 1 0 48048 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_453
timestamp 1698431365
transform 1 0 52080 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_457
timestamp 1698431365
transform 1 0 52528 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_489
timestamp 1698431365
transform 1 0 56112 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_496
timestamp 1698431365
transform 1 0 56896 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_500
timestamp 1698431365
transform 1 0 57344 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_504
timestamp 1698431365
transform 1 0 57792 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_508
timestamp 1698431365
transform 1 0 58240 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 36288
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_32_18
timestamp 1698431365
transform 1 0 3360 0 1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_22
timestamp 1698431365
transform 1 0 3808 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_32_69
timestamp 1698431365
transform 1 0 9072 0 1 36288
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_85
timestamp 1698431365
transform 1 0 10864 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_32_88
timestamp 1698431365
transform 1 0 11200 0 1 36288
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_32_111
timestamp 1698431365
transform 1 0 13776 0 1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_32_162
timestamp 1698431365
transform 1 0 19488 0 1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_166
timestamp 1698431365
transform 1 0 19936 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_193
timestamp 1698431365
transform 1 0 22960 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_207
timestamp 1698431365
transform 1 0 24528 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_32_211
timestamp 1698431365
transform 1 0 24976 0 1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_260
timestamp 1698431365
transform 1 0 30464 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_32_264
timestamp 1698431365
transform 1 0 30912 0 1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_272
timestamp 1698431365
transform 1 0 31808 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_274
timestamp 1698431365
transform 1 0 32032 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_32_295
timestamp 1698431365
transform 1 0 34384 0 1 36288
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_32_303
timestamp 1698431365
transform 1 0 35280 0 1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_307
timestamp 1698431365
transform 1 0 35728 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_360
timestamp 1698431365
transform 1 0 41664 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_364
timestamp 1698431365
transform 1 0 42112 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_366
timestamp 1698431365
transform 1 0 42336 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_384
timestamp 1698431365
transform 1 0 44352 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_389
timestamp 1698431365
transform 1 0 44912 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_403
timestamp 1698431365
transform 1 0 46480 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_427
timestamp 1698431365
transform 1 0 49168 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_429
timestamp 1698431365
transform 1 0 49392 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_32_459
timestamp 1698431365
transform 1 0 52752 0 1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_33_10
timestamp 1698431365
transform 1 0 2464 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_14
timestamp 1698431365
transform 1 0 2912 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_33_58
timestamp 1698431365
transform 1 0 7840 0 -1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 8736 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_88
timestamp 1698431365
transform 1 0 11200 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_33_123
timestamp 1698431365
transform 1 0 15120 0 -1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_33_131
timestamp 1698431365
transform 1 0 16016 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_135
timestamp 1698431365
transform 1 0 16464 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_137
timestamp 1698431365
transform 1 0 16688 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_146
timestamp 1698431365
transform 1 0 17696 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_150
timestamp 1698431365
transform 1 0 18144 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_154
timestamp 1698431365
transform 1 0 18592 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_158
timestamp 1698431365
transform 1 0 19040 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_192
timestamp 1698431365
transform 1 0 22848 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_196
timestamp 1698431365
transform 1 0 23296 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_33_200
timestamp 1698431365
transform 1 0 23744 0 -1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_208
timestamp 1698431365
transform 1 0 24640 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_33_234
timestamp 1698431365
transform 1 0 27552 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_238
timestamp 1698431365
transform 1 0 28000 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_241
timestamp 1698431365
transform 1 0 28336 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_33_245
timestamp 1698431365
transform 1 0 28784 0 -1 38304
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_277
timestamp 1698431365
transform 1 0 32368 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_308
timestamp 1698431365
transform 1 0 35840 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_310
timestamp 1698431365
transform 1 0 36064 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_33_317
timestamp 1698431365
transform 1 0 36848 0 -1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_333
timestamp 1698431365
transform 1 0 38640 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_336
timestamp 1698431365
transform 1 0 38976 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_340
timestamp 1698431365
transform 1 0 39424 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_33_344
timestamp 1698431365
transform 1 0 39872 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_33_383
timestamp 1698431365
transform 1 0 44240 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_387
timestamp 1698431365
transform 1 0 44688 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_390
timestamp 1698431365
transform 1 0 45024 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_33_394
timestamp 1698431365
transform 1 0 45472 0 -1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_415
timestamp 1698431365
transform 1 0 47824 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_417
timestamp 1698431365
transform 1 0 48048 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_426
timestamp 1698431365
transform 1 0 49056 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_430
timestamp 1698431365
transform 1 0 49504 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_434
timestamp 1698431365
transform 1 0 49952 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_438
timestamp 1698431365
transform 1 0 50400 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_442
timestamp 1698431365
transform 1 0 50848 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_446
timestamp 1698431365
transform 1 0 51296 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_482
timestamp 1698431365
transform 1 0 55328 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_486
timestamp 1698431365
transform 1 0 55776 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_496
timestamp 1698431365
transform 1 0 56896 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_33_500
timestamp 1698431365
transform 1 0 57344 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_33_504
timestamp 1698431365
transform 1 0 57792 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_33_508
timestamp 1698431365
transform 1 0 58240 0 -1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_34_18
timestamp 1698431365
transform 1 0 3360 0 1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_26
timestamp 1698431365
transform 1 0 4256 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_28
timestamp 1698431365
transform 1 0 4480 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_34_69
timestamp 1698431365
transform 1 0 9072 0 1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_34_85
timestamp 1698431365
transform 1 0 10864 0 1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_34_93
timestamp 1698431365
transform 1 0 11760 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_97
timestamp 1698431365
transform 1 0 12208 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_99
timestamp 1698431365
transform 1 0 12432 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_34_111
timestamp 1698431365
transform 1 0 13776 0 1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_34_127
timestamp 1698431365
transform 1 0 15568 0 1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_137
timestamp 1698431365
transform 1 0 16688 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_141
timestamp 1698431365
transform 1 0 17136 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_145
timestamp 1698431365
transform 1 0 17584 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_183
timestamp 1698431365
transform 1 0 21840 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_185
timestamp 1698431365
transform 1 0 22064 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_188
timestamp 1698431365
transform 1 0 22400 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_34_217
timestamp 1698431365
transform 1 0 25648 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_243
timestamp 1698431365
transform 1 0 28560 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_249
timestamp 1698431365
transform 1 0 29232 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_34_252
timestamp 1698431365
transform 1 0 29568 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_34_258
timestamp 1698431365
transform 1 0 30240 0 1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_34_274
timestamp 1698431365
transform 1 0 32032 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_293
timestamp 1698431365
transform 1 0 34160 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_34_297
timestamp 1698431365
transform 1 0 34608 0 1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_313
timestamp 1698431365
transform 1 0 36400 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_319
timestamp 1698431365
transform 1 0 37072 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_322
timestamp 1698431365
transform 1 0 37408 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_326
timestamp 1698431365
transform 1 0 37856 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_330
timestamp 1698431365
transform 1 0 38304 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_34_374
timestamp 1698431365
transform 1 0 43232 0 1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_382
timestamp 1698431365
transform 1 0 44128 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_384
timestamp 1698431365
transform 1 0 44352 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_34_391
timestamp 1698431365
transform 1 0 45136 0 1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_399
timestamp 1698431365
transform 1 0 46032 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_34_414
timestamp 1698431365
transform 1 0 47712 0 1 38304
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_34_430
timestamp 1698431365
transform 1 0 49504 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_436
timestamp 1698431365
transform 1 0 50176 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_440
timestamp 1698431365
transform 1 0 50624 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_444
timestamp 1698431365
transform 1 0 51072 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_448
timestamp 1698431365
transform 1 0 51520 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_452
timestamp 1698431365
transform 1 0 51968 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_34_454
timestamp 1698431365
transform 1 0 52192 0 1 38304
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_461
timestamp 1698431365
transform 1 0 52976 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_34_465
timestamp 1698431365
transform 1 0 53424 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_34_501
timestamp 1698431365
transform 1 0 57456 0 1 38304
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_35_6
timestamp 1698431365
transform 1 0 2016 0 -1 40320
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_35_56
timestamp 1698431365
transform 1 0 7616 0 -1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_35_64
timestamp 1698431365
transform 1 0 8512 0 -1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_68
timestamp 1698431365
transform 1 0 8960 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_80
timestamp 1698431365
transform 1 0 10304 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_35_115
timestamp 1698431365
transform 1 0 14224 0 -1 40320
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_131
timestamp 1698431365
transform 1 0 16016 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_133
timestamp 1698431365
transform 1 0 16240 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_35_197
timestamp 1698431365
transform 1 0 23408 0 -1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_201
timestamp 1698431365
transform 1 0 23856 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_203
timestamp 1698431365
transform 1 0 24080 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_315
timestamp 1698431365
transform 1 0 36624 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_319
timestamp 1698431365
transform 1 0 37072 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_321
timestamp 1698431365
transform 1 0 37296 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_328
timestamp 1698431365
transform 1 0 38080 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_348
timestamp 1698431365
transform 1 0 40320 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_383
timestamp 1698431365
transform 1 0 44240 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_387
timestamp 1698431365
transform 1 0 44688 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_426
timestamp 1698431365
transform 1 0 49056 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_468
timestamp 1698431365
transform 1 0 53760 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_489
timestamp 1698431365
transform 1 0 56112 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_35_496
timestamp 1698431365
transform 1 0 56896 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_35_500
timestamp 1698431365
transform 1 0 57344 0 -1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_35_508
timestamp 1698431365
transform 1 0 58240 0 -1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_36_45
timestamp 1698431365
transform 1 0 6384 0 1 40320
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_36_61
timestamp 1698431365
transform 1 0 8176 0 1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_69
timestamp 1698431365
transform 1 0 9072 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_36_111
timestamp 1698431365
transform 1 0 13776 0 1 40320
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_36_127
timestamp 1698431365
transform 1 0 15568 0 1 40320
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_135
timestamp 1698431365
transform 1 0 16464 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_139
timestamp 1698431365
transform 1 0 16912 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_143
timestamp 1698431365
transform 1 0 17360 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_181
timestamp 1698431365
transform 1 0 21616 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_185
timestamp 1698431365
transform 1 0 22064 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_189
timestamp 1698431365
transform 1 0 22512 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_193
timestamp 1698431365
transform 1 0 22960 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_196
timestamp 1698431365
transform 1 0 23296 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_242
timestamp 1698431365
transform 1 0 28448 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_249
timestamp 1698431365
transform 1 0 29232 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_252
timestamp 1698431365
transform 1 0 29568 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_256
timestamp 1698431365
transform 1 0 30016 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_312
timestamp 1698431365
transform 1 0 36288 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_314
timestamp 1698431365
transform 1 0 36512 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_373
timestamp 1698431365
transform 1 0 43120 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_36_377
timestamp 1698431365
transform 1 0 43568 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_383
timestamp 1698431365
transform 1 0 44240 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_410
timestamp 1698431365
transform 1 0 47264 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_36_453
timestamp 1698431365
transform 1 0 52080 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_36_492
timestamp 1698431365
transform 1 0 56448 0 1 40320
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_36_508
timestamp 1698431365
transform 1 0 58240 0 1 40320
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_37_6
timestamp 1698431365
transform 1 0 2016 0 -1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_14
timestamp 1698431365
transform 1 0 2912 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_37_53
timestamp 1698431365
transform 1 0 7280 0 -1 42336
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_80
timestamp 1698431365
transform 1 0 10304 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_37_119
timestamp 1698431365
transform 1 0 14672 0 -1 42336
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_37_135
timestamp 1698431365
transform 1 0 16464 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_139
timestamp 1698431365
transform 1 0 16912 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_180
timestamp 1698431365
transform 1 0 21504 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_37_184
timestamp 1698431365
transform 1 0 21952 0 -1 42336
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_37_200
timestamp 1698431365
transform 1 0 23744 0 -1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_208
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_254
timestamp 1698431365
transform 1 0 29792 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_258
timestamp 1698431365
transform 1 0 30240 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_37_262
timestamp 1698431365
transform 1 0 30688 0 -1 42336
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_313
timestamp 1698431365
transform 1 0 36400 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_317
timestamp 1698431365
transform 1 0 36848 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_321
timestamp 1698431365
transform 1 0 37296 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_325
timestamp 1698431365
transform 1 0 37744 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_37_329
timestamp 1698431365
transform 1 0 38192 0 -1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_37_337
timestamp 1698431365
transform 1 0 39088 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_341
timestamp 1698431365
transform 1 0 39536 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_343
timestamp 1698431365
transform 1 0 39760 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_37_360
timestamp 1698431365
transform 1 0 41664 0 -1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_37_368
timestamp 1698431365
transform 1 0 42560 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_374
timestamp 1698431365
transform 1 0 43232 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_378
timestamp 1698431365
transform 1 0 43680 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_426
timestamp 1698431365
transform 1 0 49056 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_440
timestamp 1698431365
transform 1 0 50624 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_37_444
timestamp 1698431365
transform 1 0 51072 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_37_450
timestamp 1698431365
transform 1 0 51744 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_489
timestamp 1698431365
transform 1 0 56112 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_37_508
timestamp 1698431365
transform 1 0 58240 0 -1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_45
timestamp 1698431365
transform 1 0 6384 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_38_49
timestamp 1698431365
transform 1 0 6832 0 1 42336
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_38_65
timestamp 1698431365
transform 1 0 8624 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_69
timestamp 1698431365
transform 1 0 9072 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_38_111
timestamp 1698431365
transform 1 0 13776 0 1 42336
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_38_127
timestamp 1698431365
transform 1 0 15568 0 1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_135
timestamp 1698431365
transform 1 0 16464 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_38_167
timestamp 1698431365
transform 1 0 20048 0 1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_181
timestamp 1698431365
transform 1 0 21616 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_185
timestamp 1698431365
transform 1 0 22064 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_38_227
timestamp 1698431365
transform 1 0 26768 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_231
timestamp 1698431365
transform 1 0 27216 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_234
timestamp 1698431365
transform 1 0 27552 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_38_238
timestamp 1698431365
transform 1 0 28000 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_242
timestamp 1698431365
transform 1 0 28448 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_251
timestamp 1698431365
transform 1 0 29456 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_253
timestamp 1698431365
transform 1 0 29680 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_38_256
timestamp 1698431365
transform 1 0 30016 0 1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_38_264
timestamp 1698431365
transform 1 0 30912 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_268
timestamp 1698431365
transform 1 0 31360 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_301
timestamp 1698431365
transform 1 0 35056 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_305
timestamp 1698431365
transform 1 0 35504 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_307
timestamp 1698431365
transform 1 0 35728 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_38_310
timestamp 1698431365
transform 1 0 36064 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_314
timestamp 1698431365
transform 1 0 36512 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_38_321
timestamp 1698431365
transform 1 0 37296 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_325
timestamp 1698431365
transform 1 0 37744 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_38_328
timestamp 1698431365
transform 1 0 38080 0 1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_38_336
timestamp 1698431365
transform 1 0 38976 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_340
timestamp 1698431365
transform 1 0 39424 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_38_372
timestamp 1698431365
transform 1 0 43008 0 1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_382
timestamp 1698431365
transform 1 0 44128 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_384
timestamp 1698431365
transform 1 0 44352 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_391
timestamp 1698431365
transform 1 0 45136 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_395
timestamp 1698431365
transform 1 0 45584 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_399
timestamp 1698431365
transform 1 0 46032 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_403
timestamp 1698431365
transform 1 0 46480 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_407
timestamp 1698431365
transform 1 0 46928 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_420
timestamp 1698431365
transform 1 0 48384 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_424
timestamp 1698431365
transform 1 0 48832 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_428
timestamp 1698431365
transform 1 0 49280 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_38_432
timestamp 1698431365
transform 1 0 49728 0 1 42336
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_440
timestamp 1698431365
transform 1 0 50624 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_443
timestamp 1698431365
transform 1 0 50960 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_447
timestamp 1698431365
transform 1 0 51408 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_451
timestamp 1698431365
transform 1 0 51856 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_461
timestamp 1698431365
transform 1 0 52976 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_463
timestamp 1698431365
transform 1 0 53200 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_466
timestamp 1698431365
transform 1 0 53536 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_470
timestamp 1698431365
transform 1 0 53984 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_38_474
timestamp 1698431365
transform 1 0 54432 0 1 42336
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_38_506
timestamp 1698431365
transform 1 0 58016 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_38_508
timestamp 1698431365
transform 1 0 58240 0 1 42336
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_82
timestamp 1698431365
transform 1 0 10528 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_39_120
timestamp 1698431365
transform 1 0 14784 0 -1 44352
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_39_170
timestamp 1698431365
transform 1 0 20384 0 -1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_39_202
timestamp 1698431365
transform 1 0 23968 0 -1 44352
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 44352
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_228
timestamp 1698431365
transform 1 0 26880 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_39_230
timestamp 1698431365
transform 1 0 27104 0 -1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_233
timestamp 1698431365
transform 1 0 27440 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_39_272
timestamp 1698431365
transform 1 0 31808 0 -1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_278
timestamp 1698431365
transform 1 0 32480 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_304
timestamp 1698431365
transform 1 0 35392 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_308
timestamp 1698431365
transform 1 0 35840 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_39_342
timestamp 1698431365
transform 1 0 39648 0 -1 44352
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_39_383
timestamp 1698431365
transform 1 0 44240 0 -1 44352
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_391
timestamp 1698431365
transform 1 0 45136 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_39_395
timestamp 1698431365
transform 1 0 45584 0 -1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_405
timestamp 1698431365
transform 1 0 46704 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_409
timestamp 1698431365
transform 1 0 47152 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_39_413
timestamp 1698431365
transform 1 0 47600 0 -1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_39_417
timestamp 1698431365
transform 1 0 48048 0 -1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_39_484
timestamp 1698431365
transform 1 0 55552 0 -1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_39_488
timestamp 1698431365
transform 1 0 56000 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 44352
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_39_508
timestamp 1698431365
transform 1 0 58240 0 -1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 44352
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 44352
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_40_185
timestamp 1698431365
transform 1 0 22064 0 1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_188
timestamp 1698431365
transform 1 0 22400 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_192
timestamp 1698431365
transform 1 0 22848 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_240
timestamp 1698431365
transform 1 0 28224 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_40_242
timestamp 1698431365
transform 1 0 28448 0 1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_40_291
timestamp 1698431365
transform 1 0 33936 0 1 44352
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_40_299
timestamp 1698431365
transform 1 0 34832 0 1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_303
timestamp 1698431365
transform 1 0 35280 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_40_305
timestamp 1698431365
transform 1 0 35504 0 1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_40_308
timestamp 1698431365
transform 1 0 35840 0 1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_40_319
timestamp 1698431365
transform 1 0 37072 0 1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_322
timestamp 1698431365
transform 1 0 37408 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_326
timestamp 1698431365
transform 1 0 37856 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_40_368
timestamp 1698431365
transform 1 0 42560 0 1 44352
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_40_384
timestamp 1698431365
transform 1 0 44352 0 1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_393
timestamp 1698431365
transform 1 0 45360 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_40_412
timestamp 1698431365
transform 1 0 47488 0 1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_40_444
timestamp 1698431365
transform 1 0 51072 0 1 44352
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_40_452
timestamp 1698431365
transform 1 0 51968 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_40_454
timestamp 1698431365
transform 1 0 52192 0 1 44352
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_40_489
timestamp 1698431365
transform 1 0 56112 0 1 44352
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_40_505
timestamp 1698431365
transform 1 0 57904 0 1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_41_6
timestamp 1698431365
transform 1 0 2016 0 -1 46368
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_22
timestamp 1698431365
transform 1 0 3808 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_41_24
timestamp 1698431365
transform 1 0 4032 0 -1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_59
timestamp 1698431365
transform 1 0 7952 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_41_65
timestamp 1698431365
transform 1 0 8624 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_41_69
timestamp 1698431365
transform 1 0 9072 0 -1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_41_76
timestamp 1698431365
transform 1 0 9856 0 -1 46368
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_41_84
timestamp 1698431365
transform 1 0 10752 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_88
timestamp 1698431365
transform 1 0 11200 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_41_94
timestamp 1698431365
transform 1 0 11872 0 -1 46368
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_41_126
timestamp 1698431365
transform 1 0 15456 0 -1 46368
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_41_134
timestamp 1698431365
transform 1 0 16352 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_138
timestamp 1698431365
transform 1 0 16800 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 46368
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 46368
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_41_220
timestamp 1698431365
transform 1 0 25984 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_226
timestamp 1698431365
transform 1 0 26656 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_230
timestamp 1698431365
transform 1 0 27104 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_234
timestamp 1698431365
transform 1 0 27552 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_41_275
timestamp 1698431365
transform 1 0 32144 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_41_286
timestamp 1698431365
transform 1 0 33376 0 -1 46368
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_294
timestamp 1698431365
transform 1 0 34272 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_41_296
timestamp 1698431365
transform 1 0 34496 0 -1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_299
timestamp 1698431365
transform 1 0 34832 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_303
timestamp 1698431365
transform 1 0 35280 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_41_349
timestamp 1698431365
transform 1 0 40432 0 -1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_41_354
timestamp 1698431365
transform 1 0 40992 0 -1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_357
timestamp 1698431365
transform 1 0 41328 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_41_361
timestamp 1698431365
transform 1 0 41776 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 46368
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_41_486
timestamp 1698431365
transform 1 0 55776 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 46368
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_41_508
timestamp 1698431365
transform 1 0 58240 0 -1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 46368
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_41
timestamp 1698431365
transform 1 0 5936 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_42_45
timestamp 1698431365
transform 1 0 6384 0 1 46368
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_42_77
timestamp 1698431365
transform 1 0 9968 0 1 46368
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_42_93
timestamp 1698431365
transform 1 0 11760 0 1 46368
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 46368
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_183
timestamp 1698431365
transform 1 0 21840 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_221
timestamp 1698431365
transform 1 0 26096 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_42_225
timestamp 1698431365
transform 1 0 26544 0 1 46368
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_42_233
timestamp 1698431365
transform 1 0 27440 0 1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_42_236
timestamp 1698431365
transform 1 0 27776 0 1 46368
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_42_244
timestamp 1698431365
transform 1 0 28672 0 1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_251
timestamp 1698431365
transform 1 0 29456 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_255
timestamp 1698431365
transform 1 0 29904 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 36176 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 46368
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_333
timestamp 1698431365
transform 1 0 38640 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_42_335
timestamp 1698431365
transform 1 0 38864 0 1 46368
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_338
timestamp 1698431365
transform 1 0 39200 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_42_342
timestamp 1698431365
transform 1 0 39648 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 46368
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_42_451
timestamp 1698431365
transform 1 0 51856 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_42_457
timestamp 1698431365
transform 1 0 52528 0 1 46368
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_42_489
timestamp 1698431365
transform 1 0 56112 0 1 46368
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_42_505
timestamp 1698431365
transform 1 0 57904 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 48384
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_10
timestamp 1698431365
transform 1 0 2464 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_43_14
timestamp 1698431365
transform 1 0 2912 0 -1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_43_49
timestamp 1698431365
transform 1 0 6832 0 -1 48384
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_65
timestamp 1698431365
transform 1 0 8624 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_43_69
timestamp 1698431365
transform 1 0 9072 0 -1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 48384
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 48384
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_43_248
timestamp 1698431365
transform 1 0 29120 0 -1 48384
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 48384
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_298
timestamp 1698431365
transform 1 0 34720 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_302
timestamp 1698431365
transform 1 0 35168 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_306
timestamp 1698431365
transform 1 0 35616 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_310
timestamp 1698431365
transform 1 0 36064 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_43_354
timestamp 1698431365
transform 1 0 40992 0 -1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_43_383
timestamp 1698431365
transform 1 0 44240 0 -1 48384
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_415
timestamp 1698431365
transform 1 0 47824 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_43_419
timestamp 1698431365
transform 1 0 48272 0 -1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 48384
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_43_486
timestamp 1698431365
transform 1 0 55776 0 -1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 48384
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_43_508
timestamp 1698431365
transform 1 0 58240 0 -1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 48384
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 48384
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 48384
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 48384
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 48384
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_265
timestamp 1698431365
transform 1 0 31024 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_269
timestamp 1698431365
transform 1 0 31472 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_44_308
timestamp 1698431365
transform 1 0 35840 0 1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_44_312
timestamp 1698431365
transform 1 0 36288 0 1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_44_319
timestamp 1698431365
transform 1 0 37072 0 1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_350
timestamp 1698431365
transform 1 0 40544 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_354
timestamp 1698431365
transform 1 0 40992 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_44_358
timestamp 1698431365
transform 1 0 41440 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_44_362
timestamp 1698431365
transform 1 0 41888 0 1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_44_384
timestamp 1698431365
transform 1 0 44352 0 1 48384
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 48384
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_44_451
timestamp 1698431365
transform 1 0 51856 0 1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 48384
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_44_489
timestamp 1698431365
transform 1 0 56112 0 1 48384
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_44_505
timestamp 1698431365
transform 1 0 57904 0 1 48384
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 50400
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_314
timestamp 1698431365
transform 1 0 36512 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_45_320
timestamp 1698431365
transform 1 0 37184 0 -1 50400
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_45_336
timestamp 1698431365
transform 1 0 38976 0 -1 50400
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_344
timestamp 1698431365
transform 1 0 39872 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_45_348
timestamp 1698431365
transform 1 0 40320 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_45_356
timestamp 1698431365
transform 1 0 41216 0 -1 50400
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_45_359
timestamp 1698431365
transform 1 0 41552 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_45_363
timestamp 1698431365
transform 1 0 42000 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_45_367
timestamp 1698431365
transform 1 0 42448 0 -1 50400
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_45_399
timestamp 1698431365
transform 1 0 46032 0 -1 50400
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_415
timestamp 1698431365
transform 1 0 47824 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_45_419
timestamp 1698431365
transform 1 0 48272 0 -1 50400
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_45_422
timestamp 1698431365
transform 1 0 48608 0 -1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_45_486
timestamp 1698431365
transform 1 0 55776 0 -1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 50400
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_45_508
timestamp 1698431365
transform 1 0 58240 0 -1 50400
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 50400
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 50400
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_381
timestamp 1698431365
transform 1 0 44016 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 50400
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_451
timestamp 1698431365
transform 1 0 51856 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 50400
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_46_489
timestamp 1698431365
transform 1 0 56112 0 1 50400
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_46_505
timestamp 1698431365
transform 1 0 57904 0 1 50400
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 52416
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_34
timestamp 1698431365
transform 1 0 5152 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_47_38
timestamp 1698431365
transform 1 0 5600 0 -1 52416
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_47_43
timestamp 1698431365
transform 1 0 6160 0 -1 52416
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_47_59
timestamp 1698431365
transform 1 0 7952 0 -1 52416
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_47_67
timestamp 1698431365
transform 1 0 8848 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_47_69
timestamp 1698431365
transform 1 0 9072 0 -1 52416
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698431365
transform 1 0 32256 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_346
timestamp 1698431365
transform 1 0 40096 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698431365
transform 1 0 47936 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_47_422
timestamp 1698431365
transform 1 0 48608 0 -1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_47_486
timestamp 1698431365
transform 1 0 55776 0 -1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 52416
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_47_508
timestamp 1698431365
transform 1 0 58240 0 -1 52416
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 52416
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 52416
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698431365
transform 1 0 44016 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 52416
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_451
timestamp 1698431365
transform 1 0 51856 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_48_457
timestamp 1698431365
transform 1 0 52528 0 1 52416
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_48_489
timestamp 1698431365
transform 1 0 56112 0 1 52416
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_48_505
timestamp 1698431365
transform 1 0 57904 0 1 52416
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698431365
transform 1 0 8736 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_49_136
timestamp 1698431365
transform 1 0 16576 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_49_346
timestamp 1698431365
transform 1 0 40096 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_49_416
timestamp 1698431365
transform 1 0 47936 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 54432
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_49_454
timestamp 1698431365
transform 1 0 52192 0 -1 54432
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_49_470
timestamp 1698431365
transform 1 0 53984 0 -1 54432
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_49_478
timestamp 1698431365
transform 1 0 54880 0 -1 54432
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_49_483
timestamp 1698431365
transform 1 0 55440 0 -1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_49_487
timestamp 1698431365
transform 1 0 55888 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_49_489
timestamp 1698431365
transform 1 0 56112 0 -1 54432
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 54432
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_49_508
timestamp 1698431365
transform 1 0 58240 0 -1 54432
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 54432
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 54432
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_101
timestamp 1698431365
transform 1 0 12656 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_171
timestamp 1698431365
transform 1 0 20496 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_241
timestamp 1698431365
transform 1 0 28336 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_311
timestamp 1698431365
transform 1 0 36176 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698431365
transform 1 0 44016 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 54432
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_451
timestamp 1698431365
transform 1 0 51856 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_50_457
timestamp 1698431365
transform 1 0 52528 0 1 54432
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_50_489
timestamp 1698431365
transform 1 0 56112 0 1 54432
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_50_505
timestamp 1698431365
transform 1 0 57904 0 1 54432
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_36
timestamp 1698431365
transform 1 0 5376 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_70
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_104
timestamp 1698431365
transform 1 0 12992 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_138
timestamp 1698431365
transform 1 0 16800 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_172
timestamp 1698431365
transform 1 0 20608 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_206
timestamp 1698431365
transform 1 0 24416 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_240
timestamp 1698431365
transform 1 0 28224 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_274
timestamp 1698431365
transform 1 0 32032 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_308
timestamp 1698431365
transform 1 0 35840 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_342
timestamp 1698431365
transform 1 0 39648 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_376
timestamp 1698431365
transform 1 0 43456 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_410
timestamp 1698431365
transform 1 0 47264 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_51_444
timestamp 1698431365
transform 1 0 51072 0 -1 56448
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_51_478
timestamp 1698431365
transform 1 0 54880 0 -1 56448
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_51_494
timestamp 1698431365
transform 1 0 56672 0 -1 56448
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_51_502
timestamp 1698431365
transform 1 0 57568 0 -1 56448
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_51_506
timestamp 1698431365
transform 1 0 58016 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_51_508
timestamp 1698431365
transform 1 0 58240 0 -1 56448
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_0_Left_52 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 4032
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 4032
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_1_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 6048
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 6048
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_2_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 6048
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 6048
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_3_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 8064
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 8064
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_4_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 8064
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 8064
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_5_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 10080
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 10080
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_6_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 10080
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 10080
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_7_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 12096
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 12096
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_8_Left_60
timestamp 1698431365
transform 1 0 1344 0 1 12096
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 12096
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_9_Left_61
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_10_Left_62
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_11_Left_63
timestamp 1698431365
transform 1 0 1344 0 -1 16128
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 16128
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_12_Left_64
timestamp 1698431365
transform 1 0 1344 0 1 16128
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 16128
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_13_Left_65
timestamp 1698431365
transform 1 0 1344 0 -1 18144
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 18144
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_14_Left_66
timestamp 1698431365
transform 1 0 1344 0 1 18144
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 18144
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_15_Left_67
timestamp 1698431365
transform 1 0 1344 0 -1 20160
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 20160
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_16_Left_68
timestamp 1698431365
transform 1 0 1344 0 1 20160
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 20160
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_17_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 22176
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 22176
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_18_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 22176
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 22176
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_19_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 24192
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 24192
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_20_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 24192
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 24192
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_21_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 26208
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 26208
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_22_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 26208
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 26208
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_23_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_24_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_25_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 30240
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 30240
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_26_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 30240
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 30240
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_27_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 32256
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 32256
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_28_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 32256
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 32256
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_29_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 34272
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 34272
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_30_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 34272
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 34272
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_31_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 36288
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 36288
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_32_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 36288
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 36288
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_33_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 38304
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 38304
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_34_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 38304
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 38304
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_35_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 40320
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 40320
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_36_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 40320
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 40320
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_37_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 42336
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_38_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 42336
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_39_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 44352
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 44352
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_40_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 44352
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 44352
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_41_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 46368
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 46368
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_42_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 46368
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 46368
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_43_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 48384
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 58576 0 -1 48384
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_44_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 48384
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 58576 0 1 48384
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_45_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 50400
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 58576 0 -1 50400
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_46_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 50400
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 58576 0 1 50400
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_47_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 52416
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 58576 0 -1 52416
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_48_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 52416
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 58576 0 1 52416
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_49_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 54432
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 58576 0 -1 54432
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_50_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 54432
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 58576 0 1 54432
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_51_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 58576 0 -1 56448
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__icgtp_1  ro_inst.clock_gate
timestamp 1698431365
transform 1 0 10080 0 1 34272
box -86 -90 3110 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.clock_gate_inv
timestamp 1698431365
transform -1 0 12096 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[1\].div_flop
timestamp 1698431365
transform 1 0 10640 0 -1 32256
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[1\].div_flop_inv
timestamp 1698431365
transform -1 0 14672 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[2\].div_flop
timestamp 1698431365
transform 1 0 10640 0 -1 30240
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[2\].div_flop_inv
timestamp 1698431365
transform -1 0 13776 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[3\].div_flop_inv
timestamp 1698431365
transform -1 0 10640 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[3\].div_flop
timestamp 1698431365
transform 1 0 9520 0 1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[4\].div_flop
timestamp 1698431365
transform 1 0 9520 0 1 30240
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[4\].div_flop_inv
timestamp 1698431365
transform -1 0 10192 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[5\].div_flop_inv
timestamp 1698431365
transform -1 0 9184 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[5\].div_flop
timestamp 1698431365
transform 1 0 9520 0 -1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[6\].div_flop_inv
timestamp 1698431365
transform 1 0 5936 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[6\].div_flop
timestamp 1698431365
transform -1 0 8064 0 -1 30240
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[7\].div_flop_inv
timestamp 1698431365
transform 1 0 4032 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[7\].div_flop
timestamp 1698431365
transform -1 0 7168 0 -1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[8\].div_flop_inv
timestamp 1698431365
transform -1 0 3584 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[8\].div_flop
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[9\].div_flop_inv
timestamp 1698431365
transform 1 0 3584 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[9\].div_flop
timestamp 1698431365
transform -1 0 5264 0 1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[10\].div_flop
timestamp 1698431365
transform 1 0 1680 0 1 30240
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[10\].div_flop_inv
timestamp 1698431365
transform -1 0 5936 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[11\].div_flop_inv
timestamp 1698431365
transform -1 0 5152 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[11\].div_flop
timestamp 1698431365
transform 1 0 2576 0 -1 32256
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[12\].div_flop
timestamp 1698431365
transform 1 0 2576 0 -1 34272
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[12\].div_flop_inv
timestamp 1698431365
transform -1 0 4704 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[13\].div_flop_inv
timestamp 1698431365
transform -1 0 5936 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[13\].div_flop
timestamp 1698431365
transform 1 0 1680 0 1 34272
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[14\].div_flop_inv
timestamp 1698431365
transform -1 0 5152 0 1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[14\].div_flop
timestamp 1698431365
transform 1 0 2912 0 -1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[15\].div_flop
timestamp 1698431365
transform 1 0 3360 0 -1 38304
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[15\].div_flop_inv
timestamp 1698431365
transform -1 0 4704 0 1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[16\].div_flop
timestamp 1698431365
transform 1 0 4032 0 -1 40320
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[16\].div_flop_inv
timestamp 1698431365
transform -1 0 7392 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[17\].div_flop
timestamp 1698431365
transform 1 0 5488 0 1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[17\].div_flop_inv
timestamp 1698431365
transform -1 0 7840 0 -1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[18\].div_flop_inv
timestamp 1698431365
transform -1 0 5264 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[18\].div_flop
timestamp 1698431365
transform -1 0 9072 0 1 38304
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[19\].div_flop
timestamp 1698431365
transform 1 0 3696 0 -1 42336
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[19\].div_flop_inv
timestamp 1698431365
transform -1 0 5936 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[20\].div_flop_inv
timestamp 1698431365
transform -1 0 6384 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[20\].div_flop
timestamp 1698431365
transform 1 0 1680 0 1 40320
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[21\].div_flop
timestamp 1698431365
transform 1 0 1680 0 1 42336
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[21\].div_flop_inv
timestamp 1698431365
transform -1 0 3696 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[22\].div_flop
timestamp 1698431365
transform 1 0 2016 0 -1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[22\].div_flop_inv
timestamp 1698431365
transform -1 0 5936 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[23\].div_flop
timestamp 1698431365
transform 1 0 1680 0 1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[23\].div_flop_inv
timestamp 1698431365
transform -1 0 6384 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[24\].div_flop
timestamp 1698431365
transform 1 0 3248 0 -1 48384
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[24\].div_flop_inv
timestamp 1698431365
transform -1 0 5936 0 1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[25\].div_flop
timestamp 1698431365
transform 1 0 4368 0 -1 46368
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[25\].div_flop_inv
timestamp 1698431365
transform -1 0 5936 0 1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[26\].div_flop_inv
timestamp 1698431365
transform -1 0 8624 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[26\].div_flop
timestamp 1698431365
transform 1 0 5600 0 -1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[27\].div_flop_inv
timestamp 1698431365
transform -1 0 10528 0 -1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[27\].div_flop
timestamp 1698431365
transform 1 0 5936 0 1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[28\].div_flop_inv
timestamp 1698431365
transform -1 0 11872 0 -1 46368
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[28\].div_flop
timestamp 1698431365
transform 1 0 9520 0 1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[29\].div_flop_inv
timestamp 1698431365
transform -1 0 14784 0 -1 44352
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[29\].div_flop
timestamp 1698431365
transform 1 0 9520 0 1 42336
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[30\].div_flop
timestamp 1698431365
transform 1 0 10752 0 -1 44352
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[30\].div_flop_inv
timestamp 1698431365
transform -1 0 13776 0 1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[31\].div_flop_inv
timestamp 1698431365
transform -1 0 14672 0 -1 42336
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[31\].div_flop
timestamp 1698431365
transform 1 0 10640 0 -1 42336
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[32\].div_flop_inv
timestamp 1698431365
transform -1 0 13776 0 1 40320
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[32\].div_flop
timestamp 1698431365
transform 1 0 9520 0 1 40320
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[33\].div_flop
timestamp 1698431365
transform 1 0 10640 0 -1 40320
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[33\].div_flop_inv
timestamp 1698431365
transform -1 0 12992 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.gcount\[34\].div_flop_inv
timestamp 1698431365
transform -1 0 13776 0 1 38304
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__dffrnq_1  ro_inst.gcount\[34\].div_flop
timestamp 1698431365
transform 1 0 11536 0 -1 38304
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  ro_inst.ring_osc_0
timestamp 1698431365
transform -1 0 13888 0 1 34272
box -86 -90 646 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.ring_osc_1
timestamp 1698431365
transform -1 0 13776 0 1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.ring_osc_2
timestamp 1698431365
transform 1 0 9632 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor2_1  ro_inst.sig_cmp
timestamp 1698431365
transform -1 0 11200 0 -1 36288
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__latq_1  ro_inst.sig_latch
timestamp 1698431365
transform 1 0 10192 0 -1 34272
box -86 -90 2326 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  ro_inst.slow_clock_inv
timestamp 1698431365
transform 1 0 9184 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_104 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_105
timestamp 1698431365
transform 1 0 8960 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_106
timestamp 1698431365
transform 1 0 12768 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 16576 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_108
timestamp 1698431365
transform 1 0 20384 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_109
timestamp 1698431365
transform 1 0 24192 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_110
timestamp 1698431365
transform 1 0 28000 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 31808 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 35616 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 39424 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 43232 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 47040 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 50848 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_117
timestamp 1698431365
transform 1 0 54656 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_118
timestamp 1698431365
transform 1 0 9184 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_119
timestamp 1698431365
transform 1 0 17024 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_120
timestamp 1698431365
transform 1 0 24864 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_121
timestamp 1698431365
transform 1 0 32704 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_122
timestamp 1698431365
transform 1 0 40544 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_123
timestamp 1698431365
transform 1 0 48384 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_124
timestamp 1698431365
transform 1 0 56224 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_125
timestamp 1698431365
transform 1 0 5264 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_126
timestamp 1698431365
transform 1 0 13104 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_127
timestamp 1698431365
transform 1 0 20944 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_128
timestamp 1698431365
transform 1 0 28784 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_129
timestamp 1698431365
transform 1 0 36624 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_130
timestamp 1698431365
transform 1 0 44464 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_131
timestamp 1698431365
transform 1 0 52304 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_132
timestamp 1698431365
transform 1 0 9184 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_133
timestamp 1698431365
transform 1 0 17024 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_134
timestamp 1698431365
transform 1 0 24864 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_135
timestamp 1698431365
transform 1 0 32704 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_136
timestamp 1698431365
transform 1 0 40544 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_137
timestamp 1698431365
transform 1 0 48384 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_138
timestamp 1698431365
transform 1 0 56224 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_139
timestamp 1698431365
transform 1 0 5264 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_140
timestamp 1698431365
transform 1 0 13104 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_141
timestamp 1698431365
transform 1 0 20944 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_142
timestamp 1698431365
transform 1 0 28784 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_143
timestamp 1698431365
transform 1 0 36624 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_144
timestamp 1698431365
transform 1 0 44464 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_145
timestamp 1698431365
transform 1 0 52304 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_146
timestamp 1698431365
transform 1 0 9184 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_147
timestamp 1698431365
transform 1 0 17024 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_148
timestamp 1698431365
transform 1 0 24864 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_149
timestamp 1698431365
transform 1 0 32704 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_150
timestamp 1698431365
transform 1 0 40544 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_151
timestamp 1698431365
transform 1 0 48384 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_152
timestamp 1698431365
transform 1 0 56224 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_153
timestamp 1698431365
transform 1 0 5264 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_154
timestamp 1698431365
transform 1 0 13104 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_155
timestamp 1698431365
transform 1 0 20944 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_156
timestamp 1698431365
transform 1 0 28784 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_157
timestamp 1698431365
transform 1 0 36624 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_158
timestamp 1698431365
transform 1 0 44464 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_159
timestamp 1698431365
transform 1 0 52304 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_160
timestamp 1698431365
transform 1 0 9184 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_161
timestamp 1698431365
transform 1 0 17024 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_162
timestamp 1698431365
transform 1 0 24864 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_163
timestamp 1698431365
transform 1 0 32704 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_164
timestamp 1698431365
transform 1 0 40544 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_165
timestamp 1698431365
transform 1 0 48384 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_166
timestamp 1698431365
transform 1 0 56224 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_167
timestamp 1698431365
transform 1 0 5264 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_168
timestamp 1698431365
transform 1 0 13104 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_169
timestamp 1698431365
transform 1 0 20944 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_170
timestamp 1698431365
transform 1 0 28784 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_171
timestamp 1698431365
transform 1 0 36624 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_172
timestamp 1698431365
transform 1 0 44464 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_173
timestamp 1698431365
transform 1 0 52304 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_174
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_175
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_176
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_177
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_178
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_179
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_180
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_181
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_182
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_183
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_184
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_185
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_186
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_187
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_188
timestamp 1698431365
transform 1 0 9184 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_189
timestamp 1698431365
transform 1 0 17024 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_190
timestamp 1698431365
transform 1 0 24864 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_191
timestamp 1698431365
transform 1 0 32704 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_192
timestamp 1698431365
transform 1 0 40544 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_193
timestamp 1698431365
transform 1 0 48384 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_194
timestamp 1698431365
transform 1 0 56224 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_195
timestamp 1698431365
transform 1 0 5264 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_196
timestamp 1698431365
transform 1 0 13104 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_197
timestamp 1698431365
transform 1 0 20944 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_198
timestamp 1698431365
transform 1 0 28784 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_199
timestamp 1698431365
transform 1 0 36624 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_200
timestamp 1698431365
transform 1 0 44464 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_201
timestamp 1698431365
transform 1 0 52304 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_202
timestamp 1698431365
transform 1 0 9184 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_203
timestamp 1698431365
transform 1 0 17024 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_204
timestamp 1698431365
transform 1 0 24864 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_205
timestamp 1698431365
transform 1 0 32704 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_206
timestamp 1698431365
transform 1 0 40544 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_207
timestamp 1698431365
transform 1 0 48384 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_208
timestamp 1698431365
transform 1 0 56224 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_209
timestamp 1698431365
transform 1 0 5264 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_210
timestamp 1698431365
transform 1 0 13104 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_211
timestamp 1698431365
transform 1 0 20944 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_212
timestamp 1698431365
transform 1 0 28784 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_213
timestamp 1698431365
transform 1 0 36624 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_214
timestamp 1698431365
transform 1 0 44464 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_215
timestamp 1698431365
transform 1 0 52304 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_216
timestamp 1698431365
transform 1 0 9184 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_217
timestamp 1698431365
transform 1 0 17024 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_218
timestamp 1698431365
transform 1 0 24864 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_219
timestamp 1698431365
transform 1 0 32704 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_220
timestamp 1698431365
transform 1 0 40544 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_221
timestamp 1698431365
transform 1 0 48384 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_222
timestamp 1698431365
transform 1 0 56224 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_223
timestamp 1698431365
transform 1 0 5264 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_224
timestamp 1698431365
transform 1 0 13104 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_225
timestamp 1698431365
transform 1 0 20944 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_226
timestamp 1698431365
transform 1 0 28784 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_227
timestamp 1698431365
transform 1 0 36624 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_228
timestamp 1698431365
transform 1 0 44464 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_229
timestamp 1698431365
transform 1 0 52304 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_230
timestamp 1698431365
transform 1 0 9184 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_231
timestamp 1698431365
transform 1 0 17024 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_232
timestamp 1698431365
transform 1 0 24864 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_233
timestamp 1698431365
transform 1 0 32704 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_234
timestamp 1698431365
transform 1 0 40544 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_235
timestamp 1698431365
transform 1 0 48384 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_236
timestamp 1698431365
transform 1 0 56224 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_237
timestamp 1698431365
transform 1 0 5264 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_238
timestamp 1698431365
transform 1 0 13104 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_239
timestamp 1698431365
transform 1 0 20944 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_240
timestamp 1698431365
transform 1 0 28784 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_241
timestamp 1698431365
transform 1 0 36624 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_242
timestamp 1698431365
transform 1 0 44464 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_243
timestamp 1698431365
transform 1 0 52304 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_244
timestamp 1698431365
transform 1 0 9184 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_245
timestamp 1698431365
transform 1 0 17024 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_246
timestamp 1698431365
transform 1 0 24864 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_247
timestamp 1698431365
transform 1 0 32704 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_248
timestamp 1698431365
transform 1 0 40544 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_249
timestamp 1698431365
transform 1 0 48384 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_250
timestamp 1698431365
transform 1 0 56224 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_251
timestamp 1698431365
transform 1 0 5264 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_252
timestamp 1698431365
transform 1 0 13104 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_253
timestamp 1698431365
transform 1 0 20944 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_254
timestamp 1698431365
transform 1 0 28784 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_255
timestamp 1698431365
transform 1 0 36624 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_256
timestamp 1698431365
transform 1 0 44464 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_257
timestamp 1698431365
transform 1 0 52304 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_258
timestamp 1698431365
transform 1 0 9184 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_259
timestamp 1698431365
transform 1 0 17024 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_260
timestamp 1698431365
transform 1 0 24864 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_261
timestamp 1698431365
transform 1 0 32704 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_262
timestamp 1698431365
transform 1 0 40544 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_263
timestamp 1698431365
transform 1 0 48384 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_264
timestamp 1698431365
transform 1 0 56224 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_265
timestamp 1698431365
transform 1 0 5264 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_266
timestamp 1698431365
transform 1 0 13104 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_267
timestamp 1698431365
transform 1 0 20944 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_268
timestamp 1698431365
transform 1 0 28784 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_269
timestamp 1698431365
transform 1 0 36624 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_270
timestamp 1698431365
transform 1 0 44464 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_271
timestamp 1698431365
transform 1 0 52304 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_272
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_273
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_274
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_275
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_276
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_277
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_278
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_279
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_280
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_281
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_282
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_283
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_284
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_285
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_286
timestamp 1698431365
transform 1 0 9184 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_287
timestamp 1698431365
transform 1 0 17024 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_288
timestamp 1698431365
transform 1 0 24864 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_289
timestamp 1698431365
transform 1 0 32704 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_290
timestamp 1698431365
transform 1 0 40544 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_291
timestamp 1698431365
transform 1 0 48384 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_292
timestamp 1698431365
transform 1 0 56224 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_293
timestamp 1698431365
transform 1 0 5264 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_294
timestamp 1698431365
transform 1 0 13104 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_295
timestamp 1698431365
transform 1 0 20944 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_296
timestamp 1698431365
transform 1 0 28784 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_297
timestamp 1698431365
transform 1 0 36624 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_298
timestamp 1698431365
transform 1 0 44464 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_299
timestamp 1698431365
transform 1 0 52304 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_300
timestamp 1698431365
transform 1 0 9184 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_301
timestamp 1698431365
transform 1 0 17024 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_302
timestamp 1698431365
transform 1 0 24864 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_303
timestamp 1698431365
transform 1 0 32704 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_304
timestamp 1698431365
transform 1 0 40544 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_305
timestamp 1698431365
transform 1 0 48384 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_306
timestamp 1698431365
transform 1 0 56224 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_307
timestamp 1698431365
transform 1 0 5264 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_308
timestamp 1698431365
transform 1 0 13104 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_309
timestamp 1698431365
transform 1 0 20944 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_310
timestamp 1698431365
transform 1 0 28784 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_311
timestamp 1698431365
transform 1 0 36624 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_312
timestamp 1698431365
transform 1 0 44464 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_313
timestamp 1698431365
transform 1 0 52304 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_314
timestamp 1698431365
transform 1 0 9184 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_315
timestamp 1698431365
transform 1 0 17024 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_316
timestamp 1698431365
transform 1 0 24864 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_317
timestamp 1698431365
transform 1 0 32704 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_318
timestamp 1698431365
transform 1 0 40544 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_319
timestamp 1698431365
transform 1 0 48384 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_320
timestamp 1698431365
transform 1 0 56224 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_321
timestamp 1698431365
transform 1 0 5264 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_322
timestamp 1698431365
transform 1 0 13104 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_323
timestamp 1698431365
transform 1 0 20944 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_324
timestamp 1698431365
transform 1 0 28784 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_325
timestamp 1698431365
transform 1 0 36624 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_326
timestamp 1698431365
transform 1 0 44464 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_327
timestamp 1698431365
transform 1 0 52304 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_328
timestamp 1698431365
transform 1 0 9184 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_329
timestamp 1698431365
transform 1 0 17024 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_330
timestamp 1698431365
transform 1 0 24864 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_331
timestamp 1698431365
transform 1 0 32704 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_332
timestamp 1698431365
transform 1 0 40544 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_333
timestamp 1698431365
transform 1 0 48384 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_334
timestamp 1698431365
transform 1 0 56224 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_335
timestamp 1698431365
transform 1 0 5264 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_336
timestamp 1698431365
transform 1 0 13104 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_337
timestamp 1698431365
transform 1 0 20944 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_338
timestamp 1698431365
transform 1 0 28784 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_339
timestamp 1698431365
transform 1 0 36624 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_340
timestamp 1698431365
transform 1 0 44464 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_32_341
timestamp 1698431365
transform 1 0 52304 0 1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_342
timestamp 1698431365
transform 1 0 9184 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_343
timestamp 1698431365
transform 1 0 17024 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_344
timestamp 1698431365
transform 1 0 24864 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_345
timestamp 1698431365
transform 1 0 32704 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_346
timestamp 1698431365
transform 1 0 40544 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_347
timestamp 1698431365
transform 1 0 48384 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_33_348
timestamp 1698431365
transform 1 0 56224 0 -1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_349
timestamp 1698431365
transform 1 0 5264 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_350
timestamp 1698431365
transform 1 0 13104 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_351
timestamp 1698431365
transform 1 0 20944 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_352
timestamp 1698431365
transform 1 0 28784 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_353
timestamp 1698431365
transform 1 0 36624 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_354
timestamp 1698431365
transform 1 0 44464 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_34_355
timestamp 1698431365
transform 1 0 52304 0 1 38304
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_356
timestamp 1698431365
transform 1 0 9184 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_357
timestamp 1698431365
transform 1 0 17024 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_358
timestamp 1698431365
transform 1 0 24864 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_359
timestamp 1698431365
transform 1 0 32704 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_360
timestamp 1698431365
transform 1 0 40544 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_361
timestamp 1698431365
transform 1 0 48384 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_35_362
timestamp 1698431365
transform 1 0 56224 0 -1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_363
timestamp 1698431365
transform 1 0 5264 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_364
timestamp 1698431365
transform 1 0 13104 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_365
timestamp 1698431365
transform 1 0 20944 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_366
timestamp 1698431365
transform 1 0 28784 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_367
timestamp 1698431365
transform 1 0 36624 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_368
timestamp 1698431365
transform 1 0 44464 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_36_369
timestamp 1698431365
transform 1 0 52304 0 1 40320
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_370
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_371
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_372
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_373
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_374
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_375
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_37_376
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_377
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_378
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_379
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_380
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_381
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_382
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_38_383
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_384
timestamp 1698431365
transform 1 0 9184 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_385
timestamp 1698431365
transform 1 0 17024 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_386
timestamp 1698431365
transform 1 0 24864 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_387
timestamp 1698431365
transform 1 0 32704 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_388
timestamp 1698431365
transform 1 0 40544 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_389
timestamp 1698431365
transform 1 0 48384 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_39_390
timestamp 1698431365
transform 1 0 56224 0 -1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_391
timestamp 1698431365
transform 1 0 5264 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_392
timestamp 1698431365
transform 1 0 13104 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_393
timestamp 1698431365
transform 1 0 20944 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_394
timestamp 1698431365
transform 1 0 28784 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_395
timestamp 1698431365
transform 1 0 36624 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_396
timestamp 1698431365
transform 1 0 44464 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_40_397
timestamp 1698431365
transform 1 0 52304 0 1 44352
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_398
timestamp 1698431365
transform 1 0 9184 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_399
timestamp 1698431365
transform 1 0 17024 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_400
timestamp 1698431365
transform 1 0 24864 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_401
timestamp 1698431365
transform 1 0 32704 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_402
timestamp 1698431365
transform 1 0 40544 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_403
timestamp 1698431365
transform 1 0 48384 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_41_404
timestamp 1698431365
transform 1 0 56224 0 -1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_405
timestamp 1698431365
transform 1 0 5264 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_406
timestamp 1698431365
transform 1 0 13104 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_407
timestamp 1698431365
transform 1 0 20944 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_408
timestamp 1698431365
transform 1 0 28784 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_409
timestamp 1698431365
transform 1 0 36624 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_410
timestamp 1698431365
transform 1 0 44464 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_42_411
timestamp 1698431365
transform 1 0 52304 0 1 46368
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_412
timestamp 1698431365
transform 1 0 9184 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_413
timestamp 1698431365
transform 1 0 17024 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_414
timestamp 1698431365
transform 1 0 24864 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_415
timestamp 1698431365
transform 1 0 32704 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_416
timestamp 1698431365
transform 1 0 40544 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_417
timestamp 1698431365
transform 1 0 48384 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_43_418
timestamp 1698431365
transform 1 0 56224 0 -1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_419
timestamp 1698431365
transform 1 0 5264 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_420
timestamp 1698431365
transform 1 0 13104 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_421
timestamp 1698431365
transform 1 0 20944 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_422
timestamp 1698431365
transform 1 0 28784 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_423
timestamp 1698431365
transform 1 0 36624 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_424
timestamp 1698431365
transform 1 0 44464 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_44_425
timestamp 1698431365
transform 1 0 52304 0 1 48384
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_426
timestamp 1698431365
transform 1 0 9184 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_427
timestamp 1698431365
transform 1 0 17024 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_428
timestamp 1698431365
transform 1 0 24864 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_429
timestamp 1698431365
transform 1 0 32704 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_430
timestamp 1698431365
transform 1 0 40544 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_431
timestamp 1698431365
transform 1 0 48384 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_45_432
timestamp 1698431365
transform 1 0 56224 0 -1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_433
timestamp 1698431365
transform 1 0 5264 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_434
timestamp 1698431365
transform 1 0 13104 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_435
timestamp 1698431365
transform 1 0 20944 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_436
timestamp 1698431365
transform 1 0 28784 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_437
timestamp 1698431365
transform 1 0 36624 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_438
timestamp 1698431365
transform 1 0 44464 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_46_439
timestamp 1698431365
transform 1 0 52304 0 1 50400
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_440
timestamp 1698431365
transform 1 0 9184 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_441
timestamp 1698431365
transform 1 0 17024 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_442
timestamp 1698431365
transform 1 0 24864 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_443
timestamp 1698431365
transform 1 0 32704 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_444
timestamp 1698431365
transform 1 0 40544 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_445
timestamp 1698431365
transform 1 0 48384 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_47_446
timestamp 1698431365
transform 1 0 56224 0 -1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_447
timestamp 1698431365
transform 1 0 5264 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_448
timestamp 1698431365
transform 1 0 13104 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_449
timestamp 1698431365
transform 1 0 20944 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_450
timestamp 1698431365
transform 1 0 28784 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_451
timestamp 1698431365
transform 1 0 36624 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_452
timestamp 1698431365
transform 1 0 44464 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_48_453
timestamp 1698431365
transform 1 0 52304 0 1 52416
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_454
timestamp 1698431365
transform 1 0 9184 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_455
timestamp 1698431365
transform 1 0 17024 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_456
timestamp 1698431365
transform 1 0 24864 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_457
timestamp 1698431365
transform 1 0 32704 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_458
timestamp 1698431365
transform 1 0 40544 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_459
timestamp 1698431365
transform 1 0 48384 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_49_460
timestamp 1698431365
transform 1 0 56224 0 -1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_461
timestamp 1698431365
transform 1 0 5264 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_462
timestamp 1698431365
transform 1 0 13104 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_463
timestamp 1698431365
transform 1 0 20944 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_464
timestamp 1698431365
transform 1 0 28784 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_465
timestamp 1698431365
transform 1 0 36624 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_466
timestamp 1698431365
transform 1 0 44464 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_50_467
timestamp 1698431365
transform 1 0 52304 0 1 54432
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_468
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_469
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_470
timestamp 1698431365
transform 1 0 12768 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_471
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_472
timestamp 1698431365
transform 1 0 20384 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_473
timestamp 1698431365
transform 1 0 24192 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_474
timestamp 1698431365
transform 1 0 28000 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_475
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_476
timestamp 1698431365
transform 1 0 35616 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_477
timestamp 1698431365
transform 1 0 39424 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_478
timestamp 1698431365
transform 1 0 43232 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_479
timestamp 1698431365
transform 1 0 47040 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_480
timestamp 1698431365
transform 1 0 50848 0 -1 56448
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_51_481
timestamp 1698431365
transform 1 0 54656 0 -1 56448
box -86 -90 310 1098
<< labels >>
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 44352 800 44464 0 FreeSans 448 0 0 0 in[0]
port 1 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 in[10]
port 2 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 in[11]
port 3 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 in[12]
port 4 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 in[13]
port 5 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 in[14]
port 6 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 in[15]
port 7 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 in[16]
port 8 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 in[17]
port 9 nsew signal input
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 in[1]
port 10 nsew signal input
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 in[2]
port 11 nsew signal input
flabel metal2 s 27552 59200 27664 60000 0 FreeSans 448 90 0 0 in[3]
port 12 nsew signal input
flabel metal2 s 29568 59200 29680 60000 0 FreeSans 448 90 0 0 in[4]
port 13 nsew signal input
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 in[5]
port 14 nsew signal input
flabel metal3 s 0 38976 800 39088 0 FreeSans 448 0 0 0 in[6]
port 15 nsew signal input
flabel metal3 s 0 37632 800 37744 0 FreeSans 448 0 0 0 in[7]
port 16 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 in[8]
port 17 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 in[9]
port 18 nsew signal input
flabel metal3 s 0 32256 800 32368 0 FreeSans 448 0 0 0 out[0]
port 19 nsew signal tristate
flabel metal3 s 0 51744 800 51856 0 FreeSans 448 0 0 0 out[10]
port 20 nsew signal tristate
flabel metal3 s 0 6720 800 6832 0 FreeSans 448 0 0 0 out[11]
port 21 nsew signal tristate
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 out[1]
port 22 nsew signal tristate
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 out[2]
port 23 nsew signal tristate
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 out[3]
port 24 nsew signal tristate
flabel metal3 s 0 29568 800 29680 0 FreeSans 448 0 0 0 out[4]
port 25 nsew signal tristate
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 out[5]
port 26 nsew signal tristate
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 out[6]
port 27 nsew signal tristate
flabel metal3 s 0 34272 800 34384 0 FreeSans 448 0 0 0 out[7]
port 28 nsew signal tristate
flabel metal3 s 0 6048 800 6160 0 FreeSans 448 0 0 0 out[8]
port 29 nsew signal tristate
flabel metal3 s 59200 53760 60000 53872 0 FreeSans 448 0 0 0 out[9]
port 30 nsew signal tristate
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 rst_n
port 31 nsew signal input
flabel metal4 s 4448 3972 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 35168 3972 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 19808 3972 20128 56508 0 FreeSans 1280 90 0 0 vss
port 33 nsew ground bidirectional
flabel metal4 s 50528 3972 50848 56508 0 FreeSans 1280 90 0 0 vss
port 33 nsew ground bidirectional
rlabel metal1 29960 55440 29960 55440 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal3 27496 36008 27496 36008 0 _000_
rlabel metal2 29512 34216 29512 34216 0 _001_
rlabel metal2 30072 35560 30072 35560 0 _002_
rlabel metal3 26320 35896 26320 35896 0 _003_
rlabel metal2 24024 33600 24024 33600 0 _004_
rlabel metal2 22680 34440 22680 34440 0 _005_
rlabel metal2 23128 37856 23128 37856 0 _006_
rlabel metal2 17416 41384 17416 41384 0 _007_
rlabel metal2 18200 43820 18200 43820 0 _008_
rlabel metal2 22008 41048 22008 41048 0 _009_
rlabel metal2 18816 40600 18816 40600 0 _010_
rlabel metal2 19544 39536 19544 39536 0 _011_
rlabel metal3 13328 35896 13328 35896 0 _012_
rlabel metal2 19712 31976 19712 31976 0 _013_
rlabel metal2 16632 35056 16632 35056 0 _014_
rlabel metal3 16968 36568 16968 36568 0 _015_
rlabel metal2 16184 34384 16184 34384 0 _016_
rlabel metal2 27776 29960 27776 29960 0 _017_
rlabel metal2 26040 30408 26040 30408 0 _018_
rlabel metal2 34384 21784 34384 21784 0 _019_
rlabel metal2 49784 21560 49784 21560 0 _020_
rlabel metal3 30688 20664 30688 20664 0 _021_
rlabel metal2 34720 18536 34720 18536 0 _022_
rlabel metal2 22960 5656 22960 5656 0 _023_
rlabel metal2 25032 16688 25032 16688 0 _024_
rlabel metal2 29848 18144 29848 18144 0 _025_
rlabel metal3 26684 21672 26684 21672 0 _026_
rlabel metal2 21896 7028 21896 7028 0 _027_
rlabel metal2 23800 16688 23800 16688 0 _028_
rlabel metal2 24528 16632 24528 16632 0 _029_
rlabel metal2 20776 18200 20776 18200 0 _030_
rlabel metal2 23576 18200 23576 18200 0 _031_
rlabel metal3 46704 33880 46704 33880 0 _032_
rlabel metal3 24808 11592 24808 11592 0 _033_
rlabel metal2 25256 24640 25256 24640 0 _034_
rlabel metal3 33264 30632 33264 30632 0 _035_
rlabel metal2 49336 29680 49336 29680 0 _036_
rlabel metal2 23800 26600 23800 26600 0 _037_
rlabel metal2 24080 26824 24080 26824 0 _038_
rlabel metal2 32200 28168 32200 28168 0 _039_
rlabel metal2 24248 26432 24248 26432 0 _040_
rlabel metal2 25592 25704 25592 25704 0 _041_
rlabel metal2 25256 25984 25256 25984 0 _042_
rlabel metal2 23240 25536 23240 25536 0 _043_
rlabel metal2 22512 21000 22512 21000 0 _044_
rlabel metal2 22904 25816 22904 25816 0 _045_
rlabel metal2 45248 28504 45248 28504 0 _046_
rlabel metal2 30072 28840 30072 28840 0 _047_
rlabel metal3 25788 27720 25788 27720 0 _048_
rlabel metal3 23744 29960 23744 29960 0 _049_
rlabel metal3 23296 7672 23296 7672 0 _050_
rlabel metal2 22344 11088 22344 11088 0 _051_
rlabel metal2 24696 25816 24696 25816 0 _052_
rlabel metal2 24024 27328 24024 27328 0 _053_
rlabel metal2 23800 29120 23800 29120 0 _054_
rlabel metal2 22960 32536 22960 32536 0 _055_
rlabel metal3 18648 31752 18648 31752 0 _056_
rlabel metal3 15232 33768 15232 33768 0 _057_
rlabel metal2 26376 32872 26376 32872 0 _058_
rlabel metal2 27720 30576 27720 30576 0 _059_
rlabel metal3 40096 38696 40096 38696 0 _060_
rlabel metal2 46536 39368 46536 39368 0 _061_
rlabel metal3 44632 38696 44632 38696 0 _062_
rlabel metal2 50904 42280 50904 42280 0 _063_
rlabel metal2 47544 31752 47544 31752 0 _064_
rlabel metal2 51128 40880 51128 40880 0 _065_
rlabel metal2 46760 39480 46760 39480 0 _066_
rlabel metal2 51576 34832 51576 34832 0 _067_
rlabel metal2 46088 37576 46088 37576 0 _068_
rlabel metal2 46032 39816 46032 39816 0 _069_
rlabel metal3 48720 39816 48720 39816 0 _070_
rlabel metal2 45528 36568 45528 36568 0 _071_
rlabel metal2 45192 34776 45192 34776 0 _072_
rlabel metal2 23912 32088 23912 32088 0 _073_
rlabel metal2 45752 25200 45752 25200 0 _074_
rlabel metal2 26376 26740 26376 26740 0 _075_
rlabel metal2 26936 10136 26936 10136 0 _076_
rlabel metal2 41272 9464 41272 9464 0 _077_
rlabel metal3 36736 15624 36736 15624 0 _078_
rlabel metal3 30744 7784 30744 7784 0 _079_
rlabel metal2 26376 28784 26376 28784 0 _080_
rlabel metal2 33656 24024 33656 24024 0 _081_
rlabel metal2 40376 31472 40376 31472 0 _082_
rlabel metal2 36064 26488 36064 26488 0 _083_
rlabel metal2 33880 26096 33880 26096 0 _084_
rlabel metal3 31248 22456 31248 22456 0 _085_
rlabel metal2 29960 25256 29960 25256 0 _086_
rlabel metal2 42896 26712 42896 26712 0 _087_
rlabel metal2 42280 26152 42280 26152 0 _088_
rlabel metal2 30408 25704 30408 25704 0 _089_
rlabel metal2 25480 28056 25480 28056 0 _090_
rlabel metal2 25368 31920 25368 31920 0 _091_
rlabel metal2 24584 30352 24584 30352 0 _092_
rlabel metal2 15960 31472 15960 31472 0 _093_
rlabel metal2 32872 12152 32872 12152 0 _094_
rlabel metal2 42616 21448 42616 21448 0 _095_
rlabel metal2 32200 11144 32200 11144 0 _096_
rlabel metal2 25592 26600 25592 26600 0 _097_
rlabel metal2 28056 42280 28056 42280 0 _098_
rlabel metal2 25032 26656 25032 26656 0 _099_
rlabel metal2 26152 22400 26152 22400 0 _100_
rlabel metal2 21896 26376 21896 26376 0 _101_
rlabel metal3 20328 26712 20328 26712 0 _102_
rlabel metal2 25200 28168 25200 28168 0 _103_
rlabel metal2 31472 21784 31472 21784 0 _104_
rlabel metal3 31136 24584 31136 24584 0 _105_
rlabel metal2 30128 26712 30128 26712 0 _106_
rlabel metal2 26152 25872 26152 25872 0 _107_
rlabel metal2 26824 25760 26824 25760 0 _108_
rlabel metal2 26936 25984 26936 25984 0 _109_
rlabel metal2 32704 31864 32704 31864 0 _110_
rlabel metal3 30968 32872 30968 32872 0 _111_
rlabel metal2 39928 34272 39928 34272 0 _112_
rlabel metal2 39368 35056 39368 35056 0 _113_
rlabel metal3 31304 26712 31304 26712 0 _114_
rlabel metal2 30688 27048 30688 27048 0 _115_
rlabel metal2 36568 26264 36568 26264 0 _116_
rlabel metal2 33768 26852 33768 26852 0 _117_
rlabel metal2 30576 41720 30576 41720 0 _118_
rlabel metal2 33544 30800 33544 30800 0 _119_
rlabel metal2 29904 39704 29904 39704 0 _120_
rlabel metal2 33936 28728 33936 28728 0 _121_
rlabel metal2 51016 21056 51016 21056 0 _122_
rlabel metal3 37072 26712 37072 26712 0 _123_
rlabel metal2 34664 28392 34664 28392 0 _124_
rlabel metal2 31080 28672 31080 28672 0 _125_
rlabel metal2 30744 28784 30744 28784 0 _126_
rlabel metal2 25256 29680 25256 29680 0 _127_
rlabel metal2 18312 30520 18312 30520 0 _128_
rlabel metal2 36232 19544 36232 19544 0 _129_
rlabel metal3 41328 21672 41328 21672 0 _130_
rlabel metal2 41608 18984 41608 18984 0 _131_
rlabel metal2 37016 39368 37016 39368 0 _132_
rlabel metal2 26264 23520 26264 23520 0 _133_
rlabel metal2 25816 25872 25816 25872 0 _134_
rlabel metal2 26152 26852 26152 26852 0 _135_
rlabel metal2 49784 35224 49784 35224 0 _136_
rlabel metal2 51688 30744 51688 30744 0 _137_
rlabel metal3 48944 24360 48944 24360 0 _138_
rlabel metal2 53928 33152 53928 33152 0 _139_
rlabel metal2 49672 34216 49672 34216 0 _140_
rlabel metal2 51912 35616 51912 35616 0 _141_
rlabel metal2 53256 34328 53256 34328 0 _142_
rlabel metal2 49112 34160 49112 34160 0 _143_
rlabel metal2 48664 33096 48664 33096 0 _144_
rlabel metal2 27160 30632 27160 30632 0 _145_
rlabel metal2 14504 30576 14504 30576 0 _146_
rlabel metal2 14952 30240 14952 30240 0 _147_
rlabel metal2 41048 23464 41048 23464 0 _148_
rlabel metal3 40656 43848 40656 43848 0 _149_
rlabel metal2 42504 43764 42504 43764 0 _150_
rlabel metal2 41608 38808 41608 38808 0 _151_
rlabel metal2 40152 29680 40152 29680 0 _152_
rlabel metal3 23576 26824 23576 26824 0 _153_
rlabel metal3 26376 38808 26376 38808 0 _154_
rlabel metal2 24808 29344 24808 29344 0 _155_
rlabel metal2 32536 21784 32536 21784 0 _156_
rlabel metal2 31192 24920 31192 24920 0 _157_
rlabel metal2 25928 23856 25928 23856 0 _158_
rlabel metal3 28784 25032 28784 25032 0 _159_
rlabel metal3 33768 31864 33768 31864 0 _160_
rlabel metal2 31416 28672 31416 28672 0 _161_
rlabel metal2 29736 28448 29736 28448 0 _162_
rlabel metal2 33768 24472 33768 24472 0 _163_
rlabel metal2 33152 28728 33152 28728 0 _164_
rlabel metal2 33208 32088 33208 32088 0 _165_
rlabel metal2 32872 29792 32872 29792 0 _166_
rlabel metal2 39480 26768 39480 26768 0 _167_
rlabel metal2 33544 28448 33544 28448 0 _168_
rlabel metal3 31584 28728 31584 28728 0 _169_
rlabel metal2 24248 29512 24248 29512 0 _170_
rlabel metal3 15092 28616 15092 28616 0 _171_
rlabel metal2 25816 36904 25816 36904 0 _172_
rlabel metal2 35560 39872 35560 39872 0 _173_
rlabel metal2 35000 40544 35000 40544 0 _174_
rlabel metal2 26040 38024 26040 38024 0 _175_
rlabel metal2 25480 38248 25480 38248 0 _176_
rlabel metal2 25536 31864 25536 31864 0 _177_
rlabel metal2 51912 28896 51912 28896 0 _178_
rlabel metal2 46872 22680 46872 22680 0 _179_
rlabel metal2 55160 23072 55160 23072 0 _180_
rlabel metal3 52248 27944 52248 27944 0 _181_
rlabel metal2 51016 24752 51016 24752 0 _182_
rlabel metal2 50904 29456 50904 29456 0 _183_
rlabel metal2 51240 24528 51240 24528 0 _184_
rlabel metal2 50456 22400 50456 22400 0 _185_
rlabel metal2 50232 24976 50232 24976 0 _186_
rlabel metal2 48664 30240 48664 30240 0 _187_
rlabel metal2 26264 31360 26264 31360 0 _188_
rlabel metal2 19208 30800 19208 30800 0 _189_
rlabel metal3 42056 15848 42056 15848 0 _190_
rlabel metal2 40768 42616 40768 42616 0 _191_
rlabel metal2 29064 29848 29064 29848 0 _192_
rlabel metal2 22680 29288 22680 29288 0 _193_
rlabel metal3 26656 30632 26656 30632 0 _194_
rlabel metal3 30072 20888 30072 20888 0 _195_
rlabel metal2 29904 24696 29904 24696 0 _196_
rlabel metal2 24920 25368 24920 25368 0 _197_
rlabel metal2 26040 26432 26040 26432 0 _198_
rlabel metal3 31416 30072 31416 30072 0 _199_
rlabel metal2 30296 28392 30296 28392 0 _200_
rlabel metal2 29624 28784 29624 28784 0 _201_
rlabel metal2 32592 25928 32592 25928 0 _202_
rlabel metal2 33376 29736 33376 29736 0 _203_
rlabel metal2 33096 31976 33096 31976 0 _204_
rlabel metal2 33096 30128 33096 30128 0 _205_
rlabel metal2 35784 30296 35784 30296 0 _206_
rlabel metal3 34608 29736 34608 29736 0 _207_
rlabel metal3 31584 29736 31584 29736 0 _208_
rlabel metal2 25704 30408 25704 30408 0 _209_
rlabel metal2 18984 33376 18984 33376 0 _210_
rlabel metal2 29848 40152 29848 40152 0 _211_
rlabel metal3 28504 39928 28504 39928 0 _212_
rlabel metal2 28560 38808 28560 38808 0 _213_
rlabel metal2 27496 38360 27496 38360 0 _214_
rlabel metal2 28000 38920 28000 38920 0 _215_
rlabel metal2 47656 23072 47656 23072 0 _216_
rlabel metal2 47656 24584 47656 24584 0 _217_
rlabel metal2 47432 25088 47432 25088 0 _218_
rlabel metal2 51912 22512 51912 22512 0 _219_
rlabel metal3 52136 21336 52136 21336 0 _220_
rlabel metal2 50904 24360 50904 24360 0 _221_
rlabel metal2 45864 26096 45864 26096 0 _222_
rlabel metal2 26712 31864 26712 31864 0 _223_
rlabel metal2 18424 33264 18424 33264 0 _224_
rlabel metal2 19600 34664 19600 34664 0 _225_
rlabel metal3 23016 31864 23016 31864 0 _226_
rlabel via1 21336 31755 21336 31755 0 _227_
rlabel metal3 20608 31864 20608 31864 0 _228_
rlabel metal2 18760 31864 18760 31864 0 _229_
rlabel metal2 17248 31080 17248 31080 0 _230_
rlabel metal2 17640 33096 17640 33096 0 _231_
rlabel metal2 12824 32592 12824 32592 0 _232_
rlabel metal3 23800 36680 23800 36680 0 _233_
rlabel metal2 22456 35672 22456 35672 0 _234_
rlabel metal2 22232 35448 22232 35448 0 _235_
rlabel metal2 22904 36008 22904 36008 0 _236_
rlabel metal3 25032 35784 25032 35784 0 _237_
rlabel metal2 20720 38696 20720 38696 0 _238_
rlabel metal2 24248 36624 24248 36624 0 _239_
rlabel metal2 21672 39424 21672 39424 0 _240_
rlabel metal3 17136 35784 17136 35784 0 _241_
rlabel metal3 20328 36904 20328 36904 0 _242_
rlabel metal3 9576 34552 9576 34552 0 _243_
rlabel metal2 20664 6664 20664 6664 0 cm_inst.cc_inst.in\[0\]
rlabel metal2 20496 5768 20496 5768 0 cm_inst.cc_inst.in\[1\]
rlabel metal2 20216 6160 20216 6160 0 cm_inst.cc_inst.in\[2\]
rlabel metal2 25928 5040 25928 5040 0 cm_inst.cc_inst.in\[3\]
rlabel metal2 24696 7840 24696 7840 0 cm_inst.cc_inst.in\[4\]
rlabel metal3 22792 24696 22792 24696 0 cm_inst.cc_inst.in\[5\]
rlabel metal2 21784 15792 21784 15792 0 cm_inst.cc_inst.out_notouch_\[0\]
rlabel metal2 45696 33880 45696 33880 0 cm_inst.cc_inst.out_notouch_\[100\]
rlabel metal2 54152 29456 54152 29456 0 cm_inst.cc_inst.out_notouch_\[101\]
rlabel metal2 45192 30240 45192 30240 0 cm_inst.cc_inst.out_notouch_\[102\]
rlabel metal2 49224 21728 49224 21728 0 cm_inst.cc_inst.out_notouch_\[103\]
rlabel metal2 28616 17640 28616 17640 0 cm_inst.cc_inst.out_notouch_\[104\]
rlabel metal2 43960 36120 43960 36120 0 cm_inst.cc_inst.out_notouch_\[105\]
rlabel metal2 40824 36344 40824 36344 0 cm_inst.cc_inst.out_notouch_\[106\]
rlabel metal2 50904 35224 50904 35224 0 cm_inst.cc_inst.out_notouch_\[107\]
rlabel metal3 45528 32984 45528 32984 0 cm_inst.cc_inst.out_notouch_\[108\]
rlabel metal2 49896 29288 49896 29288 0 cm_inst.cc_inst.out_notouch_\[109\]
rlabel metal2 33544 33096 33544 33096 0 cm_inst.cc_inst.out_notouch_\[10\]
rlabel metal2 46200 29288 46200 29288 0 cm_inst.cc_inst.out_notouch_\[110\]
rlabel metal2 48776 21364 48776 21364 0 cm_inst.cc_inst.out_notouch_\[111\]
rlabel metal2 46648 18872 46648 18872 0 cm_inst.cc_inst.out_notouch_\[112\]
rlabel metal2 39816 36960 39816 36960 0 cm_inst.cc_inst.out_notouch_\[113\]
rlabel metal2 38024 36400 38024 36400 0 cm_inst.cc_inst.out_notouch_\[114\]
rlabel metal3 47600 35784 47600 35784 0 cm_inst.cc_inst.out_notouch_\[115\]
rlabel metal2 42840 34272 42840 34272 0 cm_inst.cc_inst.out_notouch_\[116\]
rlabel metal2 51352 30128 51352 30128 0 cm_inst.cc_inst.out_notouch_\[117\]
rlabel metal2 42448 29848 42448 29848 0 cm_inst.cc_inst.out_notouch_\[118\]
rlabel metal2 46648 23016 46648 23016 0 cm_inst.cc_inst.out_notouch_\[119\]
rlabel metal2 54376 33936 54376 33936 0 cm_inst.cc_inst.out_notouch_\[11\]
rlabel metal2 30184 17136 30184 17136 0 cm_inst.cc_inst.out_notouch_\[120\]
rlabel metal2 41608 38248 41608 38248 0 cm_inst.cc_inst.out_notouch_\[121\]
rlabel metal2 38808 35784 38808 35784 0 cm_inst.cc_inst.out_notouch_\[122\]
rlabel metal2 49448 36176 49448 36176 0 cm_inst.cc_inst.out_notouch_\[123\]
rlabel metal2 43512 34216 43512 34216 0 cm_inst.cc_inst.out_notouch_\[124\]
rlabel metal2 52024 30128 52024 30128 0 cm_inst.cc_inst.out_notouch_\[125\]
rlabel metal2 43064 30184 43064 30184 0 cm_inst.cc_inst.out_notouch_\[126\]
rlabel metal2 47320 22232 47320 22232 0 cm_inst.cc_inst.out_notouch_\[127\]
rlabel metal2 22456 10136 22456 10136 0 cm_inst.cc_inst.out_notouch_\[128\]
rlabel metal2 35840 6888 35840 6888 0 cm_inst.cc_inst.out_notouch_\[129\]
rlabel metal3 34216 33768 34216 33768 0 cm_inst.cc_inst.out_notouch_\[12\]
rlabel metal2 44072 9296 44072 9296 0 cm_inst.cc_inst.out_notouch_\[130\]
rlabel metal3 43512 20440 43512 20440 0 cm_inst.cc_inst.out_notouch_\[131\]
rlabel metal2 43792 44072 43792 44072 0 cm_inst.cc_inst.out_notouch_\[132\]
rlabel metal2 35112 43820 35112 43820 0 cm_inst.cc_inst.out_notouch_\[133\]
rlabel metal2 42168 45640 42168 45640 0 cm_inst.cc_inst.out_notouch_\[134\]
rlabel metal2 28728 45724 28728 45724 0 cm_inst.cc_inst.out_notouch_\[135\]
rlabel metal2 23464 11032 23464 11032 0 cm_inst.cc_inst.out_notouch_\[136\]
rlabel metal2 35168 7560 35168 7560 0 cm_inst.cc_inst.out_notouch_\[137\]
rlabel metal2 43064 10248 43064 10248 0 cm_inst.cc_inst.out_notouch_\[138\]
rlabel metal2 42728 19040 42728 19040 0 cm_inst.cc_inst.out_notouch_\[139\]
rlabel metal2 51576 20916 51576 20916 0 cm_inst.cc_inst.out_notouch_\[13\]
rlabel metal2 43064 45248 43064 45248 0 cm_inst.cc_inst.out_notouch_\[140\]
rlabel metal2 33656 44156 33656 44156 0 cm_inst.cc_inst.out_notouch_\[141\]
rlabel metal2 42056 44632 42056 44632 0 cm_inst.cc_inst.out_notouch_\[142\]
rlabel metal2 28616 42392 28616 42392 0 cm_inst.cc_inst.out_notouch_\[143\]
rlabel metal3 20748 10472 20748 10472 0 cm_inst.cc_inst.out_notouch_\[144\]
rlabel metal2 32872 7168 32872 7168 0 cm_inst.cc_inst.out_notouch_\[145\]
rlabel metal3 40600 9576 40600 9576 0 cm_inst.cc_inst.out_notouch_\[146\]
rlabel metal2 40600 18760 40600 18760 0 cm_inst.cc_inst.out_notouch_\[147\]
rlabel metal2 40936 45080 40936 45080 0 cm_inst.cc_inst.out_notouch_\[148\]
rlabel metal2 31752 43232 31752 43232 0 cm_inst.cc_inst.out_notouch_\[149\]
rlabel metal2 33208 38668 33208 38668 0 cm_inst.cc_inst.out_notouch_\[14\]
rlabel metal2 39704 43232 39704 43232 0 cm_inst.cc_inst.out_notouch_\[150\]
rlabel metal2 25816 45164 25816 45164 0 cm_inst.cc_inst.out_notouch_\[151\]
rlabel metal3 21560 10584 21560 10584 0 cm_inst.cc_inst.out_notouch_\[152\]
rlabel metal2 32480 5768 32480 5768 0 cm_inst.cc_inst.out_notouch_\[153\]
rlabel metal2 41160 8904 41160 8904 0 cm_inst.cc_inst.out_notouch_\[154\]
rlabel metal2 41272 19040 41272 19040 0 cm_inst.cc_inst.out_notouch_\[155\]
rlabel metal2 41608 44744 41608 44744 0 cm_inst.cc_inst.out_notouch_\[156\]
rlabel metal2 31864 44968 31864 44968 0 cm_inst.cc_inst.out_notouch_\[157\]
rlabel metal2 40096 45640 40096 45640 0 cm_inst.cc_inst.out_notouch_\[158\]
rlabel metal3 26768 41944 26768 41944 0 cm_inst.cc_inst.out_notouch_\[159\]
rlabel metal2 54040 18816 54040 18816 0 cm_inst.cc_inst.out_notouch_\[15\]
rlabel metal2 24360 6048 24360 6048 0 cm_inst.cc_inst.out_notouch_\[160\]
rlabel metal2 28728 8680 28728 8680 0 cm_inst.cc_inst.out_notouch_\[161\]
rlabel metal2 35560 10304 35560 10304 0 cm_inst.cc_inst.out_notouch_\[162\]
rlabel metal3 38808 15736 38808 15736 0 cm_inst.cc_inst.out_notouch_\[163\]
rlabel metal2 44520 13328 44520 13328 0 cm_inst.cc_inst.out_notouch_\[164\]
rlabel metal2 42392 40320 42392 40320 0 cm_inst.cc_inst.out_notouch_\[165\]
rlabel metal2 44184 16072 44184 16072 0 cm_inst.cc_inst.out_notouch_\[166\]
rlabel metal2 35896 41440 35896 41440 0 cm_inst.cc_inst.out_notouch_\[167\]
rlabel metal2 23688 6496 23688 6496 0 cm_inst.cc_inst.out_notouch_\[168\]
rlabel metal2 28280 9184 28280 9184 0 cm_inst.cc_inst.out_notouch_\[169\]
rlabel metal2 19040 15624 19040 15624 0 cm_inst.cc_inst.out_notouch_\[16\]
rlabel metal2 34552 10640 34552 10640 0 cm_inst.cc_inst.out_notouch_\[170\]
rlabel metal2 38920 15176 38920 15176 0 cm_inst.cc_inst.out_notouch_\[171\]
rlabel metal2 47768 13160 47768 13160 0 cm_inst.cc_inst.out_notouch_\[172\]
rlabel metal2 46536 44240 46536 44240 0 cm_inst.cc_inst.out_notouch_\[173\]
rlabel metal2 44968 15792 44968 15792 0 cm_inst.cc_inst.out_notouch_\[174\]
rlabel metal2 34888 47936 34888 47936 0 cm_inst.cc_inst.out_notouch_\[175\]
rlabel metal2 21504 5656 21504 5656 0 cm_inst.cc_inst.out_notouch_\[176\]
rlabel metal2 25928 10192 25928 10192 0 cm_inst.cc_inst.out_notouch_\[177\]
rlabel metal2 32704 11592 32704 11592 0 cm_inst.cc_inst.out_notouch_\[178\]
rlabel metal2 36792 16240 36792 16240 0 cm_inst.cc_inst.out_notouch_\[179\]
rlabel metal2 49560 40208 49560 40208 0 cm_inst.cc_inst.out_notouch_\[17\]
rlabel metal2 41720 14224 41720 14224 0 cm_inst.cc_inst.out_notouch_\[180\]
rlabel metal2 40936 39984 40936 39984 0 cm_inst.cc_inst.out_notouch_\[181\]
rlabel metal2 41384 15848 41384 15848 0 cm_inst.cc_inst.out_notouch_\[182\]
rlabel metal2 33096 41160 33096 41160 0 cm_inst.cc_inst.out_notouch_\[183\]
rlabel metal2 22232 5992 22232 5992 0 cm_inst.cc_inst.out_notouch_\[184\]
rlabel metal2 25704 7532 25704 7532 0 cm_inst.cc_inst.out_notouch_\[185\]
rlabel metal2 32536 9912 32536 9912 0 cm_inst.cc_inst.out_notouch_\[186\]
rlabel metal3 36848 15736 36848 15736 0 cm_inst.cc_inst.out_notouch_\[187\]
rlabel metal2 42392 13776 42392 13776 0 cm_inst.cc_inst.out_notouch_\[188\]
rlabel metal2 41552 39928 41552 39928 0 cm_inst.cc_inst.out_notouch_\[189\]
rlabel metal2 33544 26544 33544 26544 0 cm_inst.cc_inst.out_notouch_\[18\]
rlabel metal2 42112 15736 42112 15736 0 cm_inst.cc_inst.out_notouch_\[190\]
rlabel metal2 34048 40040 34048 40040 0 cm_inst.cc_inst.out_notouch_\[191\]
rlabel metal3 20440 20552 20440 20552 0 cm_inst.cc_inst.out_notouch_\[192\]
rlabel metal2 43176 26320 43176 26320 0 cm_inst.cc_inst.out_notouch_\[193\]
rlabel metal2 16968 25704 16968 25704 0 cm_inst.cc_inst.out_notouch_\[194\]
rlabel metal2 14616 24808 14616 24808 0 cm_inst.cc_inst.out_notouch_\[195\]
rlabel metal3 22288 27384 22288 27384 0 cm_inst.cc_inst.out_notouch_\[196\]
rlabel metal2 27160 38976 27160 38976 0 cm_inst.cc_inst.out_notouch_\[197\]
rlabel metal2 21672 28168 21672 28168 0 cm_inst.cc_inst.out_notouch_\[198\]
rlabel metal3 27048 39816 27048 39816 0 cm_inst.cc_inst.out_notouch_\[199\]
rlabel metal2 52024 33768 52024 33768 0 cm_inst.cc_inst.out_notouch_\[19\]
rlabel metal2 52360 41048 52360 41048 0 cm_inst.cc_inst.out_notouch_\[1\]
rlabel metal3 22120 20496 22120 20496 0 cm_inst.cc_inst.out_notouch_\[200\]
rlabel metal2 42728 27048 42728 27048 0 cm_inst.cc_inst.out_notouch_\[201\]
rlabel metal2 16408 24808 16408 24808 0 cm_inst.cc_inst.out_notouch_\[202\]
rlabel metal2 18200 25872 18200 25872 0 cm_inst.cc_inst.out_notouch_\[203\]
rlabel metal2 22120 26544 22120 26544 0 cm_inst.cc_inst.out_notouch_\[204\]
rlabel metal2 26600 39592 26600 39592 0 cm_inst.cc_inst.out_notouch_\[205\]
rlabel metal3 21560 27720 21560 27720 0 cm_inst.cc_inst.out_notouch_\[206\]
rlabel metal2 27496 39592 27496 39592 0 cm_inst.cc_inst.out_notouch_\[207\]
rlabel metal2 21784 24192 21784 24192 0 cm_inst.cc_inst.out_notouch_\[208\]
rlabel metal3 30016 24024 30016 24024 0 cm_inst.cc_inst.out_notouch_\[209\]
rlabel metal2 35560 26264 35560 26264 0 cm_inst.cc_inst.out_notouch_\[20\]
rlabel metal2 49504 21784 49504 21784 0 cm_inst.cc_inst.out_notouch_\[21\]
rlabel metal2 33152 26936 33152 26936 0 cm_inst.cc_inst.out_notouch_\[22\]
rlabel metal2 51912 19208 51912 19208 0 cm_inst.cc_inst.out_notouch_\[23\]
rlabel metal2 20216 18144 20216 18144 0 cm_inst.cc_inst.out_notouch_\[24\]
rlabel metal2 50232 40768 50232 40768 0 cm_inst.cc_inst.out_notouch_\[25\]
rlabel metal2 36232 25536 36232 25536 0 cm_inst.cc_inst.out_notouch_\[26\]
rlabel metal2 52920 34216 52920 34216 0 cm_inst.cc_inst.out_notouch_\[27\]
rlabel metal2 33432 24640 33432 24640 0 cm_inst.cc_inst.out_notouch_\[28\]
rlabel metal2 50120 20552 50120 20552 0 cm_inst.cc_inst.out_notouch_\[29\]
rlabel metal2 34104 33152 34104 33152 0 cm_inst.cc_inst.out_notouch_\[2\]
rlabel metal3 31976 25704 31976 25704 0 cm_inst.cc_inst.out_notouch_\[30\]
rlabel metal2 50008 18816 50008 18816 0 cm_inst.cc_inst.out_notouch_\[31\]
rlabel metal2 22568 18592 22568 18592 0 cm_inst.cc_inst.out_notouch_\[32\]
rlabel metal2 47992 40040 47992 40040 0 cm_inst.cc_inst.out_notouch_\[33\]
rlabel metal2 40040 23632 40040 23632 0 cm_inst.cc_inst.out_notouch_\[34\]
rlabel metal2 55832 35840 55832 35840 0 cm_inst.cc_inst.out_notouch_\[35\]
rlabel metal2 41160 26264 41160 26264 0 cm_inst.cc_inst.out_notouch_\[36\]
rlabel metal2 56336 24472 56336 24472 0 cm_inst.cc_inst.out_notouch_\[37\]
rlabel metal2 39144 31192 39144 31192 0 cm_inst.cc_inst.out_notouch_\[38\]
rlabel metal3 56840 22456 56840 22456 0 cm_inst.cc_inst.out_notouch_\[39\]
rlabel metal2 55048 34720 55048 34720 0 cm_inst.cc_inst.out_notouch_\[3\]
rlabel metal2 21840 17640 21840 17640 0 cm_inst.cc_inst.out_notouch_\[40\]
rlabel metal2 47208 40992 47208 40992 0 cm_inst.cc_inst.out_notouch_\[41\]
rlabel metal2 39368 23352 39368 23352 0 cm_inst.cc_inst.out_notouch_\[42\]
rlabel metal3 55160 36624 55160 36624 0 cm_inst.cc_inst.out_notouch_\[43\]
rlabel metal2 40600 25480 40600 25480 0 cm_inst.cc_inst.out_notouch_\[44\]
rlabel metal2 55272 25312 55272 25312 0 cm_inst.cc_inst.out_notouch_\[45\]
rlabel metal2 38472 32144 38472 32144 0 cm_inst.cc_inst.out_notouch_\[46\]
rlabel metal2 55832 23296 55832 23296 0 cm_inst.cc_inst.out_notouch_\[47\]
rlabel metal2 19768 17864 19768 17864 0 cm_inst.cc_inst.out_notouch_\[48\]
rlabel metal2 45080 40712 45080 40712 0 cm_inst.cc_inst.out_notouch_\[49\]
rlabel metal2 34104 34272 34104 34272 0 cm_inst.cc_inst.out_notouch_\[4\]
rlabel metal2 37240 24136 37240 24136 0 cm_inst.cc_inst.out_notouch_\[50\]
rlabel metal2 52584 36680 52584 36680 0 cm_inst.cc_inst.out_notouch_\[51\]
rlabel metal2 38528 25592 38528 25592 0 cm_inst.cc_inst.out_notouch_\[52\]
rlabel metal2 53256 24192 53256 24192 0 cm_inst.cc_inst.out_notouch_\[53\]
rlabel metal2 36344 31360 36344 31360 0 cm_inst.cc_inst.out_notouch_\[54\]
rlabel metal2 53704 21504 53704 21504 0 cm_inst.cc_inst.out_notouch_\[55\]
rlabel metal3 20440 17584 20440 17584 0 cm_inst.cc_inst.out_notouch_\[56\]
rlabel metal3 45360 39928 45360 39928 0 cm_inst.cc_inst.out_notouch_\[57\]
rlabel metal2 37352 23072 37352 23072 0 cm_inst.cc_inst.out_notouch_\[58\]
rlabel metal2 53704 37128 53704 37128 0 cm_inst.cc_inst.out_notouch_\[59\]
rlabel metal2 51912 21392 51912 21392 0 cm_inst.cc_inst.out_notouch_\[5\]
rlabel metal2 39144 26152 39144 26152 0 cm_inst.cc_inst.out_notouch_\[60\]
rlabel metal2 53760 24696 53760 24696 0 cm_inst.cc_inst.out_notouch_\[61\]
rlabel metal2 35784 31808 35784 31808 0 cm_inst.cc_inst.out_notouch_\[62\]
rlabel metal2 53480 22064 53480 22064 0 cm_inst.cc_inst.out_notouch_\[63\]
rlabel metal2 26544 12824 26544 12824 0 cm_inst.cc_inst.out_notouch_\[64\]
rlabel metal2 54712 39648 54712 39648 0 cm_inst.cc_inst.out_notouch_\[65\]
rlabel metal2 24472 24752 24472 24752 0 cm_inst.cc_inst.out_notouch_\[66\]
rlabel metal2 55720 33152 55720 33152 0 cm_inst.cc_inst.out_notouch_\[67\]
rlabel metal3 26264 22568 26264 22568 0 cm_inst.cc_inst.out_notouch_\[68\]
rlabel metal3 55944 27832 55944 27832 0 cm_inst.cc_inst.out_notouch_\[69\]
rlabel metal2 33768 38416 33768 38416 0 cm_inst.cc_inst.out_notouch_\[6\]
rlabel metal2 25816 24304 25816 24304 0 cm_inst.cc_inst.out_notouch_\[70\]
rlabel metal2 52360 16856 52360 16856 0 cm_inst.cc_inst.out_notouch_\[71\]
rlabel metal2 25592 16240 25592 16240 0 cm_inst.cc_inst.out_notouch_\[72\]
rlabel metal2 54936 40936 54936 40936 0 cm_inst.cc_inst.out_notouch_\[73\]
rlabel metal2 23856 25704 23856 25704 0 cm_inst.cc_inst.out_notouch_\[74\]
rlabel metal3 55048 32592 55048 32592 0 cm_inst.cc_inst.out_notouch_\[75\]
rlabel metal2 26376 23072 26376 23072 0 cm_inst.cc_inst.out_notouch_\[76\]
rlabel metal2 54320 27720 54320 27720 0 cm_inst.cc_inst.out_notouch_\[77\]
rlabel metal3 24976 24584 24976 24584 0 cm_inst.cc_inst.out_notouch_\[78\]
rlabel metal2 51688 17024 51688 17024 0 cm_inst.cc_inst.out_notouch_\[79\]
rlabel metal2 54712 19376 54712 19376 0 cm_inst.cc_inst.out_notouch_\[7\]
rlabel metal2 22680 15008 22680 15008 0 cm_inst.cc_inst.out_notouch_\[80\]
rlabel metal2 52976 40040 52976 40040 0 cm_inst.cc_inst.out_notouch_\[81\]
rlabel metal2 31080 24248 31080 24248 0 cm_inst.cc_inst.out_notouch_\[82\]
rlabel metal2 52920 32312 52920 32312 0 cm_inst.cc_inst.out_notouch_\[83\]
rlabel metal2 31304 23632 31304 23632 0 cm_inst.cc_inst.out_notouch_\[84\]
rlabel metal2 52136 27888 52136 27888 0 cm_inst.cc_inst.out_notouch_\[85\]
rlabel metal2 30520 22232 30520 22232 0 cm_inst.cc_inst.out_notouch_\[86\]
rlabel metal2 49560 17808 49560 17808 0 cm_inst.cc_inst.out_notouch_\[87\]
rlabel metal2 24136 16184 24136 16184 0 cm_inst.cc_inst.out_notouch_\[88\]
rlabel metal2 53424 41832 53424 41832 0 cm_inst.cc_inst.out_notouch_\[89\]
rlabel metal2 21112 16016 21112 16016 0 cm_inst.cc_inst.out_notouch_\[8\]
rlabel metal2 31976 21168 31976 21168 0 cm_inst.cc_inst.out_notouch_\[90\]
rlabel metal2 53592 34160 53592 34160 0 cm_inst.cc_inst.out_notouch_\[91\]
rlabel metal2 32872 20384 32872 20384 0 cm_inst.cc_inst.out_notouch_\[92\]
rlabel metal3 52416 27720 52416 27720 0 cm_inst.cc_inst.out_notouch_\[93\]
rlabel metal2 30744 20272 30744 20272 0 cm_inst.cc_inst.out_notouch_\[94\]
rlabel metal2 50232 17192 50232 17192 0 cm_inst.cc_inst.out_notouch_\[95\]
rlabel metal3 29288 16632 29288 16632 0 cm_inst.cc_inst.out_notouch_\[96\]
rlabel metal2 43792 37912 43792 37912 0 cm_inst.cc_inst.out_notouch_\[97\]
rlabel metal2 41160 34832 41160 34832 0 cm_inst.cc_inst.out_notouch_\[98\]
rlabel metal2 51576 36456 51576 36456 0 cm_inst.cc_inst.out_notouch_\[99\]
rlabel metal2 51744 39928 51744 39928 0 cm_inst.cc_inst.out_notouch_\[9\]
rlabel metal3 35616 35784 35616 35784 0 cm_inst.page\[0\]
rlabel metal2 44016 31864 44016 31864 0 cm_inst.page\[1\]
rlabel metal2 32928 34776 32928 34776 0 cm_inst.page\[2\]
rlabel metal2 30744 32200 30744 32200 0 cm_inst.page\[3\]
rlabel metal2 25256 31696 25256 31696 0 cm_inst.page\[4\]
rlabel metal2 22792 32200 22792 32200 0 cm_inst.page\[5\]
rlabel metal2 4312 27888 4312 27888 0 in[0]
rlabel metal2 18872 37352 18872 37352 0 in[1]
rlabel metal3 2478 36344 2478 36344 0 in[2]
rlabel metal2 28112 38696 28112 38696 0 in[3]
rlabel metal2 18984 38668 18984 38668 0 in[4]
rlabel metal3 2534 39704 2534 39704 0 in[5]
rlabel metal2 17416 38976 17416 38976 0 in[6]
rlabel metal2 16632 38668 16632 38668 0 in[7]
rlabel metal2 16072 32872 16072 32872 0 out[0]
rlabel metal3 2086 51800 2086 51800 0 out[10]
rlabel metal3 2702 6776 2702 6776 0 out[11]
rlabel metal3 7854 31640 7854 31640 0 out[1]
rlabel metal3 7910 30968 7910 30968 0 out[2]
rlabel metal3 2198 28952 2198 28952 0 out[3]
rlabel metal2 14000 28728 14000 28728 0 out[4]
rlabel metal3 2478 30296 2478 30296 0 out[5]
rlabel metal3 7742 32984 7742 32984 0 out[6]
rlabel metal2 12600 34216 12600 34216 0 out[7]
rlabel metal3 2478 6104 2478 6104 0 out[8]
rlabel metal2 55272 53984 55272 53984 0 out[9]
rlabel metal3 12432 34440 12432 34440 0 ro_inst.counter\[0\]
rlabel metal3 5376 30520 5376 30520 0 ro_inst.counter\[10\]
rlabel metal3 5432 31864 5432 31864 0 ro_inst.counter\[11\]
rlabel metal2 4536 32872 4536 32872 0 ro_inst.counter\[12\]
rlabel metal3 5376 34552 5376 34552 0 ro_inst.counter\[13\]
rlabel metal2 6216 36288 6216 36288 0 ro_inst.counter\[14\]
rlabel metal2 4536 36960 4536 36960 0 ro_inst.counter\[15\]
rlabel metal2 7280 38024 7280 38024 0 ro_inst.counter\[16\]
rlabel metal2 7672 37352 7672 37352 0 ro_inst.counter\[17\]
rlabel metal2 5432 38696 5432 38696 0 ro_inst.counter\[18\]
rlabel metal2 5768 41216 5768 41216 0 ro_inst.counter\[19\]
rlabel metal3 14224 31752 14224 31752 0 ro_inst.counter\[1\]
rlabel metal3 5600 40600 5600 40600 0 ro_inst.counter\[20\]
rlabel metal2 3528 42168 3528 42168 0 ro_inst.counter\[21\]
rlabel metal2 5320 43232 5320 43232 0 ro_inst.counter\[22\]
rlabel metal3 5600 42840 5600 42840 0 ro_inst.counter\[23\]
rlabel metal2 5768 46928 5768 46928 0 ro_inst.counter\[24\]
rlabel metal2 5768 45248 5768 45248 0 ro_inst.counter\[25\]
rlabel metal2 8904 44968 8904 44968 0 ro_inst.counter\[26\]
rlabel metal2 10360 44352 10360 44352 0 ro_inst.counter\[27\]
rlabel metal3 12264 45080 12264 45080 0 ro_inst.counter\[28\]
rlabel metal3 13720 43848 13720 43848 0 ro_inst.counter\[29\]
rlabel metal2 13944 30296 13944 30296 0 ro_inst.counter\[2\]
rlabel metal2 14056 43232 14056 43232 0 ro_inst.counter\[30\]
rlabel metal2 14224 41832 14224 41832 0 ro_inst.counter\[31\]
rlabel metal3 13216 40600 13216 40600 0 ro_inst.counter\[32\]
rlabel metal2 12824 39200 12824 39200 0 ro_inst.counter\[33\]
rlabel via2 14840 36904 14840 36904 0 ro_inst.counter\[34\]
rlabel metal3 13440 28952 13440 28952 0 ro_inst.counter\[3\]
rlabel metal2 12880 30520 12880 30520 0 ro_inst.counter\[4\]
rlabel metal2 12824 28280 12824 28280 0 ro_inst.counter\[5\]
rlabel metal2 4760 30128 4760 30128 0 ro_inst.counter\[6\]
rlabel metal2 3920 27944 3920 27944 0 ro_inst.counter\[7\]
rlabel metal2 3416 29624 3416 29624 0 ro_inst.counter\[8\]
rlabel metal2 1960 29344 1960 29344 0 ro_inst.counter\[9\]
rlabel metal3 11312 32424 11312 32424 0 ro_inst.counter_n\[0\]
rlabel metal2 2408 30800 2408 30800 0 ro_inst.counter_n\[10\]
rlabel metal3 3808 33096 3808 33096 0 ro_inst.counter_n\[11\]
rlabel metal2 3304 33936 3304 33936 0 ro_inst.counter_n\[12\]
rlabel metal2 2408 34832 2408 34832 0 ro_inst.counter_n\[13\]
rlabel metal2 3584 35784 3584 35784 0 ro_inst.counter_n\[14\]
rlabel metal2 4144 37800 4144 37800 0 ro_inst.counter_n\[15\]
rlabel metal2 5656 37520 5656 37520 0 ro_inst.counter_n\[16\]
rlabel metal2 6272 36792 6272 36792 0 ro_inst.counter_n\[17\]
rlabel metal2 4984 39536 4984 39536 0 ro_inst.counter_n\[18\]
rlabel metal2 4424 41664 4424 41664 0 ro_inst.counter_n\[19\]
rlabel metal2 11368 31808 11368 31808 0 ro_inst.counter_n\[1\]
rlabel metal2 2408 40880 2408 40880 0 ro_inst.counter_n\[20\]
rlabel metal2 2184 43764 2184 43764 0 ro_inst.counter_n\[21\]
rlabel metal2 1904 44856 1904 44856 0 ro_inst.counter_n\[22\]
rlabel metal2 2408 44744 2408 44744 0 ro_inst.counter_n\[23\]
rlabel metal3 4816 46984 4816 46984 0 ro_inst.counter_n\[24\]
rlabel metal2 5656 45528 5656 45528 0 ro_inst.counter_n\[25\]
rlabel metal2 6104 45192 6104 45192 0 ro_inst.counter_n\[26\]
rlabel metal2 10192 44184 10192 44184 0 ro_inst.counter_n\[27\]
rlabel metal2 10248 44912 10248 44912 0 ro_inst.counter_n\[28\]
rlabel metal3 12712 43960 12712 43960 0 ro_inst.counter_n\[29\]
rlabel metal2 11368 29400 11368 29400 0 ro_inst.counter_n\[2\]
rlabel metal3 12488 43176 12488 43176 0 ro_inst.counter_n\[30\]
rlabel metal2 11368 41720 11368 41720 0 ro_inst.counter_n\[31\]
rlabel metal2 10248 40768 10248 40768 0 ro_inst.counter_n\[32\]
rlabel metal2 12712 39480 12712 39480 0 ro_inst.counter_n\[33\]
rlabel metal2 12264 38248 12264 38248 0 ro_inst.counter_n\[34\]
rlabel metal3 10024 30072 10024 30072 0 ro_inst.counter_n\[3\]
rlabel metal2 9912 28560 9912 28560 0 ro_inst.counter_n\[4\]
rlabel metal2 7896 29568 7896 29568 0 ro_inst.counter_n\[5\]
rlabel metal2 7336 29792 7336 29792 0 ro_inst.counter_n\[6\]
rlabel metal2 5656 28896 5656 28896 0 ro_inst.counter_n\[7\]
rlabel metal2 5096 29064 5096 29064 0 ro_inst.counter_n\[8\]
rlabel metal3 2856 30072 2856 30072 0 ro_inst.counter_n\[9\]
rlabel metal2 13720 35168 13720 35168 0 ro_inst.enable
rlabel metal3 11032 34664 11032 34664 0 ro_inst.ring\[0\]
rlabel metal2 13608 35784 13608 35784 0 ro_inst.ring\[1\]
rlabel metal2 9800 35616 9800 35616 0 ro_inst.ring\[2\]
rlabel metal2 10472 34944 10472 34944 0 ro_inst.running
rlabel metal3 11536 34104 11536 34104 0 ro_inst.saved_signal
rlabel metal2 10920 33880 10920 33880 0 ro_inst.signal
rlabel metal2 10360 34160 10360 34160 0 ro_inst.slow_clk_n
rlabel metal2 17808 31528 17808 31528 0 ro_sel\[0\]
rlabel metal2 18592 34776 18592 34776 0 ro_sel\[1\]
rlabel metal2 17864 36064 17864 36064 0 ro_sel\[2\]
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
