magic
tech gf180mcuD
magscale 1 10
timestamp 1702448218
<< metal1 >>
rect 1344 36314 38800 36348
rect 1344 36262 10538 36314
rect 10590 36262 10642 36314
rect 10694 36262 10746 36314
rect 10798 36262 19862 36314
rect 19914 36262 19966 36314
rect 20018 36262 20070 36314
rect 20122 36262 29186 36314
rect 29238 36262 29290 36314
rect 29342 36262 29394 36314
rect 29446 36262 38510 36314
rect 38562 36262 38614 36314
rect 38666 36262 38718 36314
rect 38770 36262 38800 36314
rect 1344 36228 38800 36262
rect 1344 35306 38640 35340
rect 1344 35254 5876 35306
rect 5928 35254 5980 35306
rect 6032 35254 6084 35306
rect 6136 35254 15200 35306
rect 15252 35254 15304 35306
rect 15356 35254 15408 35306
rect 15460 35254 24524 35306
rect 24576 35254 24628 35306
rect 24680 35254 24732 35306
rect 24784 35254 33848 35306
rect 33900 35254 33952 35306
rect 34004 35254 34056 35306
rect 34108 35254 38640 35306
rect 1344 35220 38640 35254
rect 1344 34298 38800 34332
rect 1344 34246 10538 34298
rect 10590 34246 10642 34298
rect 10694 34246 10746 34298
rect 10798 34246 19862 34298
rect 19914 34246 19966 34298
rect 20018 34246 20070 34298
rect 20122 34246 29186 34298
rect 29238 34246 29290 34298
rect 29342 34246 29394 34298
rect 29446 34246 38510 34298
rect 38562 34246 38614 34298
rect 38666 34246 38718 34298
rect 38770 34246 38800 34298
rect 1344 34212 38800 34246
rect 1344 33290 38640 33324
rect 1344 33238 5876 33290
rect 5928 33238 5980 33290
rect 6032 33238 6084 33290
rect 6136 33238 15200 33290
rect 15252 33238 15304 33290
rect 15356 33238 15408 33290
rect 15460 33238 24524 33290
rect 24576 33238 24628 33290
rect 24680 33238 24732 33290
rect 24784 33238 33848 33290
rect 33900 33238 33952 33290
rect 34004 33238 34056 33290
rect 34108 33238 38640 33290
rect 1344 33204 38640 33238
rect 1344 32282 38800 32316
rect 1344 32230 10538 32282
rect 10590 32230 10642 32282
rect 10694 32230 10746 32282
rect 10798 32230 19862 32282
rect 19914 32230 19966 32282
rect 20018 32230 20070 32282
rect 20122 32230 29186 32282
rect 29238 32230 29290 32282
rect 29342 32230 29394 32282
rect 29446 32230 38510 32282
rect 38562 32230 38614 32282
rect 38666 32230 38718 32282
rect 38770 32230 38800 32282
rect 1344 32196 38800 32230
rect 15474 32062 15486 32114
rect 15538 32062 15550 32114
rect 14926 31890 14978 31902
rect 14926 31826 14978 31838
rect 15150 31890 15202 31902
rect 15150 31826 15202 31838
rect 1344 31274 38640 31308
rect 1344 31222 5876 31274
rect 5928 31222 5980 31274
rect 6032 31222 6084 31274
rect 6136 31222 15200 31274
rect 15252 31222 15304 31274
rect 15356 31222 15408 31274
rect 15460 31222 24524 31274
rect 24576 31222 24628 31274
rect 24680 31222 24732 31274
rect 24784 31222 33848 31274
rect 33900 31222 33952 31274
rect 34004 31222 34056 31274
rect 34108 31222 38640 31274
rect 1344 31188 38640 31222
rect 1344 30266 38800 30300
rect 1344 30214 10538 30266
rect 10590 30214 10642 30266
rect 10694 30214 10746 30266
rect 10798 30214 19862 30266
rect 19914 30214 19966 30266
rect 20018 30214 20070 30266
rect 20122 30214 29186 30266
rect 29238 30214 29290 30266
rect 29342 30214 29394 30266
rect 29446 30214 38510 30266
rect 38562 30214 38614 30266
rect 38666 30214 38718 30266
rect 38770 30214 38800 30266
rect 1344 30180 38800 30214
rect 1344 29258 38640 29292
rect 1344 29206 5876 29258
rect 5928 29206 5980 29258
rect 6032 29206 6084 29258
rect 6136 29206 15200 29258
rect 15252 29206 15304 29258
rect 15356 29206 15408 29258
rect 15460 29206 24524 29258
rect 24576 29206 24628 29258
rect 24680 29206 24732 29258
rect 24784 29206 33848 29258
rect 33900 29206 33952 29258
rect 34004 29206 34056 29258
rect 34108 29206 38640 29258
rect 1344 29172 38640 29206
rect 1344 28250 38800 28284
rect 1344 28198 10538 28250
rect 10590 28198 10642 28250
rect 10694 28198 10746 28250
rect 10798 28198 19862 28250
rect 19914 28198 19966 28250
rect 20018 28198 20070 28250
rect 20122 28198 29186 28250
rect 29238 28198 29290 28250
rect 29342 28198 29394 28250
rect 29446 28198 38510 28250
rect 38562 28198 38614 28250
rect 38666 28198 38718 28250
rect 38770 28198 38800 28250
rect 1344 28164 38800 28198
rect 1344 27242 38640 27276
rect 1344 27190 5876 27242
rect 5928 27190 5980 27242
rect 6032 27190 6084 27242
rect 6136 27190 15200 27242
rect 15252 27190 15304 27242
rect 15356 27190 15408 27242
rect 15460 27190 24524 27242
rect 24576 27190 24628 27242
rect 24680 27190 24732 27242
rect 24784 27190 33848 27242
rect 33900 27190 33952 27242
rect 34004 27190 34056 27242
rect 34108 27190 38640 27242
rect 1344 27156 38640 27190
rect 1344 26234 38800 26268
rect 1344 26182 10538 26234
rect 10590 26182 10642 26234
rect 10694 26182 10746 26234
rect 10798 26182 19862 26234
rect 19914 26182 19966 26234
rect 20018 26182 20070 26234
rect 20122 26182 29186 26234
rect 29238 26182 29290 26234
rect 29342 26182 29394 26234
rect 29446 26182 38510 26234
rect 38562 26182 38614 26234
rect 38666 26182 38718 26234
rect 38770 26182 38800 26234
rect 1344 26148 38800 26182
rect 1344 25226 38640 25260
rect 1344 25174 5876 25226
rect 5928 25174 5980 25226
rect 6032 25174 6084 25226
rect 6136 25174 15200 25226
rect 15252 25174 15304 25226
rect 15356 25174 15408 25226
rect 15460 25174 24524 25226
rect 24576 25174 24628 25226
rect 24680 25174 24732 25226
rect 24784 25174 33848 25226
rect 33900 25174 33952 25226
rect 34004 25174 34056 25226
rect 34108 25174 38640 25226
rect 1344 25140 38640 25174
rect 1344 24218 38800 24252
rect 1344 24166 10538 24218
rect 10590 24166 10642 24218
rect 10694 24166 10746 24218
rect 10798 24166 19862 24218
rect 19914 24166 19966 24218
rect 20018 24166 20070 24218
rect 20122 24166 29186 24218
rect 29238 24166 29290 24218
rect 29342 24166 29394 24218
rect 29446 24166 38510 24218
rect 38562 24166 38614 24218
rect 38666 24166 38718 24218
rect 38770 24166 38800 24218
rect 1344 24132 38800 24166
rect 1344 23210 38640 23244
rect 1344 23158 5876 23210
rect 5928 23158 5980 23210
rect 6032 23158 6084 23210
rect 6136 23158 15200 23210
rect 15252 23158 15304 23210
rect 15356 23158 15408 23210
rect 15460 23158 24524 23210
rect 24576 23158 24628 23210
rect 24680 23158 24732 23210
rect 24784 23158 33848 23210
rect 33900 23158 33952 23210
rect 34004 23158 34056 23210
rect 34108 23158 38640 23210
rect 1344 23124 38640 23158
rect 1344 22202 38800 22236
rect 1344 22150 10538 22202
rect 10590 22150 10642 22202
rect 10694 22150 10746 22202
rect 10798 22150 19862 22202
rect 19914 22150 19966 22202
rect 20018 22150 20070 22202
rect 20122 22150 29186 22202
rect 29238 22150 29290 22202
rect 29342 22150 29394 22202
rect 29446 22150 38510 22202
rect 38562 22150 38614 22202
rect 38666 22150 38718 22202
rect 38770 22150 38800 22202
rect 1344 22116 38800 22150
rect 1344 21194 38640 21228
rect 1344 21142 5876 21194
rect 5928 21142 5980 21194
rect 6032 21142 6084 21194
rect 6136 21142 15200 21194
rect 15252 21142 15304 21194
rect 15356 21142 15408 21194
rect 15460 21142 24524 21194
rect 24576 21142 24628 21194
rect 24680 21142 24732 21194
rect 24784 21142 33848 21194
rect 33900 21142 33952 21194
rect 34004 21142 34056 21194
rect 34108 21142 38640 21194
rect 1344 21108 38640 21142
rect 19282 20974 19294 21026
rect 19346 20974 19358 21026
rect 31054 20914 31106 20926
rect 18050 20862 18062 20914
rect 18114 20862 18126 20914
rect 31054 20850 31106 20862
rect 13694 20802 13746 20814
rect 13694 20738 13746 20750
rect 13918 20690 13970 20702
rect 13918 20626 13970 20638
rect 14926 20690 14978 20702
rect 14926 20626 14978 20638
rect 18398 20690 18450 20702
rect 18398 20626 18450 20638
rect 18846 20690 18898 20702
rect 21858 20638 21870 20690
rect 21922 20638 21934 20690
rect 22082 20638 22094 20690
rect 22146 20638 22158 20690
rect 22306 20638 22318 20690
rect 22370 20638 22382 20690
rect 18846 20626 18898 20638
rect 19406 20578 19458 20590
rect 19406 20514 19458 20526
rect 20414 20578 20466 20590
rect 20414 20514 20466 20526
rect 23438 20578 23490 20590
rect 23438 20514 23490 20526
rect 24334 20578 24386 20590
rect 24334 20514 24386 20526
rect 26126 20578 26178 20590
rect 26126 20514 26178 20526
rect 29150 20578 29202 20590
rect 29150 20514 29202 20526
rect 30718 20578 30770 20590
rect 30718 20514 30770 20526
rect 12462 20466 12514 20478
rect 12462 20402 12514 20414
rect 12910 20466 12962 20478
rect 12910 20402 12962 20414
rect 13470 20466 13522 20478
rect 13470 20402 13522 20414
rect 17614 20466 17666 20478
rect 17614 20402 17666 20414
rect 22878 20466 22930 20478
rect 22878 20402 22930 20414
rect 30046 20466 30098 20478
rect 30046 20402 30098 20414
rect 20738 20302 20750 20354
rect 20802 20302 20814 20354
rect 23762 20302 23774 20354
rect 23826 20302 23838 20354
rect 26450 20302 26462 20354
rect 26514 20302 26526 20354
rect 29474 20302 29486 20354
rect 29538 20302 29550 20354
rect 1344 20186 38800 20220
rect 1344 20134 10538 20186
rect 10590 20134 10642 20186
rect 10694 20134 10746 20186
rect 10798 20134 19862 20186
rect 19914 20134 19966 20186
rect 20018 20134 20070 20186
rect 20122 20134 29186 20186
rect 29238 20134 29290 20186
rect 29342 20134 29394 20186
rect 29446 20134 38510 20186
rect 38562 20134 38614 20186
rect 38666 20134 38718 20186
rect 38770 20134 38800 20186
rect 1344 20100 38800 20134
rect 17614 19906 17666 19918
rect 16706 19854 16718 19906
rect 16770 19854 16782 19906
rect 17614 19842 17666 19854
rect 20078 19906 20130 19918
rect 20078 19842 20130 19854
rect 25342 19906 25394 19918
rect 31950 19906 32002 19918
rect 25342 19842 25394 19854
rect 26898 19829 26910 19881
rect 26962 19829 26974 19881
rect 31950 19842 32002 19854
rect 12910 19794 12962 19806
rect 22654 19794 22706 19806
rect 12674 19742 12686 19794
rect 12738 19742 12750 19794
rect 16482 19742 16494 19794
rect 16546 19742 16558 19794
rect 12910 19730 12962 19742
rect 22654 19730 22706 19742
rect 30718 19794 30770 19806
rect 30718 19730 30770 19742
rect 14254 19682 14306 19694
rect 21534 19682 21586 19694
rect 13794 19630 13806 19682
rect 13858 19630 13870 19682
rect 14690 19630 14702 19682
rect 14754 19630 14766 19682
rect 14914 19630 14926 19682
rect 14978 19630 14990 19682
rect 18274 19630 18286 19682
rect 18338 19630 18350 19682
rect 19506 19630 19518 19682
rect 19570 19630 19582 19682
rect 14254 19618 14306 19630
rect 21534 19618 21586 19630
rect 23662 19682 23714 19694
rect 24210 19630 24222 19682
rect 24274 19630 24286 19682
rect 24658 19630 24670 19682
rect 24722 19630 24734 19682
rect 28018 19630 28030 19682
rect 28082 19630 28094 19682
rect 29362 19630 29374 19682
rect 29426 19630 29438 19682
rect 23662 19618 23714 19630
rect 22878 19570 22930 19582
rect 18162 19518 18174 19570
rect 18226 19518 18238 19570
rect 20850 19518 20862 19570
rect 20914 19518 20926 19570
rect 22878 19506 22930 19518
rect 25790 19570 25842 19582
rect 25790 19506 25842 19518
rect 26350 19570 26402 19582
rect 30942 19570 30994 19582
rect 28466 19518 28478 19570
rect 28530 19518 28542 19570
rect 28914 19518 28926 19570
rect 28978 19518 28990 19570
rect 26350 19506 26402 19518
rect 30942 19506 30994 19518
rect 31502 19570 31554 19582
rect 31502 19506 31554 19518
rect 1344 19178 38640 19212
rect 1344 19126 5876 19178
rect 5928 19126 5980 19178
rect 6032 19126 6084 19178
rect 6136 19126 15200 19178
rect 15252 19126 15304 19178
rect 15356 19126 15408 19178
rect 15460 19126 24524 19178
rect 24576 19126 24628 19178
rect 24680 19126 24732 19178
rect 24784 19126 33848 19178
rect 33900 19126 33952 19178
rect 34004 19126 34056 19178
rect 34108 19126 38640 19178
rect 1344 19092 38640 19126
rect 12674 18846 12686 18898
rect 12738 18846 12750 18898
rect 13806 18786 13858 18798
rect 13806 18722 13858 18734
rect 15934 18786 15986 18798
rect 15934 18722 15986 18734
rect 16270 18786 16322 18798
rect 16270 18722 16322 18734
rect 16830 18786 16882 18798
rect 16830 18722 16882 18734
rect 18174 18786 18226 18798
rect 18174 18722 18226 18734
rect 23438 18786 23490 18798
rect 26014 18786 26066 18798
rect 25554 18734 25566 18786
rect 25618 18734 25630 18786
rect 23438 18722 23490 18734
rect 26014 18722 26066 18734
rect 27358 18786 27410 18798
rect 29362 18734 29374 18786
rect 29426 18734 29438 18786
rect 27358 18722 27410 18734
rect 11566 18674 11618 18686
rect 11566 18610 11618 18622
rect 12014 18674 12066 18686
rect 12014 18610 12066 18622
rect 12126 18674 12178 18686
rect 16606 18674 16658 18686
rect 13906 18622 13918 18674
rect 13970 18622 13982 18674
rect 14130 18622 14142 18674
rect 14194 18622 14206 18674
rect 12126 18610 12178 18622
rect 16606 18610 16658 18622
rect 17054 18674 17106 18686
rect 30606 18674 30658 18686
rect 25106 18622 25118 18674
rect 25170 18622 25182 18674
rect 26898 18622 26910 18674
rect 26962 18622 26974 18674
rect 27234 18622 27246 18674
rect 27298 18622 27310 18674
rect 29698 18622 29710 18674
rect 29762 18622 29774 18674
rect 17054 18610 17106 18622
rect 30606 18610 30658 18622
rect 11118 18562 11170 18574
rect 11118 18498 11170 18510
rect 23662 18562 23714 18574
rect 23662 18498 23714 18510
rect 27918 18562 27970 18574
rect 27918 18498 27970 18510
rect 28590 18562 28642 18574
rect 28590 18498 28642 18510
rect 30034 18398 30046 18450
rect 30098 18398 30110 18450
rect 1344 18170 38800 18204
rect 1344 18118 10538 18170
rect 10590 18118 10642 18170
rect 10694 18118 10746 18170
rect 10798 18118 19862 18170
rect 19914 18118 19966 18170
rect 20018 18118 20070 18170
rect 20122 18118 29186 18170
rect 29238 18118 29290 18170
rect 29342 18118 29394 18170
rect 29446 18118 38510 18170
rect 38562 18118 38614 18170
rect 38666 18118 38718 18170
rect 38770 18118 38800 18170
rect 1344 18084 38800 18118
rect 13470 17890 13522 17902
rect 13470 17826 13522 17838
rect 13918 17890 13970 17902
rect 13918 17826 13970 17838
rect 26014 17554 26066 17566
rect 26014 17490 26066 17502
rect 1344 17162 38640 17196
rect 1344 17110 5876 17162
rect 5928 17110 5980 17162
rect 6032 17110 6084 17162
rect 6136 17110 15200 17162
rect 15252 17110 15304 17162
rect 15356 17110 15408 17162
rect 15460 17110 24524 17162
rect 24576 17110 24628 17162
rect 24680 17110 24732 17162
rect 24784 17110 33848 17162
rect 33900 17110 33952 17162
rect 34004 17110 34056 17162
rect 34108 17110 38640 17162
rect 1344 17076 38640 17110
rect 1344 16154 38800 16188
rect 1344 16102 10538 16154
rect 10590 16102 10642 16154
rect 10694 16102 10746 16154
rect 10798 16102 19862 16154
rect 19914 16102 19966 16154
rect 20018 16102 20070 16154
rect 20122 16102 29186 16154
rect 29238 16102 29290 16154
rect 29342 16102 29394 16154
rect 29446 16102 38510 16154
rect 38562 16102 38614 16154
rect 38666 16102 38718 16154
rect 38770 16102 38800 16154
rect 1344 16068 38800 16102
rect 1344 15146 38640 15180
rect 1344 15094 5876 15146
rect 5928 15094 5980 15146
rect 6032 15094 6084 15146
rect 6136 15094 15200 15146
rect 15252 15094 15304 15146
rect 15356 15094 15408 15146
rect 15460 15094 24524 15146
rect 24576 15094 24628 15146
rect 24680 15094 24732 15146
rect 24784 15094 33848 15146
rect 33900 15094 33952 15146
rect 34004 15094 34056 15146
rect 34108 15094 38640 15146
rect 1344 15060 38640 15094
rect 1344 14138 38800 14172
rect 1344 14086 10538 14138
rect 10590 14086 10642 14138
rect 10694 14086 10746 14138
rect 10798 14086 19862 14138
rect 19914 14086 19966 14138
rect 20018 14086 20070 14138
rect 20122 14086 29186 14138
rect 29238 14086 29290 14138
rect 29342 14086 29394 14138
rect 29446 14086 38510 14138
rect 38562 14086 38614 14138
rect 38666 14086 38718 14138
rect 38770 14086 38800 14138
rect 1344 14052 38800 14086
rect 1344 13130 38640 13164
rect 1344 13078 5876 13130
rect 5928 13078 5980 13130
rect 6032 13078 6084 13130
rect 6136 13078 15200 13130
rect 15252 13078 15304 13130
rect 15356 13078 15408 13130
rect 15460 13078 24524 13130
rect 24576 13078 24628 13130
rect 24680 13078 24732 13130
rect 24784 13078 33848 13130
rect 33900 13078 33952 13130
rect 34004 13078 34056 13130
rect 34108 13078 38640 13130
rect 1344 13044 38640 13078
rect 1344 12122 38800 12156
rect 1344 12070 10538 12122
rect 10590 12070 10642 12122
rect 10694 12070 10746 12122
rect 10798 12070 19862 12122
rect 19914 12070 19966 12122
rect 20018 12070 20070 12122
rect 20122 12070 29186 12122
rect 29238 12070 29290 12122
rect 29342 12070 29394 12122
rect 29446 12070 38510 12122
rect 38562 12070 38614 12122
rect 38666 12070 38718 12122
rect 38770 12070 38800 12122
rect 1344 12036 38800 12070
rect 1344 11114 38640 11148
rect 1344 11062 5876 11114
rect 5928 11062 5980 11114
rect 6032 11062 6084 11114
rect 6136 11062 15200 11114
rect 15252 11062 15304 11114
rect 15356 11062 15408 11114
rect 15460 11062 24524 11114
rect 24576 11062 24628 11114
rect 24680 11062 24732 11114
rect 24784 11062 33848 11114
rect 33900 11062 33952 11114
rect 34004 11062 34056 11114
rect 34108 11062 38640 11114
rect 1344 11028 38640 11062
rect 1344 10106 38800 10140
rect 1344 10054 10538 10106
rect 10590 10054 10642 10106
rect 10694 10054 10746 10106
rect 10798 10054 19862 10106
rect 19914 10054 19966 10106
rect 20018 10054 20070 10106
rect 20122 10054 29186 10106
rect 29238 10054 29290 10106
rect 29342 10054 29394 10106
rect 29446 10054 38510 10106
rect 38562 10054 38614 10106
rect 38666 10054 38718 10106
rect 38770 10054 38800 10106
rect 1344 10020 38800 10054
rect 1344 9098 38640 9132
rect 1344 9046 5876 9098
rect 5928 9046 5980 9098
rect 6032 9046 6084 9098
rect 6136 9046 15200 9098
rect 15252 9046 15304 9098
rect 15356 9046 15408 9098
rect 15460 9046 24524 9098
rect 24576 9046 24628 9098
rect 24680 9046 24732 9098
rect 24784 9046 33848 9098
rect 33900 9046 33952 9098
rect 34004 9046 34056 9098
rect 34108 9046 38640 9098
rect 1344 9012 38640 9046
rect 1344 8090 38800 8124
rect 1344 8038 10538 8090
rect 10590 8038 10642 8090
rect 10694 8038 10746 8090
rect 10798 8038 19862 8090
rect 19914 8038 19966 8090
rect 20018 8038 20070 8090
rect 20122 8038 29186 8090
rect 29238 8038 29290 8090
rect 29342 8038 29394 8090
rect 29446 8038 38510 8090
rect 38562 8038 38614 8090
rect 38666 8038 38718 8090
rect 38770 8038 38800 8090
rect 1344 8004 38800 8038
rect 1344 7082 38640 7116
rect 1344 7030 5876 7082
rect 5928 7030 5980 7082
rect 6032 7030 6084 7082
rect 6136 7030 15200 7082
rect 15252 7030 15304 7082
rect 15356 7030 15408 7082
rect 15460 7030 24524 7082
rect 24576 7030 24628 7082
rect 24680 7030 24732 7082
rect 24784 7030 33848 7082
rect 33900 7030 33952 7082
rect 34004 7030 34056 7082
rect 34108 7030 38640 7082
rect 1344 6996 38640 7030
rect 1344 6074 38800 6108
rect 1344 6022 10538 6074
rect 10590 6022 10642 6074
rect 10694 6022 10746 6074
rect 10798 6022 19862 6074
rect 19914 6022 19966 6074
rect 20018 6022 20070 6074
rect 20122 6022 29186 6074
rect 29238 6022 29290 6074
rect 29342 6022 29394 6074
rect 29446 6022 38510 6074
rect 38562 6022 38614 6074
rect 38666 6022 38718 6074
rect 38770 6022 38800 6074
rect 1344 5988 38800 6022
rect 1344 5066 38640 5100
rect 1344 5014 5876 5066
rect 5928 5014 5980 5066
rect 6032 5014 6084 5066
rect 6136 5014 15200 5066
rect 15252 5014 15304 5066
rect 15356 5014 15408 5066
rect 15460 5014 24524 5066
rect 24576 5014 24628 5066
rect 24680 5014 24732 5066
rect 24784 5014 33848 5066
rect 33900 5014 33952 5066
rect 34004 5014 34056 5066
rect 34108 5014 38640 5066
rect 1344 4980 38640 5014
rect 1344 4058 38800 4092
rect 1344 4006 10538 4058
rect 10590 4006 10642 4058
rect 10694 4006 10746 4058
rect 10798 4006 19862 4058
rect 19914 4006 19966 4058
rect 20018 4006 20070 4058
rect 20122 4006 29186 4058
rect 29238 4006 29290 4058
rect 29342 4006 29394 4058
rect 29446 4006 38510 4058
rect 38562 4006 38614 4058
rect 38666 4006 38718 4058
rect 38770 4006 38800 4058
rect 1344 3972 38800 4006
<< via1 >>
rect 10538 36262 10590 36314
rect 10642 36262 10694 36314
rect 10746 36262 10798 36314
rect 19862 36262 19914 36314
rect 19966 36262 20018 36314
rect 20070 36262 20122 36314
rect 29186 36262 29238 36314
rect 29290 36262 29342 36314
rect 29394 36262 29446 36314
rect 38510 36262 38562 36314
rect 38614 36262 38666 36314
rect 38718 36262 38770 36314
rect 5876 35254 5928 35306
rect 5980 35254 6032 35306
rect 6084 35254 6136 35306
rect 15200 35254 15252 35306
rect 15304 35254 15356 35306
rect 15408 35254 15460 35306
rect 24524 35254 24576 35306
rect 24628 35254 24680 35306
rect 24732 35254 24784 35306
rect 33848 35254 33900 35306
rect 33952 35254 34004 35306
rect 34056 35254 34108 35306
rect 10538 34246 10590 34298
rect 10642 34246 10694 34298
rect 10746 34246 10798 34298
rect 19862 34246 19914 34298
rect 19966 34246 20018 34298
rect 20070 34246 20122 34298
rect 29186 34246 29238 34298
rect 29290 34246 29342 34298
rect 29394 34246 29446 34298
rect 38510 34246 38562 34298
rect 38614 34246 38666 34298
rect 38718 34246 38770 34298
rect 5876 33238 5928 33290
rect 5980 33238 6032 33290
rect 6084 33238 6136 33290
rect 15200 33238 15252 33290
rect 15304 33238 15356 33290
rect 15408 33238 15460 33290
rect 24524 33238 24576 33290
rect 24628 33238 24680 33290
rect 24732 33238 24784 33290
rect 33848 33238 33900 33290
rect 33952 33238 34004 33290
rect 34056 33238 34108 33290
rect 10538 32230 10590 32282
rect 10642 32230 10694 32282
rect 10746 32230 10798 32282
rect 19862 32230 19914 32282
rect 19966 32230 20018 32282
rect 20070 32230 20122 32282
rect 29186 32230 29238 32282
rect 29290 32230 29342 32282
rect 29394 32230 29446 32282
rect 38510 32230 38562 32282
rect 38614 32230 38666 32282
rect 38718 32230 38770 32282
rect 15486 32062 15538 32114
rect 14926 31838 14978 31890
rect 15150 31838 15202 31890
rect 5876 31222 5928 31274
rect 5980 31222 6032 31274
rect 6084 31222 6136 31274
rect 15200 31222 15252 31274
rect 15304 31222 15356 31274
rect 15408 31222 15460 31274
rect 24524 31222 24576 31274
rect 24628 31222 24680 31274
rect 24732 31222 24784 31274
rect 33848 31222 33900 31274
rect 33952 31222 34004 31274
rect 34056 31222 34108 31274
rect 10538 30214 10590 30266
rect 10642 30214 10694 30266
rect 10746 30214 10798 30266
rect 19862 30214 19914 30266
rect 19966 30214 20018 30266
rect 20070 30214 20122 30266
rect 29186 30214 29238 30266
rect 29290 30214 29342 30266
rect 29394 30214 29446 30266
rect 38510 30214 38562 30266
rect 38614 30214 38666 30266
rect 38718 30214 38770 30266
rect 5876 29206 5928 29258
rect 5980 29206 6032 29258
rect 6084 29206 6136 29258
rect 15200 29206 15252 29258
rect 15304 29206 15356 29258
rect 15408 29206 15460 29258
rect 24524 29206 24576 29258
rect 24628 29206 24680 29258
rect 24732 29206 24784 29258
rect 33848 29206 33900 29258
rect 33952 29206 34004 29258
rect 34056 29206 34108 29258
rect 10538 28198 10590 28250
rect 10642 28198 10694 28250
rect 10746 28198 10798 28250
rect 19862 28198 19914 28250
rect 19966 28198 20018 28250
rect 20070 28198 20122 28250
rect 29186 28198 29238 28250
rect 29290 28198 29342 28250
rect 29394 28198 29446 28250
rect 38510 28198 38562 28250
rect 38614 28198 38666 28250
rect 38718 28198 38770 28250
rect 5876 27190 5928 27242
rect 5980 27190 6032 27242
rect 6084 27190 6136 27242
rect 15200 27190 15252 27242
rect 15304 27190 15356 27242
rect 15408 27190 15460 27242
rect 24524 27190 24576 27242
rect 24628 27190 24680 27242
rect 24732 27190 24784 27242
rect 33848 27190 33900 27242
rect 33952 27190 34004 27242
rect 34056 27190 34108 27242
rect 10538 26182 10590 26234
rect 10642 26182 10694 26234
rect 10746 26182 10798 26234
rect 19862 26182 19914 26234
rect 19966 26182 20018 26234
rect 20070 26182 20122 26234
rect 29186 26182 29238 26234
rect 29290 26182 29342 26234
rect 29394 26182 29446 26234
rect 38510 26182 38562 26234
rect 38614 26182 38666 26234
rect 38718 26182 38770 26234
rect 5876 25174 5928 25226
rect 5980 25174 6032 25226
rect 6084 25174 6136 25226
rect 15200 25174 15252 25226
rect 15304 25174 15356 25226
rect 15408 25174 15460 25226
rect 24524 25174 24576 25226
rect 24628 25174 24680 25226
rect 24732 25174 24784 25226
rect 33848 25174 33900 25226
rect 33952 25174 34004 25226
rect 34056 25174 34108 25226
rect 10538 24166 10590 24218
rect 10642 24166 10694 24218
rect 10746 24166 10798 24218
rect 19862 24166 19914 24218
rect 19966 24166 20018 24218
rect 20070 24166 20122 24218
rect 29186 24166 29238 24218
rect 29290 24166 29342 24218
rect 29394 24166 29446 24218
rect 38510 24166 38562 24218
rect 38614 24166 38666 24218
rect 38718 24166 38770 24218
rect 5876 23158 5928 23210
rect 5980 23158 6032 23210
rect 6084 23158 6136 23210
rect 15200 23158 15252 23210
rect 15304 23158 15356 23210
rect 15408 23158 15460 23210
rect 24524 23158 24576 23210
rect 24628 23158 24680 23210
rect 24732 23158 24784 23210
rect 33848 23158 33900 23210
rect 33952 23158 34004 23210
rect 34056 23158 34108 23210
rect 10538 22150 10590 22202
rect 10642 22150 10694 22202
rect 10746 22150 10798 22202
rect 19862 22150 19914 22202
rect 19966 22150 20018 22202
rect 20070 22150 20122 22202
rect 29186 22150 29238 22202
rect 29290 22150 29342 22202
rect 29394 22150 29446 22202
rect 38510 22150 38562 22202
rect 38614 22150 38666 22202
rect 38718 22150 38770 22202
rect 5876 21142 5928 21194
rect 5980 21142 6032 21194
rect 6084 21142 6136 21194
rect 15200 21142 15252 21194
rect 15304 21142 15356 21194
rect 15408 21142 15460 21194
rect 24524 21142 24576 21194
rect 24628 21142 24680 21194
rect 24732 21142 24784 21194
rect 33848 21142 33900 21194
rect 33952 21142 34004 21194
rect 34056 21142 34108 21194
rect 19294 20974 19346 21026
rect 18062 20862 18114 20914
rect 31054 20862 31106 20914
rect 13694 20750 13746 20802
rect 13918 20638 13970 20690
rect 14926 20638 14978 20690
rect 18398 20638 18450 20690
rect 18846 20638 18898 20690
rect 21870 20638 21922 20690
rect 22094 20638 22146 20690
rect 22318 20638 22370 20690
rect 19406 20526 19458 20578
rect 20414 20526 20466 20578
rect 23438 20526 23490 20578
rect 24334 20526 24386 20578
rect 26126 20526 26178 20578
rect 29150 20526 29202 20578
rect 30718 20526 30770 20578
rect 12462 20414 12514 20466
rect 12910 20414 12962 20466
rect 13470 20414 13522 20466
rect 17614 20414 17666 20466
rect 22878 20414 22930 20466
rect 30046 20414 30098 20466
rect 20750 20302 20802 20354
rect 23774 20302 23826 20354
rect 26462 20302 26514 20354
rect 29486 20302 29538 20354
rect 10538 20134 10590 20186
rect 10642 20134 10694 20186
rect 10746 20134 10798 20186
rect 19862 20134 19914 20186
rect 19966 20134 20018 20186
rect 20070 20134 20122 20186
rect 29186 20134 29238 20186
rect 29290 20134 29342 20186
rect 29394 20134 29446 20186
rect 38510 20134 38562 20186
rect 38614 20134 38666 20186
rect 38718 20134 38770 20186
rect 16718 19854 16770 19906
rect 17614 19854 17666 19906
rect 20078 19854 20130 19906
rect 25342 19854 25394 19906
rect 26910 19829 26962 19881
rect 31950 19854 32002 19906
rect 12686 19742 12738 19794
rect 12910 19742 12962 19794
rect 16494 19742 16546 19794
rect 22654 19742 22706 19794
rect 30718 19742 30770 19794
rect 13806 19630 13858 19682
rect 14254 19630 14306 19682
rect 14702 19630 14754 19682
rect 14926 19630 14978 19682
rect 18286 19630 18338 19682
rect 19518 19630 19570 19682
rect 21534 19630 21586 19682
rect 23662 19630 23714 19682
rect 24222 19630 24274 19682
rect 24670 19630 24722 19682
rect 28030 19630 28082 19682
rect 29374 19630 29426 19682
rect 18174 19518 18226 19570
rect 20862 19518 20914 19570
rect 22878 19518 22930 19570
rect 25790 19518 25842 19570
rect 26350 19518 26402 19570
rect 28478 19518 28530 19570
rect 28926 19518 28978 19570
rect 30942 19518 30994 19570
rect 31502 19518 31554 19570
rect 5876 19126 5928 19178
rect 5980 19126 6032 19178
rect 6084 19126 6136 19178
rect 15200 19126 15252 19178
rect 15304 19126 15356 19178
rect 15408 19126 15460 19178
rect 24524 19126 24576 19178
rect 24628 19126 24680 19178
rect 24732 19126 24784 19178
rect 33848 19126 33900 19178
rect 33952 19126 34004 19178
rect 34056 19126 34108 19178
rect 12686 18846 12738 18898
rect 13806 18734 13858 18786
rect 15934 18734 15986 18786
rect 16270 18734 16322 18786
rect 16830 18734 16882 18786
rect 18174 18734 18226 18786
rect 23438 18734 23490 18786
rect 25566 18734 25618 18786
rect 26014 18734 26066 18786
rect 27358 18734 27410 18786
rect 29374 18734 29426 18786
rect 11566 18622 11618 18674
rect 12014 18622 12066 18674
rect 12126 18622 12178 18674
rect 13918 18622 13970 18674
rect 14142 18622 14194 18674
rect 16606 18622 16658 18674
rect 17054 18622 17106 18674
rect 25118 18622 25170 18674
rect 26910 18622 26962 18674
rect 27246 18622 27298 18674
rect 29710 18622 29762 18674
rect 30606 18622 30658 18674
rect 11118 18510 11170 18562
rect 23662 18510 23714 18562
rect 27918 18510 27970 18562
rect 28590 18510 28642 18562
rect 30046 18398 30098 18450
rect 10538 18118 10590 18170
rect 10642 18118 10694 18170
rect 10746 18118 10798 18170
rect 19862 18118 19914 18170
rect 19966 18118 20018 18170
rect 20070 18118 20122 18170
rect 29186 18118 29238 18170
rect 29290 18118 29342 18170
rect 29394 18118 29446 18170
rect 38510 18118 38562 18170
rect 38614 18118 38666 18170
rect 38718 18118 38770 18170
rect 13470 17838 13522 17890
rect 13918 17838 13970 17890
rect 26014 17502 26066 17554
rect 5876 17110 5928 17162
rect 5980 17110 6032 17162
rect 6084 17110 6136 17162
rect 15200 17110 15252 17162
rect 15304 17110 15356 17162
rect 15408 17110 15460 17162
rect 24524 17110 24576 17162
rect 24628 17110 24680 17162
rect 24732 17110 24784 17162
rect 33848 17110 33900 17162
rect 33952 17110 34004 17162
rect 34056 17110 34108 17162
rect 10538 16102 10590 16154
rect 10642 16102 10694 16154
rect 10746 16102 10798 16154
rect 19862 16102 19914 16154
rect 19966 16102 20018 16154
rect 20070 16102 20122 16154
rect 29186 16102 29238 16154
rect 29290 16102 29342 16154
rect 29394 16102 29446 16154
rect 38510 16102 38562 16154
rect 38614 16102 38666 16154
rect 38718 16102 38770 16154
rect 5876 15094 5928 15146
rect 5980 15094 6032 15146
rect 6084 15094 6136 15146
rect 15200 15094 15252 15146
rect 15304 15094 15356 15146
rect 15408 15094 15460 15146
rect 24524 15094 24576 15146
rect 24628 15094 24680 15146
rect 24732 15094 24784 15146
rect 33848 15094 33900 15146
rect 33952 15094 34004 15146
rect 34056 15094 34108 15146
rect 10538 14086 10590 14138
rect 10642 14086 10694 14138
rect 10746 14086 10798 14138
rect 19862 14086 19914 14138
rect 19966 14086 20018 14138
rect 20070 14086 20122 14138
rect 29186 14086 29238 14138
rect 29290 14086 29342 14138
rect 29394 14086 29446 14138
rect 38510 14086 38562 14138
rect 38614 14086 38666 14138
rect 38718 14086 38770 14138
rect 5876 13078 5928 13130
rect 5980 13078 6032 13130
rect 6084 13078 6136 13130
rect 15200 13078 15252 13130
rect 15304 13078 15356 13130
rect 15408 13078 15460 13130
rect 24524 13078 24576 13130
rect 24628 13078 24680 13130
rect 24732 13078 24784 13130
rect 33848 13078 33900 13130
rect 33952 13078 34004 13130
rect 34056 13078 34108 13130
rect 10538 12070 10590 12122
rect 10642 12070 10694 12122
rect 10746 12070 10798 12122
rect 19862 12070 19914 12122
rect 19966 12070 20018 12122
rect 20070 12070 20122 12122
rect 29186 12070 29238 12122
rect 29290 12070 29342 12122
rect 29394 12070 29446 12122
rect 38510 12070 38562 12122
rect 38614 12070 38666 12122
rect 38718 12070 38770 12122
rect 5876 11062 5928 11114
rect 5980 11062 6032 11114
rect 6084 11062 6136 11114
rect 15200 11062 15252 11114
rect 15304 11062 15356 11114
rect 15408 11062 15460 11114
rect 24524 11062 24576 11114
rect 24628 11062 24680 11114
rect 24732 11062 24784 11114
rect 33848 11062 33900 11114
rect 33952 11062 34004 11114
rect 34056 11062 34108 11114
rect 10538 10054 10590 10106
rect 10642 10054 10694 10106
rect 10746 10054 10798 10106
rect 19862 10054 19914 10106
rect 19966 10054 20018 10106
rect 20070 10054 20122 10106
rect 29186 10054 29238 10106
rect 29290 10054 29342 10106
rect 29394 10054 29446 10106
rect 38510 10054 38562 10106
rect 38614 10054 38666 10106
rect 38718 10054 38770 10106
rect 5876 9046 5928 9098
rect 5980 9046 6032 9098
rect 6084 9046 6136 9098
rect 15200 9046 15252 9098
rect 15304 9046 15356 9098
rect 15408 9046 15460 9098
rect 24524 9046 24576 9098
rect 24628 9046 24680 9098
rect 24732 9046 24784 9098
rect 33848 9046 33900 9098
rect 33952 9046 34004 9098
rect 34056 9046 34108 9098
rect 10538 8038 10590 8090
rect 10642 8038 10694 8090
rect 10746 8038 10798 8090
rect 19862 8038 19914 8090
rect 19966 8038 20018 8090
rect 20070 8038 20122 8090
rect 29186 8038 29238 8090
rect 29290 8038 29342 8090
rect 29394 8038 29446 8090
rect 38510 8038 38562 8090
rect 38614 8038 38666 8090
rect 38718 8038 38770 8090
rect 5876 7030 5928 7082
rect 5980 7030 6032 7082
rect 6084 7030 6136 7082
rect 15200 7030 15252 7082
rect 15304 7030 15356 7082
rect 15408 7030 15460 7082
rect 24524 7030 24576 7082
rect 24628 7030 24680 7082
rect 24732 7030 24784 7082
rect 33848 7030 33900 7082
rect 33952 7030 34004 7082
rect 34056 7030 34108 7082
rect 10538 6022 10590 6074
rect 10642 6022 10694 6074
rect 10746 6022 10798 6074
rect 19862 6022 19914 6074
rect 19966 6022 20018 6074
rect 20070 6022 20122 6074
rect 29186 6022 29238 6074
rect 29290 6022 29342 6074
rect 29394 6022 29446 6074
rect 38510 6022 38562 6074
rect 38614 6022 38666 6074
rect 38718 6022 38770 6074
rect 5876 5014 5928 5066
rect 5980 5014 6032 5066
rect 6084 5014 6136 5066
rect 15200 5014 15252 5066
rect 15304 5014 15356 5066
rect 15408 5014 15460 5066
rect 24524 5014 24576 5066
rect 24628 5014 24680 5066
rect 24732 5014 24784 5066
rect 33848 5014 33900 5066
rect 33952 5014 34004 5066
rect 34056 5014 34108 5066
rect 10538 4006 10590 4058
rect 10642 4006 10694 4058
rect 10746 4006 10798 4058
rect 19862 4006 19914 4058
rect 19966 4006 20018 4058
rect 20070 4006 20122 4058
rect 29186 4006 29238 4058
rect 29290 4006 29342 4058
rect 29394 4006 29446 4058
rect 38510 4006 38562 4058
rect 38614 4006 38666 4058
rect 38718 4006 38770 4058
<< metal2 >>
rect 14784 39200 14896 40000
rect 15456 39200 15568 40000
rect 10536 36316 10800 36326
rect 10592 36260 10640 36316
rect 10696 36260 10744 36316
rect 10536 36250 10800 36260
rect 5874 35308 6138 35318
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 5874 35242 6138 35252
rect 10536 34300 10800 34310
rect 10592 34244 10640 34300
rect 10696 34244 10744 34300
rect 10536 34234 10800 34244
rect 5874 33292 6138 33302
rect 5930 33236 5978 33292
rect 6034 33236 6082 33292
rect 5874 33226 6138 33236
rect 10536 32284 10800 32294
rect 10592 32228 10640 32284
rect 10696 32228 10744 32284
rect 10536 32218 10800 32228
rect 14812 31948 14868 39200
rect 15484 35700 15540 39200
rect 19860 36316 20124 36326
rect 19916 36260 19964 36316
rect 20020 36260 20068 36316
rect 19860 36250 20124 36260
rect 29184 36316 29448 36326
rect 29240 36260 29288 36316
rect 29344 36260 29392 36316
rect 29184 36250 29448 36260
rect 38508 36316 38772 36326
rect 38564 36260 38612 36316
rect 38668 36260 38716 36316
rect 38508 36250 38772 36260
rect 15484 35644 15652 35700
rect 15198 35308 15462 35318
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15198 35242 15462 35252
rect 15198 33292 15462 33302
rect 15254 33236 15302 33292
rect 15358 33236 15406 33292
rect 15198 33226 15462 33236
rect 15484 32116 15540 32126
rect 15596 32116 15652 35644
rect 24522 35308 24786 35318
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24522 35242 24786 35252
rect 33846 35308 34110 35318
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 33846 35242 34110 35252
rect 19860 34300 20124 34310
rect 19916 34244 19964 34300
rect 20020 34244 20068 34300
rect 19860 34234 20124 34244
rect 29184 34300 29448 34310
rect 29240 34244 29288 34300
rect 29344 34244 29392 34300
rect 29184 34234 29448 34244
rect 38508 34300 38772 34310
rect 38564 34244 38612 34300
rect 38668 34244 38716 34300
rect 38508 34234 38772 34244
rect 24522 33292 24786 33302
rect 24578 33236 24626 33292
rect 24682 33236 24730 33292
rect 24522 33226 24786 33236
rect 33846 33292 34110 33302
rect 33902 33236 33950 33292
rect 34006 33236 34054 33292
rect 33846 33226 34110 33236
rect 19860 32284 20124 32294
rect 19916 32228 19964 32284
rect 20020 32228 20068 32284
rect 19860 32218 20124 32228
rect 29184 32284 29448 32294
rect 29240 32228 29288 32284
rect 29344 32228 29392 32284
rect 29184 32218 29448 32228
rect 38508 32284 38772 32294
rect 38564 32228 38612 32284
rect 38668 32228 38716 32284
rect 38508 32218 38772 32228
rect 15484 32114 15652 32116
rect 15484 32062 15486 32114
rect 15538 32062 15652 32114
rect 15484 32060 15652 32062
rect 15484 32050 15540 32060
rect 14812 31892 14980 31948
rect 15148 31892 15204 31902
rect 14924 31890 15204 31892
rect 14924 31838 14926 31890
rect 14978 31838 15150 31890
rect 15202 31838 15204 31890
rect 14924 31836 15204 31838
rect 14924 31826 14980 31836
rect 15148 31826 15204 31836
rect 5874 31276 6138 31286
rect 5930 31220 5978 31276
rect 6034 31220 6082 31276
rect 5874 31210 6138 31220
rect 15198 31276 15462 31286
rect 15254 31220 15302 31276
rect 15358 31220 15406 31276
rect 15198 31210 15462 31220
rect 24522 31276 24786 31286
rect 24578 31220 24626 31276
rect 24682 31220 24730 31276
rect 24522 31210 24786 31220
rect 33846 31276 34110 31286
rect 33902 31220 33950 31276
rect 34006 31220 34054 31276
rect 33846 31210 34110 31220
rect 10536 30268 10800 30278
rect 10592 30212 10640 30268
rect 10696 30212 10744 30268
rect 10536 30202 10800 30212
rect 19860 30268 20124 30278
rect 19916 30212 19964 30268
rect 20020 30212 20068 30268
rect 19860 30202 20124 30212
rect 29184 30268 29448 30278
rect 29240 30212 29288 30268
rect 29344 30212 29392 30268
rect 29184 30202 29448 30212
rect 38508 30268 38772 30278
rect 38564 30212 38612 30268
rect 38668 30212 38716 30268
rect 38508 30202 38772 30212
rect 5874 29260 6138 29270
rect 5930 29204 5978 29260
rect 6034 29204 6082 29260
rect 5874 29194 6138 29204
rect 15198 29260 15462 29270
rect 15254 29204 15302 29260
rect 15358 29204 15406 29260
rect 15198 29194 15462 29204
rect 24522 29260 24786 29270
rect 24578 29204 24626 29260
rect 24682 29204 24730 29260
rect 24522 29194 24786 29204
rect 33846 29260 34110 29270
rect 33902 29204 33950 29260
rect 34006 29204 34054 29260
rect 33846 29194 34110 29204
rect 10536 28252 10800 28262
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10536 28186 10800 28196
rect 19860 28252 20124 28262
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 19860 28186 20124 28196
rect 29184 28252 29448 28262
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29184 28186 29448 28196
rect 38508 28252 38772 28262
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38508 28186 38772 28196
rect 5874 27244 6138 27254
rect 5930 27188 5978 27244
rect 6034 27188 6082 27244
rect 5874 27178 6138 27188
rect 15198 27244 15462 27254
rect 15254 27188 15302 27244
rect 15358 27188 15406 27244
rect 15198 27178 15462 27188
rect 24522 27244 24786 27254
rect 24578 27188 24626 27244
rect 24682 27188 24730 27244
rect 24522 27178 24786 27188
rect 33846 27244 34110 27254
rect 33902 27188 33950 27244
rect 34006 27188 34054 27244
rect 33846 27178 34110 27188
rect 10536 26236 10800 26246
rect 10592 26180 10640 26236
rect 10696 26180 10744 26236
rect 10536 26170 10800 26180
rect 19860 26236 20124 26246
rect 19916 26180 19964 26236
rect 20020 26180 20068 26236
rect 19860 26170 20124 26180
rect 29184 26236 29448 26246
rect 29240 26180 29288 26236
rect 29344 26180 29392 26236
rect 29184 26170 29448 26180
rect 38508 26236 38772 26246
rect 38564 26180 38612 26236
rect 38668 26180 38716 26236
rect 38508 26170 38772 26180
rect 34524 25620 34580 25630
rect 5874 25228 6138 25238
rect 5930 25172 5978 25228
rect 6034 25172 6082 25228
rect 5874 25162 6138 25172
rect 15198 25228 15462 25238
rect 15254 25172 15302 25228
rect 15358 25172 15406 25228
rect 15198 25162 15462 25172
rect 24522 25228 24786 25238
rect 24578 25172 24626 25228
rect 24682 25172 24730 25228
rect 24522 25162 24786 25172
rect 33846 25228 34110 25238
rect 33902 25172 33950 25228
rect 34006 25172 34054 25228
rect 33846 25162 34110 25172
rect 4172 24276 4228 24286
rect 4060 23604 4116 23614
rect 4060 20580 4116 23548
rect 4172 22708 4228 24220
rect 10536 24220 10800 24230
rect 10592 24164 10640 24220
rect 10696 24164 10744 24220
rect 10536 24154 10800 24164
rect 19860 24220 20124 24230
rect 19916 24164 19964 24220
rect 20020 24164 20068 24220
rect 19860 24154 20124 24164
rect 29184 24220 29448 24230
rect 29240 24164 29288 24220
rect 29344 24164 29392 24220
rect 29184 24154 29448 24164
rect 5874 23212 6138 23222
rect 5930 23156 5978 23212
rect 6034 23156 6082 23212
rect 5874 23146 6138 23156
rect 15198 23212 15462 23222
rect 15254 23156 15302 23212
rect 15358 23156 15406 23212
rect 15198 23146 15462 23156
rect 24522 23212 24786 23222
rect 24578 23156 24626 23212
rect 24682 23156 24730 23212
rect 24522 23146 24786 23156
rect 33846 23212 34110 23222
rect 33902 23156 33950 23212
rect 34006 23156 34054 23212
rect 33846 23146 34110 23156
rect 4172 22642 4228 22652
rect 4284 22932 4340 22942
rect 4284 20692 4340 22876
rect 13580 22708 13636 22718
rect 10536 22204 10800 22214
rect 10592 22148 10640 22204
rect 10696 22148 10744 22204
rect 10536 22138 10800 22148
rect 5874 21196 6138 21206
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 5874 21130 6138 21140
rect 4284 20626 4340 20636
rect 4060 20514 4116 20524
rect 12460 20468 12516 20478
rect 12460 20374 12516 20412
rect 12908 20466 12964 20478
rect 12908 20414 12910 20466
rect 12962 20414 12964 20466
rect 4620 20356 4676 20366
rect 4060 18788 4116 18798
rect 4060 16212 4116 18732
rect 4284 18676 4340 18686
rect 4172 18564 4228 18574
rect 4172 17556 4228 18508
rect 4172 17490 4228 17500
rect 4284 16884 4340 18620
rect 4620 18228 4676 20300
rect 12908 20356 12964 20414
rect 12908 20290 12964 20300
rect 13468 20466 13524 20478
rect 13468 20414 13470 20466
rect 13522 20414 13524 20466
rect 10536 20188 10800 20198
rect 13468 20188 13524 20414
rect 10592 20132 10640 20188
rect 10696 20132 10744 20188
rect 10536 20122 10800 20132
rect 12908 20132 13524 20188
rect 13580 20188 13636 22652
rect 19860 22204 20124 22214
rect 19916 22148 19964 22204
rect 20020 22148 20068 22204
rect 19860 22138 20124 22148
rect 29184 22204 29448 22214
rect 29240 22148 29288 22204
rect 29344 22148 29392 22204
rect 29184 22138 29448 22148
rect 17948 21924 18004 21934
rect 15198 21196 15462 21206
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15198 21130 15462 21140
rect 13692 20802 13748 20814
rect 13692 20750 13694 20802
rect 13746 20750 13748 20802
rect 13692 20468 13748 20750
rect 13692 20402 13748 20412
rect 13916 20690 13972 20702
rect 13916 20638 13918 20690
rect 13970 20638 13972 20690
rect 13804 20356 13860 20366
rect 13916 20356 13972 20638
rect 13860 20300 13972 20356
rect 14924 20692 14980 20702
rect 13804 20290 13860 20300
rect 13580 20132 13972 20188
rect 12684 19794 12740 19806
rect 12684 19742 12686 19794
rect 12738 19742 12740 19794
rect 5874 19180 6138 19190
rect 5930 19124 5978 19180
rect 6034 19124 6082 19180
rect 5874 19114 6138 19124
rect 12684 18898 12740 19742
rect 12908 19794 12964 20132
rect 12908 19742 12910 19794
rect 12962 19742 12964 19794
rect 12908 19730 12964 19742
rect 13804 19682 13860 19694
rect 13804 19630 13806 19682
rect 13858 19630 13860 19682
rect 12684 18846 12686 18898
rect 12738 18846 12740 18898
rect 12684 18834 12740 18846
rect 13468 19572 13524 19582
rect 11564 18676 11620 18686
rect 11564 18582 11620 18620
rect 12012 18674 12068 18686
rect 12012 18622 12014 18674
rect 12066 18622 12068 18674
rect 11116 18564 11172 18574
rect 11116 18470 11172 18508
rect 12012 18564 12068 18622
rect 12124 18676 12180 18686
rect 12124 18582 12180 18620
rect 12012 18498 12068 18508
rect 4620 18162 4676 18172
rect 10536 18172 10800 18182
rect 10592 18116 10640 18172
rect 10696 18116 10744 18172
rect 10536 18106 10800 18116
rect 13468 17890 13524 19516
rect 13804 18786 13860 19630
rect 13804 18734 13806 18786
rect 13858 18734 13860 18786
rect 13804 18722 13860 18734
rect 13468 17838 13470 17890
rect 13522 17838 13524 17890
rect 13468 17826 13524 17838
rect 13916 18674 13972 20132
rect 14252 19684 14308 19694
rect 14700 19684 14756 19694
rect 14252 19682 14756 19684
rect 14252 19630 14254 19682
rect 14306 19630 14702 19682
rect 14754 19630 14756 19682
rect 14252 19628 14756 19630
rect 14252 19618 14308 19628
rect 14700 19618 14756 19628
rect 14924 19682 14980 20636
rect 17612 20580 17668 20590
rect 17612 20466 17668 20524
rect 17612 20414 17614 20466
rect 17666 20414 17668 20466
rect 16716 19908 16772 19918
rect 16716 19814 16772 19852
rect 17612 19906 17668 20414
rect 17948 20188 18004 21868
rect 31052 21924 31108 21934
rect 22092 21812 22148 21822
rect 19292 21588 19348 21598
rect 19292 21026 19348 21532
rect 19292 20974 19294 21026
rect 19346 20974 19348 21026
rect 19292 20962 19348 20974
rect 18060 20916 18116 20926
rect 18060 20822 18116 20860
rect 18396 20692 18452 20702
rect 18284 20690 18452 20692
rect 18284 20638 18398 20690
rect 18450 20638 18452 20690
rect 18284 20636 18452 20638
rect 18284 20580 18340 20636
rect 18396 20626 18452 20636
rect 18844 20690 18900 20702
rect 18844 20638 18846 20690
rect 18898 20638 18900 20690
rect 17948 20132 18228 20188
rect 17612 19854 17614 19906
rect 17666 19854 17668 19906
rect 17612 19842 17668 19854
rect 16492 19796 16548 19806
rect 16492 19794 16660 19796
rect 16492 19742 16494 19794
rect 16546 19742 16660 19794
rect 16492 19740 16660 19742
rect 16492 19730 16548 19740
rect 14924 19630 14926 19682
rect 14978 19630 14980 19682
rect 14924 19618 14980 19630
rect 14028 19572 14084 19582
rect 14084 19516 14196 19572
rect 14028 19506 14084 19516
rect 13916 18622 13918 18674
rect 13970 18622 13972 18674
rect 13916 17890 13972 18622
rect 14140 18674 14196 19516
rect 15198 19180 15462 19190
rect 15254 19124 15302 19180
rect 15358 19124 15406 19180
rect 15198 19114 15462 19124
rect 15932 18900 15988 18910
rect 15932 18786 15988 18844
rect 15932 18734 15934 18786
rect 15986 18734 15988 18786
rect 15932 18722 15988 18734
rect 16268 18788 16324 18798
rect 16268 18694 16324 18732
rect 14140 18622 14142 18674
rect 14194 18622 14196 18674
rect 14140 18610 14196 18622
rect 16604 18674 16660 19740
rect 18172 19570 18228 20132
rect 18284 19682 18340 20524
rect 18844 20580 18900 20638
rect 21868 20690 21924 20702
rect 21868 20638 21870 20690
rect 21922 20638 21924 20690
rect 19404 20580 19460 20590
rect 18844 20578 19460 20580
rect 18844 20526 19406 20578
rect 19458 20526 19460 20578
rect 18844 20524 19460 20526
rect 18844 19908 18900 20524
rect 19404 20188 19460 20524
rect 20412 20578 20468 20590
rect 20412 20526 20414 20578
rect 20466 20526 20468 20578
rect 19860 20188 20124 20198
rect 20412 20188 20468 20526
rect 20860 20580 20916 20590
rect 20748 20356 20804 20366
rect 20748 20262 20804 20300
rect 19404 20132 19572 20188
rect 18844 19842 18900 19852
rect 18284 19630 18286 19682
rect 18338 19630 18340 19682
rect 18284 19618 18340 19630
rect 19516 19682 19572 20132
rect 19916 20132 19964 20188
rect 20020 20132 20068 20188
rect 19860 20122 20124 20132
rect 20188 20132 20468 20188
rect 20188 20020 20244 20132
rect 20076 19964 20244 20020
rect 20076 19906 20132 19964
rect 20076 19854 20078 19906
rect 20130 19854 20132 19906
rect 20076 19842 20132 19854
rect 19516 19630 19518 19682
rect 19570 19630 19572 19682
rect 19516 19618 19572 19630
rect 18172 19518 18174 19570
rect 18226 19518 18228 19570
rect 16828 18900 16884 18910
rect 16828 18786 16884 18844
rect 16828 18734 16830 18786
rect 16882 18734 16884 18786
rect 16828 18722 16884 18734
rect 16940 18788 16996 18798
rect 16996 18732 17108 18788
rect 16940 18722 16996 18732
rect 16604 18622 16606 18674
rect 16658 18622 16660 18674
rect 16604 18610 16660 18622
rect 17052 18674 17108 18732
rect 18172 18786 18228 19518
rect 20860 19570 20916 20524
rect 21868 20468 21924 20638
rect 22092 20690 22148 21756
rect 27356 21588 27412 21598
rect 24522 21196 24786 21206
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24522 21130 24786 21140
rect 25116 20916 25172 20926
rect 22092 20638 22094 20690
rect 22146 20638 22148 20690
rect 21980 20468 22036 20478
rect 21868 20412 21980 20468
rect 21980 20402 22036 20412
rect 21532 20356 21588 20366
rect 21532 20188 21588 20300
rect 22092 20188 22148 20638
rect 22316 20692 22372 20702
rect 22316 20598 22372 20636
rect 23436 20580 23492 20590
rect 23436 20486 23492 20524
rect 24332 20580 24388 20590
rect 24332 20486 24388 20524
rect 22876 20468 22932 20478
rect 22876 20188 22932 20412
rect 23772 20356 23828 20366
rect 21532 20132 22148 20188
rect 22652 20132 22932 20188
rect 23660 20354 23828 20356
rect 23660 20302 23774 20354
rect 23826 20302 23828 20354
rect 23660 20300 23828 20302
rect 23660 20244 23716 20300
rect 23772 20290 23828 20300
rect 21532 19682 21588 20132
rect 22652 19794 22708 20132
rect 22652 19742 22654 19794
rect 22706 19742 22708 19794
rect 22652 19730 22708 19742
rect 22876 19908 22932 19918
rect 21532 19630 21534 19682
rect 21586 19630 21588 19682
rect 21532 19618 21588 19630
rect 20860 19518 20862 19570
rect 20914 19518 20916 19570
rect 20860 19506 20916 19518
rect 22876 19570 22932 19852
rect 23660 19682 23716 20188
rect 25116 20244 25172 20860
rect 26124 20578 26180 20590
rect 26124 20526 26126 20578
rect 26178 20526 26180 20578
rect 26124 20188 26180 20526
rect 23660 19630 23662 19682
rect 23714 19630 23716 19682
rect 23660 19618 23716 19630
rect 24220 19682 24276 19694
rect 24220 19630 24222 19682
rect 24274 19630 24276 19682
rect 24220 19572 24276 19630
rect 24668 19684 24724 19694
rect 24668 19682 24948 19684
rect 24668 19630 24670 19682
rect 24722 19630 24948 19682
rect 24668 19628 24948 19630
rect 24668 19618 24724 19628
rect 24332 19572 24388 19582
rect 22876 19518 22878 19570
rect 22930 19518 22932 19570
rect 22876 19506 22932 19518
rect 23772 19516 24332 19572
rect 18172 18734 18174 18786
rect 18226 18734 18228 18786
rect 18172 18722 18228 18734
rect 23436 18786 23492 18798
rect 23436 18734 23438 18786
rect 23490 18734 23492 18786
rect 17052 18622 17054 18674
rect 17106 18622 17108 18674
rect 17052 18610 17108 18622
rect 19860 18172 20124 18182
rect 19916 18116 19964 18172
rect 20020 18116 20068 18172
rect 19860 18106 20124 18116
rect 13916 17838 13918 17890
rect 13970 17838 13972 17890
rect 13916 17826 13972 17838
rect 23436 17556 23492 18734
rect 23660 18564 23716 18574
rect 23772 18564 23828 19516
rect 24332 19506 24388 19516
rect 24522 19180 24786 19190
rect 24578 19124 24626 19180
rect 24682 19124 24730 19180
rect 24522 19114 24786 19124
rect 23660 18562 23828 18564
rect 23660 18510 23662 18562
rect 23714 18510 23828 18562
rect 23660 18508 23828 18510
rect 23660 18498 23716 18508
rect 23436 17490 23492 17500
rect 5874 17164 6138 17174
rect 5930 17108 5978 17164
rect 6034 17108 6082 17164
rect 5874 17098 6138 17108
rect 15198 17164 15462 17174
rect 15254 17108 15302 17164
rect 15358 17108 15406 17164
rect 15198 17098 15462 17108
rect 24522 17164 24786 17174
rect 24578 17108 24626 17164
rect 24682 17108 24730 17164
rect 24522 17098 24786 17108
rect 4284 16818 4340 16828
rect 4060 16146 4116 16156
rect 10536 16156 10800 16166
rect 10592 16100 10640 16156
rect 10696 16100 10744 16156
rect 10536 16090 10800 16100
rect 19860 16156 20124 16166
rect 19916 16100 19964 16156
rect 20020 16100 20068 16156
rect 19860 16090 20124 16100
rect 24892 15540 24948 19628
rect 25116 18674 25172 20188
rect 25564 20132 26180 20188
rect 26460 20354 26516 20366
rect 26460 20302 26462 20354
rect 26514 20302 26516 20354
rect 26460 20244 26516 20302
rect 26460 20178 26516 20188
rect 27244 20244 27300 20254
rect 25340 19908 25396 19918
rect 25340 19814 25396 19852
rect 25564 18786 25620 20132
rect 26908 19881 26964 19893
rect 26908 19829 26910 19881
rect 26962 19829 26964 19881
rect 25564 18734 25566 18786
rect 25618 18734 25620 18786
rect 25564 18722 25620 18734
rect 25788 19572 25844 19582
rect 25788 18788 25844 19516
rect 26348 19572 26404 19582
rect 26348 19478 26404 19516
rect 26012 18788 26068 18798
rect 25788 18732 26012 18788
rect 26012 18694 26068 18732
rect 25116 18622 25118 18674
rect 25170 18622 25172 18674
rect 25116 18610 25172 18622
rect 26908 18674 26964 19829
rect 26908 18622 26910 18674
rect 26962 18622 26964 18674
rect 26908 18564 26964 18622
rect 27244 18674 27300 20188
rect 27356 18786 27412 21532
rect 31052 20914 31108 21868
rect 33846 21196 34110 21206
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 33846 21130 34110 21140
rect 31052 20862 31054 20914
rect 31106 20862 31108 20914
rect 31052 20850 31108 20862
rect 28140 20804 28196 20814
rect 28140 20244 28196 20748
rect 29148 20580 29204 20590
rect 28028 20132 28196 20188
rect 28476 20578 29204 20580
rect 28476 20526 29150 20578
rect 29202 20526 29204 20578
rect 28476 20524 29204 20526
rect 28028 19682 28084 20132
rect 28028 19630 28030 19682
rect 28082 19630 28084 19682
rect 28028 19618 28084 19630
rect 28476 19570 28532 20524
rect 29148 20514 29204 20524
rect 30716 20578 30772 20590
rect 30716 20526 30718 20578
rect 30770 20526 30772 20578
rect 30044 20466 30100 20478
rect 30044 20414 30046 20466
rect 30098 20414 30100 20466
rect 28476 19518 28478 19570
rect 28530 19518 28532 19570
rect 28476 19506 28532 19518
rect 28924 20356 28980 20366
rect 28924 19570 28980 20300
rect 29484 20356 29540 20366
rect 29596 20356 29652 20366
rect 29484 20354 29596 20356
rect 29484 20302 29486 20354
rect 29538 20302 29596 20354
rect 29484 20300 29596 20302
rect 29484 20290 29540 20300
rect 29184 20188 29448 20198
rect 29240 20132 29288 20188
rect 29344 20132 29392 20188
rect 29184 20122 29448 20132
rect 28924 19518 28926 19570
rect 28978 19518 28980 19570
rect 28924 19506 28980 19518
rect 29372 19684 29428 19694
rect 29596 19684 29652 20300
rect 29372 19682 29652 19684
rect 29372 19630 29374 19682
rect 29426 19630 29652 19682
rect 29372 19628 29652 19630
rect 27356 18734 27358 18786
rect 27410 18734 27412 18786
rect 27356 18722 27412 18734
rect 29372 18786 29428 19628
rect 30044 19572 30100 20414
rect 30716 20468 30772 20526
rect 30716 20402 30772 20412
rect 34300 20580 34356 20590
rect 30940 20020 30996 20030
rect 30044 18900 30100 19516
rect 30044 18834 30100 18844
rect 30716 19794 30772 19806
rect 30716 19742 30718 19794
rect 30770 19742 30772 19794
rect 30716 19572 30772 19742
rect 29372 18734 29374 18786
rect 29426 18734 29428 18786
rect 29372 18722 29428 18734
rect 27244 18622 27246 18674
rect 27298 18622 27300 18674
rect 27244 18610 27300 18622
rect 29708 18676 29764 18686
rect 29708 18582 29764 18620
rect 30604 18676 30660 18686
rect 30716 18676 30772 19516
rect 30940 19570 30996 19964
rect 31948 20020 32004 20030
rect 31948 19906 32004 19964
rect 31948 19854 31950 19906
rect 32002 19854 32004 19906
rect 31948 19842 32004 19854
rect 30940 19518 30942 19570
rect 30994 19518 30996 19570
rect 30940 19506 30996 19518
rect 31500 19572 31556 19582
rect 31500 19478 31556 19516
rect 33846 19180 34110 19190
rect 33902 19124 33950 19180
rect 34006 19124 34054 19180
rect 33846 19114 34110 19124
rect 30660 18620 30772 18676
rect 30604 18582 30660 18620
rect 26908 18498 26964 18508
rect 27916 18564 27972 18574
rect 27916 18470 27972 18508
rect 28588 18564 28644 18574
rect 28588 18470 28644 18508
rect 30044 18452 30100 18462
rect 30044 18358 30100 18396
rect 29184 18172 29448 18182
rect 29240 18116 29288 18172
rect 29344 18116 29392 18172
rect 29184 18106 29448 18116
rect 26012 17556 26068 17566
rect 26012 17462 26068 17500
rect 33846 17164 34110 17174
rect 33902 17108 33950 17164
rect 34006 17108 34054 17164
rect 33846 17098 34110 17108
rect 29184 16156 29448 16166
rect 29240 16100 29288 16156
rect 29344 16100 29392 16156
rect 29184 16090 29448 16100
rect 24892 15474 24948 15484
rect 5874 15148 6138 15158
rect 5930 15092 5978 15148
rect 6034 15092 6082 15148
rect 5874 15082 6138 15092
rect 15198 15148 15462 15158
rect 15254 15092 15302 15148
rect 15358 15092 15406 15148
rect 15198 15082 15462 15092
rect 24522 15148 24786 15158
rect 24578 15092 24626 15148
rect 24682 15092 24730 15148
rect 24522 15082 24786 15092
rect 33846 15148 34110 15158
rect 33902 15092 33950 15148
rect 34006 15092 34054 15148
rect 33846 15082 34110 15092
rect 34300 14868 34356 20524
rect 34524 19908 34580 25564
rect 34748 24948 34804 24958
rect 34748 20804 34804 24892
rect 38508 24220 38772 24230
rect 38564 24164 38612 24220
rect 38668 24164 38716 24220
rect 38508 24154 38772 24164
rect 35084 24052 35140 24062
rect 34972 22932 35028 22942
rect 34748 20738 34804 20748
rect 34860 22036 34916 22046
rect 34860 20692 34916 21980
rect 34972 20916 35028 22876
rect 35084 21812 35140 23996
rect 35196 23604 35252 23614
rect 35196 21924 35252 23548
rect 38508 22204 38772 22214
rect 38564 22148 38612 22204
rect 38668 22148 38716 22204
rect 38508 22138 38772 22148
rect 35196 21858 35252 21868
rect 35084 21746 35140 21756
rect 34972 20850 35028 20860
rect 34860 20626 34916 20636
rect 34636 20356 34692 20366
rect 34636 20020 34692 20300
rect 38508 20188 38772 20198
rect 38564 20132 38612 20188
rect 38668 20132 38716 20188
rect 38508 20122 38772 20132
rect 34636 19954 34692 19964
rect 34524 19842 34580 19852
rect 35084 18900 35140 18910
rect 35084 16324 35140 18844
rect 35196 18788 35252 18798
rect 35196 16884 35252 18732
rect 38508 18172 38772 18182
rect 38564 18116 38612 18172
rect 38668 18116 38716 18172
rect 38508 18106 38772 18116
rect 35196 16818 35252 16828
rect 35084 16258 35140 16268
rect 38508 16156 38772 16166
rect 38564 16100 38612 16156
rect 38668 16100 38716 16156
rect 38508 16090 38772 16100
rect 34300 14802 34356 14812
rect 10536 14140 10800 14150
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10536 14074 10800 14084
rect 19860 14140 20124 14150
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 19860 14074 20124 14084
rect 29184 14140 29448 14150
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29184 14074 29448 14084
rect 38508 14140 38772 14150
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38508 14074 38772 14084
rect 5874 13132 6138 13142
rect 5930 13076 5978 13132
rect 6034 13076 6082 13132
rect 5874 13066 6138 13076
rect 15198 13132 15462 13142
rect 15254 13076 15302 13132
rect 15358 13076 15406 13132
rect 15198 13066 15462 13076
rect 24522 13132 24786 13142
rect 24578 13076 24626 13132
rect 24682 13076 24730 13132
rect 24522 13066 24786 13076
rect 33846 13132 34110 13142
rect 33902 13076 33950 13132
rect 34006 13076 34054 13132
rect 33846 13066 34110 13076
rect 10536 12124 10800 12134
rect 10592 12068 10640 12124
rect 10696 12068 10744 12124
rect 10536 12058 10800 12068
rect 19860 12124 20124 12134
rect 19916 12068 19964 12124
rect 20020 12068 20068 12124
rect 19860 12058 20124 12068
rect 29184 12124 29448 12134
rect 29240 12068 29288 12124
rect 29344 12068 29392 12124
rect 29184 12058 29448 12068
rect 38508 12124 38772 12134
rect 38564 12068 38612 12124
rect 38668 12068 38716 12124
rect 38508 12058 38772 12068
rect 5874 11116 6138 11126
rect 5930 11060 5978 11116
rect 6034 11060 6082 11116
rect 5874 11050 6138 11060
rect 15198 11116 15462 11126
rect 15254 11060 15302 11116
rect 15358 11060 15406 11116
rect 15198 11050 15462 11060
rect 24522 11116 24786 11126
rect 24578 11060 24626 11116
rect 24682 11060 24730 11116
rect 24522 11050 24786 11060
rect 33846 11116 34110 11126
rect 33902 11060 33950 11116
rect 34006 11060 34054 11116
rect 33846 11050 34110 11060
rect 10536 10108 10800 10118
rect 10592 10052 10640 10108
rect 10696 10052 10744 10108
rect 10536 10042 10800 10052
rect 19860 10108 20124 10118
rect 19916 10052 19964 10108
rect 20020 10052 20068 10108
rect 19860 10042 20124 10052
rect 29184 10108 29448 10118
rect 29240 10052 29288 10108
rect 29344 10052 29392 10108
rect 29184 10042 29448 10052
rect 38508 10108 38772 10118
rect 38564 10052 38612 10108
rect 38668 10052 38716 10108
rect 38508 10042 38772 10052
rect 5874 9100 6138 9110
rect 5930 9044 5978 9100
rect 6034 9044 6082 9100
rect 5874 9034 6138 9044
rect 15198 9100 15462 9110
rect 15254 9044 15302 9100
rect 15358 9044 15406 9100
rect 15198 9034 15462 9044
rect 24522 9100 24786 9110
rect 24578 9044 24626 9100
rect 24682 9044 24730 9100
rect 24522 9034 24786 9044
rect 33846 9100 34110 9110
rect 33902 9044 33950 9100
rect 34006 9044 34054 9100
rect 33846 9034 34110 9044
rect 10536 8092 10800 8102
rect 10592 8036 10640 8092
rect 10696 8036 10744 8092
rect 10536 8026 10800 8036
rect 19860 8092 20124 8102
rect 19916 8036 19964 8092
rect 20020 8036 20068 8092
rect 19860 8026 20124 8036
rect 29184 8092 29448 8102
rect 29240 8036 29288 8092
rect 29344 8036 29392 8092
rect 29184 8026 29448 8036
rect 38508 8092 38772 8102
rect 38564 8036 38612 8092
rect 38668 8036 38716 8092
rect 38508 8026 38772 8036
rect 5874 7084 6138 7094
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 5874 7018 6138 7028
rect 15198 7084 15462 7094
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15198 7018 15462 7028
rect 24522 7084 24786 7094
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24522 7018 24786 7028
rect 33846 7084 34110 7094
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 33846 7018 34110 7028
rect 10536 6076 10800 6086
rect 10592 6020 10640 6076
rect 10696 6020 10744 6076
rect 10536 6010 10800 6020
rect 19860 6076 20124 6086
rect 19916 6020 19964 6076
rect 20020 6020 20068 6076
rect 19860 6010 20124 6020
rect 29184 6076 29448 6086
rect 29240 6020 29288 6076
rect 29344 6020 29392 6076
rect 29184 6010 29448 6020
rect 38508 6076 38772 6086
rect 38564 6020 38612 6076
rect 38668 6020 38716 6076
rect 38508 6010 38772 6020
rect 5874 5068 6138 5078
rect 5930 5012 5978 5068
rect 6034 5012 6082 5068
rect 5874 5002 6138 5012
rect 15198 5068 15462 5078
rect 15254 5012 15302 5068
rect 15358 5012 15406 5068
rect 15198 5002 15462 5012
rect 24522 5068 24786 5078
rect 24578 5012 24626 5068
rect 24682 5012 24730 5068
rect 24522 5002 24786 5012
rect 33846 5068 34110 5078
rect 33902 5012 33950 5068
rect 34006 5012 34054 5068
rect 33846 5002 34110 5012
rect 10536 4060 10800 4070
rect 10592 4004 10640 4060
rect 10696 4004 10744 4060
rect 10536 3994 10800 4004
rect 19860 4060 20124 4070
rect 19916 4004 19964 4060
rect 20020 4004 20068 4060
rect 19860 3994 20124 4004
rect 29184 4060 29448 4070
rect 29240 4004 29288 4060
rect 29344 4004 29392 4060
rect 29184 3994 29448 4004
rect 38508 4060 38772 4070
rect 38564 4004 38612 4060
rect 38668 4004 38716 4060
rect 38508 3994 38772 4004
<< via2 >>
rect 10536 36314 10592 36316
rect 10536 36262 10538 36314
rect 10538 36262 10590 36314
rect 10590 36262 10592 36314
rect 10536 36260 10592 36262
rect 10640 36314 10696 36316
rect 10640 36262 10642 36314
rect 10642 36262 10694 36314
rect 10694 36262 10696 36314
rect 10640 36260 10696 36262
rect 10744 36314 10800 36316
rect 10744 36262 10746 36314
rect 10746 36262 10798 36314
rect 10798 36262 10800 36314
rect 10744 36260 10800 36262
rect 5874 35306 5930 35308
rect 5874 35254 5876 35306
rect 5876 35254 5928 35306
rect 5928 35254 5930 35306
rect 5874 35252 5930 35254
rect 5978 35306 6034 35308
rect 5978 35254 5980 35306
rect 5980 35254 6032 35306
rect 6032 35254 6034 35306
rect 5978 35252 6034 35254
rect 6082 35306 6138 35308
rect 6082 35254 6084 35306
rect 6084 35254 6136 35306
rect 6136 35254 6138 35306
rect 6082 35252 6138 35254
rect 10536 34298 10592 34300
rect 10536 34246 10538 34298
rect 10538 34246 10590 34298
rect 10590 34246 10592 34298
rect 10536 34244 10592 34246
rect 10640 34298 10696 34300
rect 10640 34246 10642 34298
rect 10642 34246 10694 34298
rect 10694 34246 10696 34298
rect 10640 34244 10696 34246
rect 10744 34298 10800 34300
rect 10744 34246 10746 34298
rect 10746 34246 10798 34298
rect 10798 34246 10800 34298
rect 10744 34244 10800 34246
rect 5874 33290 5930 33292
rect 5874 33238 5876 33290
rect 5876 33238 5928 33290
rect 5928 33238 5930 33290
rect 5874 33236 5930 33238
rect 5978 33290 6034 33292
rect 5978 33238 5980 33290
rect 5980 33238 6032 33290
rect 6032 33238 6034 33290
rect 5978 33236 6034 33238
rect 6082 33290 6138 33292
rect 6082 33238 6084 33290
rect 6084 33238 6136 33290
rect 6136 33238 6138 33290
rect 6082 33236 6138 33238
rect 10536 32282 10592 32284
rect 10536 32230 10538 32282
rect 10538 32230 10590 32282
rect 10590 32230 10592 32282
rect 10536 32228 10592 32230
rect 10640 32282 10696 32284
rect 10640 32230 10642 32282
rect 10642 32230 10694 32282
rect 10694 32230 10696 32282
rect 10640 32228 10696 32230
rect 10744 32282 10800 32284
rect 10744 32230 10746 32282
rect 10746 32230 10798 32282
rect 10798 32230 10800 32282
rect 10744 32228 10800 32230
rect 19860 36314 19916 36316
rect 19860 36262 19862 36314
rect 19862 36262 19914 36314
rect 19914 36262 19916 36314
rect 19860 36260 19916 36262
rect 19964 36314 20020 36316
rect 19964 36262 19966 36314
rect 19966 36262 20018 36314
rect 20018 36262 20020 36314
rect 19964 36260 20020 36262
rect 20068 36314 20124 36316
rect 20068 36262 20070 36314
rect 20070 36262 20122 36314
rect 20122 36262 20124 36314
rect 20068 36260 20124 36262
rect 29184 36314 29240 36316
rect 29184 36262 29186 36314
rect 29186 36262 29238 36314
rect 29238 36262 29240 36314
rect 29184 36260 29240 36262
rect 29288 36314 29344 36316
rect 29288 36262 29290 36314
rect 29290 36262 29342 36314
rect 29342 36262 29344 36314
rect 29288 36260 29344 36262
rect 29392 36314 29448 36316
rect 29392 36262 29394 36314
rect 29394 36262 29446 36314
rect 29446 36262 29448 36314
rect 29392 36260 29448 36262
rect 38508 36314 38564 36316
rect 38508 36262 38510 36314
rect 38510 36262 38562 36314
rect 38562 36262 38564 36314
rect 38508 36260 38564 36262
rect 38612 36314 38668 36316
rect 38612 36262 38614 36314
rect 38614 36262 38666 36314
rect 38666 36262 38668 36314
rect 38612 36260 38668 36262
rect 38716 36314 38772 36316
rect 38716 36262 38718 36314
rect 38718 36262 38770 36314
rect 38770 36262 38772 36314
rect 38716 36260 38772 36262
rect 15198 35306 15254 35308
rect 15198 35254 15200 35306
rect 15200 35254 15252 35306
rect 15252 35254 15254 35306
rect 15198 35252 15254 35254
rect 15302 35306 15358 35308
rect 15302 35254 15304 35306
rect 15304 35254 15356 35306
rect 15356 35254 15358 35306
rect 15302 35252 15358 35254
rect 15406 35306 15462 35308
rect 15406 35254 15408 35306
rect 15408 35254 15460 35306
rect 15460 35254 15462 35306
rect 15406 35252 15462 35254
rect 15198 33290 15254 33292
rect 15198 33238 15200 33290
rect 15200 33238 15252 33290
rect 15252 33238 15254 33290
rect 15198 33236 15254 33238
rect 15302 33290 15358 33292
rect 15302 33238 15304 33290
rect 15304 33238 15356 33290
rect 15356 33238 15358 33290
rect 15302 33236 15358 33238
rect 15406 33290 15462 33292
rect 15406 33238 15408 33290
rect 15408 33238 15460 33290
rect 15460 33238 15462 33290
rect 15406 33236 15462 33238
rect 24522 35306 24578 35308
rect 24522 35254 24524 35306
rect 24524 35254 24576 35306
rect 24576 35254 24578 35306
rect 24522 35252 24578 35254
rect 24626 35306 24682 35308
rect 24626 35254 24628 35306
rect 24628 35254 24680 35306
rect 24680 35254 24682 35306
rect 24626 35252 24682 35254
rect 24730 35306 24786 35308
rect 24730 35254 24732 35306
rect 24732 35254 24784 35306
rect 24784 35254 24786 35306
rect 24730 35252 24786 35254
rect 33846 35306 33902 35308
rect 33846 35254 33848 35306
rect 33848 35254 33900 35306
rect 33900 35254 33902 35306
rect 33846 35252 33902 35254
rect 33950 35306 34006 35308
rect 33950 35254 33952 35306
rect 33952 35254 34004 35306
rect 34004 35254 34006 35306
rect 33950 35252 34006 35254
rect 34054 35306 34110 35308
rect 34054 35254 34056 35306
rect 34056 35254 34108 35306
rect 34108 35254 34110 35306
rect 34054 35252 34110 35254
rect 19860 34298 19916 34300
rect 19860 34246 19862 34298
rect 19862 34246 19914 34298
rect 19914 34246 19916 34298
rect 19860 34244 19916 34246
rect 19964 34298 20020 34300
rect 19964 34246 19966 34298
rect 19966 34246 20018 34298
rect 20018 34246 20020 34298
rect 19964 34244 20020 34246
rect 20068 34298 20124 34300
rect 20068 34246 20070 34298
rect 20070 34246 20122 34298
rect 20122 34246 20124 34298
rect 20068 34244 20124 34246
rect 29184 34298 29240 34300
rect 29184 34246 29186 34298
rect 29186 34246 29238 34298
rect 29238 34246 29240 34298
rect 29184 34244 29240 34246
rect 29288 34298 29344 34300
rect 29288 34246 29290 34298
rect 29290 34246 29342 34298
rect 29342 34246 29344 34298
rect 29288 34244 29344 34246
rect 29392 34298 29448 34300
rect 29392 34246 29394 34298
rect 29394 34246 29446 34298
rect 29446 34246 29448 34298
rect 29392 34244 29448 34246
rect 38508 34298 38564 34300
rect 38508 34246 38510 34298
rect 38510 34246 38562 34298
rect 38562 34246 38564 34298
rect 38508 34244 38564 34246
rect 38612 34298 38668 34300
rect 38612 34246 38614 34298
rect 38614 34246 38666 34298
rect 38666 34246 38668 34298
rect 38612 34244 38668 34246
rect 38716 34298 38772 34300
rect 38716 34246 38718 34298
rect 38718 34246 38770 34298
rect 38770 34246 38772 34298
rect 38716 34244 38772 34246
rect 24522 33290 24578 33292
rect 24522 33238 24524 33290
rect 24524 33238 24576 33290
rect 24576 33238 24578 33290
rect 24522 33236 24578 33238
rect 24626 33290 24682 33292
rect 24626 33238 24628 33290
rect 24628 33238 24680 33290
rect 24680 33238 24682 33290
rect 24626 33236 24682 33238
rect 24730 33290 24786 33292
rect 24730 33238 24732 33290
rect 24732 33238 24784 33290
rect 24784 33238 24786 33290
rect 24730 33236 24786 33238
rect 33846 33290 33902 33292
rect 33846 33238 33848 33290
rect 33848 33238 33900 33290
rect 33900 33238 33902 33290
rect 33846 33236 33902 33238
rect 33950 33290 34006 33292
rect 33950 33238 33952 33290
rect 33952 33238 34004 33290
rect 34004 33238 34006 33290
rect 33950 33236 34006 33238
rect 34054 33290 34110 33292
rect 34054 33238 34056 33290
rect 34056 33238 34108 33290
rect 34108 33238 34110 33290
rect 34054 33236 34110 33238
rect 19860 32282 19916 32284
rect 19860 32230 19862 32282
rect 19862 32230 19914 32282
rect 19914 32230 19916 32282
rect 19860 32228 19916 32230
rect 19964 32282 20020 32284
rect 19964 32230 19966 32282
rect 19966 32230 20018 32282
rect 20018 32230 20020 32282
rect 19964 32228 20020 32230
rect 20068 32282 20124 32284
rect 20068 32230 20070 32282
rect 20070 32230 20122 32282
rect 20122 32230 20124 32282
rect 20068 32228 20124 32230
rect 29184 32282 29240 32284
rect 29184 32230 29186 32282
rect 29186 32230 29238 32282
rect 29238 32230 29240 32282
rect 29184 32228 29240 32230
rect 29288 32282 29344 32284
rect 29288 32230 29290 32282
rect 29290 32230 29342 32282
rect 29342 32230 29344 32282
rect 29288 32228 29344 32230
rect 29392 32282 29448 32284
rect 29392 32230 29394 32282
rect 29394 32230 29446 32282
rect 29446 32230 29448 32282
rect 29392 32228 29448 32230
rect 38508 32282 38564 32284
rect 38508 32230 38510 32282
rect 38510 32230 38562 32282
rect 38562 32230 38564 32282
rect 38508 32228 38564 32230
rect 38612 32282 38668 32284
rect 38612 32230 38614 32282
rect 38614 32230 38666 32282
rect 38666 32230 38668 32282
rect 38612 32228 38668 32230
rect 38716 32282 38772 32284
rect 38716 32230 38718 32282
rect 38718 32230 38770 32282
rect 38770 32230 38772 32282
rect 38716 32228 38772 32230
rect 5874 31274 5930 31276
rect 5874 31222 5876 31274
rect 5876 31222 5928 31274
rect 5928 31222 5930 31274
rect 5874 31220 5930 31222
rect 5978 31274 6034 31276
rect 5978 31222 5980 31274
rect 5980 31222 6032 31274
rect 6032 31222 6034 31274
rect 5978 31220 6034 31222
rect 6082 31274 6138 31276
rect 6082 31222 6084 31274
rect 6084 31222 6136 31274
rect 6136 31222 6138 31274
rect 6082 31220 6138 31222
rect 15198 31274 15254 31276
rect 15198 31222 15200 31274
rect 15200 31222 15252 31274
rect 15252 31222 15254 31274
rect 15198 31220 15254 31222
rect 15302 31274 15358 31276
rect 15302 31222 15304 31274
rect 15304 31222 15356 31274
rect 15356 31222 15358 31274
rect 15302 31220 15358 31222
rect 15406 31274 15462 31276
rect 15406 31222 15408 31274
rect 15408 31222 15460 31274
rect 15460 31222 15462 31274
rect 15406 31220 15462 31222
rect 24522 31274 24578 31276
rect 24522 31222 24524 31274
rect 24524 31222 24576 31274
rect 24576 31222 24578 31274
rect 24522 31220 24578 31222
rect 24626 31274 24682 31276
rect 24626 31222 24628 31274
rect 24628 31222 24680 31274
rect 24680 31222 24682 31274
rect 24626 31220 24682 31222
rect 24730 31274 24786 31276
rect 24730 31222 24732 31274
rect 24732 31222 24784 31274
rect 24784 31222 24786 31274
rect 24730 31220 24786 31222
rect 33846 31274 33902 31276
rect 33846 31222 33848 31274
rect 33848 31222 33900 31274
rect 33900 31222 33902 31274
rect 33846 31220 33902 31222
rect 33950 31274 34006 31276
rect 33950 31222 33952 31274
rect 33952 31222 34004 31274
rect 34004 31222 34006 31274
rect 33950 31220 34006 31222
rect 34054 31274 34110 31276
rect 34054 31222 34056 31274
rect 34056 31222 34108 31274
rect 34108 31222 34110 31274
rect 34054 31220 34110 31222
rect 10536 30266 10592 30268
rect 10536 30214 10538 30266
rect 10538 30214 10590 30266
rect 10590 30214 10592 30266
rect 10536 30212 10592 30214
rect 10640 30266 10696 30268
rect 10640 30214 10642 30266
rect 10642 30214 10694 30266
rect 10694 30214 10696 30266
rect 10640 30212 10696 30214
rect 10744 30266 10800 30268
rect 10744 30214 10746 30266
rect 10746 30214 10798 30266
rect 10798 30214 10800 30266
rect 10744 30212 10800 30214
rect 19860 30266 19916 30268
rect 19860 30214 19862 30266
rect 19862 30214 19914 30266
rect 19914 30214 19916 30266
rect 19860 30212 19916 30214
rect 19964 30266 20020 30268
rect 19964 30214 19966 30266
rect 19966 30214 20018 30266
rect 20018 30214 20020 30266
rect 19964 30212 20020 30214
rect 20068 30266 20124 30268
rect 20068 30214 20070 30266
rect 20070 30214 20122 30266
rect 20122 30214 20124 30266
rect 20068 30212 20124 30214
rect 29184 30266 29240 30268
rect 29184 30214 29186 30266
rect 29186 30214 29238 30266
rect 29238 30214 29240 30266
rect 29184 30212 29240 30214
rect 29288 30266 29344 30268
rect 29288 30214 29290 30266
rect 29290 30214 29342 30266
rect 29342 30214 29344 30266
rect 29288 30212 29344 30214
rect 29392 30266 29448 30268
rect 29392 30214 29394 30266
rect 29394 30214 29446 30266
rect 29446 30214 29448 30266
rect 29392 30212 29448 30214
rect 38508 30266 38564 30268
rect 38508 30214 38510 30266
rect 38510 30214 38562 30266
rect 38562 30214 38564 30266
rect 38508 30212 38564 30214
rect 38612 30266 38668 30268
rect 38612 30214 38614 30266
rect 38614 30214 38666 30266
rect 38666 30214 38668 30266
rect 38612 30212 38668 30214
rect 38716 30266 38772 30268
rect 38716 30214 38718 30266
rect 38718 30214 38770 30266
rect 38770 30214 38772 30266
rect 38716 30212 38772 30214
rect 5874 29258 5930 29260
rect 5874 29206 5876 29258
rect 5876 29206 5928 29258
rect 5928 29206 5930 29258
rect 5874 29204 5930 29206
rect 5978 29258 6034 29260
rect 5978 29206 5980 29258
rect 5980 29206 6032 29258
rect 6032 29206 6034 29258
rect 5978 29204 6034 29206
rect 6082 29258 6138 29260
rect 6082 29206 6084 29258
rect 6084 29206 6136 29258
rect 6136 29206 6138 29258
rect 6082 29204 6138 29206
rect 15198 29258 15254 29260
rect 15198 29206 15200 29258
rect 15200 29206 15252 29258
rect 15252 29206 15254 29258
rect 15198 29204 15254 29206
rect 15302 29258 15358 29260
rect 15302 29206 15304 29258
rect 15304 29206 15356 29258
rect 15356 29206 15358 29258
rect 15302 29204 15358 29206
rect 15406 29258 15462 29260
rect 15406 29206 15408 29258
rect 15408 29206 15460 29258
rect 15460 29206 15462 29258
rect 15406 29204 15462 29206
rect 24522 29258 24578 29260
rect 24522 29206 24524 29258
rect 24524 29206 24576 29258
rect 24576 29206 24578 29258
rect 24522 29204 24578 29206
rect 24626 29258 24682 29260
rect 24626 29206 24628 29258
rect 24628 29206 24680 29258
rect 24680 29206 24682 29258
rect 24626 29204 24682 29206
rect 24730 29258 24786 29260
rect 24730 29206 24732 29258
rect 24732 29206 24784 29258
rect 24784 29206 24786 29258
rect 24730 29204 24786 29206
rect 33846 29258 33902 29260
rect 33846 29206 33848 29258
rect 33848 29206 33900 29258
rect 33900 29206 33902 29258
rect 33846 29204 33902 29206
rect 33950 29258 34006 29260
rect 33950 29206 33952 29258
rect 33952 29206 34004 29258
rect 34004 29206 34006 29258
rect 33950 29204 34006 29206
rect 34054 29258 34110 29260
rect 34054 29206 34056 29258
rect 34056 29206 34108 29258
rect 34108 29206 34110 29258
rect 34054 29204 34110 29206
rect 10536 28250 10592 28252
rect 10536 28198 10538 28250
rect 10538 28198 10590 28250
rect 10590 28198 10592 28250
rect 10536 28196 10592 28198
rect 10640 28250 10696 28252
rect 10640 28198 10642 28250
rect 10642 28198 10694 28250
rect 10694 28198 10696 28250
rect 10640 28196 10696 28198
rect 10744 28250 10800 28252
rect 10744 28198 10746 28250
rect 10746 28198 10798 28250
rect 10798 28198 10800 28250
rect 10744 28196 10800 28198
rect 19860 28250 19916 28252
rect 19860 28198 19862 28250
rect 19862 28198 19914 28250
rect 19914 28198 19916 28250
rect 19860 28196 19916 28198
rect 19964 28250 20020 28252
rect 19964 28198 19966 28250
rect 19966 28198 20018 28250
rect 20018 28198 20020 28250
rect 19964 28196 20020 28198
rect 20068 28250 20124 28252
rect 20068 28198 20070 28250
rect 20070 28198 20122 28250
rect 20122 28198 20124 28250
rect 20068 28196 20124 28198
rect 29184 28250 29240 28252
rect 29184 28198 29186 28250
rect 29186 28198 29238 28250
rect 29238 28198 29240 28250
rect 29184 28196 29240 28198
rect 29288 28250 29344 28252
rect 29288 28198 29290 28250
rect 29290 28198 29342 28250
rect 29342 28198 29344 28250
rect 29288 28196 29344 28198
rect 29392 28250 29448 28252
rect 29392 28198 29394 28250
rect 29394 28198 29446 28250
rect 29446 28198 29448 28250
rect 29392 28196 29448 28198
rect 38508 28250 38564 28252
rect 38508 28198 38510 28250
rect 38510 28198 38562 28250
rect 38562 28198 38564 28250
rect 38508 28196 38564 28198
rect 38612 28250 38668 28252
rect 38612 28198 38614 28250
rect 38614 28198 38666 28250
rect 38666 28198 38668 28250
rect 38612 28196 38668 28198
rect 38716 28250 38772 28252
rect 38716 28198 38718 28250
rect 38718 28198 38770 28250
rect 38770 28198 38772 28250
rect 38716 28196 38772 28198
rect 5874 27242 5930 27244
rect 5874 27190 5876 27242
rect 5876 27190 5928 27242
rect 5928 27190 5930 27242
rect 5874 27188 5930 27190
rect 5978 27242 6034 27244
rect 5978 27190 5980 27242
rect 5980 27190 6032 27242
rect 6032 27190 6034 27242
rect 5978 27188 6034 27190
rect 6082 27242 6138 27244
rect 6082 27190 6084 27242
rect 6084 27190 6136 27242
rect 6136 27190 6138 27242
rect 6082 27188 6138 27190
rect 15198 27242 15254 27244
rect 15198 27190 15200 27242
rect 15200 27190 15252 27242
rect 15252 27190 15254 27242
rect 15198 27188 15254 27190
rect 15302 27242 15358 27244
rect 15302 27190 15304 27242
rect 15304 27190 15356 27242
rect 15356 27190 15358 27242
rect 15302 27188 15358 27190
rect 15406 27242 15462 27244
rect 15406 27190 15408 27242
rect 15408 27190 15460 27242
rect 15460 27190 15462 27242
rect 15406 27188 15462 27190
rect 24522 27242 24578 27244
rect 24522 27190 24524 27242
rect 24524 27190 24576 27242
rect 24576 27190 24578 27242
rect 24522 27188 24578 27190
rect 24626 27242 24682 27244
rect 24626 27190 24628 27242
rect 24628 27190 24680 27242
rect 24680 27190 24682 27242
rect 24626 27188 24682 27190
rect 24730 27242 24786 27244
rect 24730 27190 24732 27242
rect 24732 27190 24784 27242
rect 24784 27190 24786 27242
rect 24730 27188 24786 27190
rect 33846 27242 33902 27244
rect 33846 27190 33848 27242
rect 33848 27190 33900 27242
rect 33900 27190 33902 27242
rect 33846 27188 33902 27190
rect 33950 27242 34006 27244
rect 33950 27190 33952 27242
rect 33952 27190 34004 27242
rect 34004 27190 34006 27242
rect 33950 27188 34006 27190
rect 34054 27242 34110 27244
rect 34054 27190 34056 27242
rect 34056 27190 34108 27242
rect 34108 27190 34110 27242
rect 34054 27188 34110 27190
rect 10536 26234 10592 26236
rect 10536 26182 10538 26234
rect 10538 26182 10590 26234
rect 10590 26182 10592 26234
rect 10536 26180 10592 26182
rect 10640 26234 10696 26236
rect 10640 26182 10642 26234
rect 10642 26182 10694 26234
rect 10694 26182 10696 26234
rect 10640 26180 10696 26182
rect 10744 26234 10800 26236
rect 10744 26182 10746 26234
rect 10746 26182 10798 26234
rect 10798 26182 10800 26234
rect 10744 26180 10800 26182
rect 19860 26234 19916 26236
rect 19860 26182 19862 26234
rect 19862 26182 19914 26234
rect 19914 26182 19916 26234
rect 19860 26180 19916 26182
rect 19964 26234 20020 26236
rect 19964 26182 19966 26234
rect 19966 26182 20018 26234
rect 20018 26182 20020 26234
rect 19964 26180 20020 26182
rect 20068 26234 20124 26236
rect 20068 26182 20070 26234
rect 20070 26182 20122 26234
rect 20122 26182 20124 26234
rect 20068 26180 20124 26182
rect 29184 26234 29240 26236
rect 29184 26182 29186 26234
rect 29186 26182 29238 26234
rect 29238 26182 29240 26234
rect 29184 26180 29240 26182
rect 29288 26234 29344 26236
rect 29288 26182 29290 26234
rect 29290 26182 29342 26234
rect 29342 26182 29344 26234
rect 29288 26180 29344 26182
rect 29392 26234 29448 26236
rect 29392 26182 29394 26234
rect 29394 26182 29446 26234
rect 29446 26182 29448 26234
rect 29392 26180 29448 26182
rect 38508 26234 38564 26236
rect 38508 26182 38510 26234
rect 38510 26182 38562 26234
rect 38562 26182 38564 26234
rect 38508 26180 38564 26182
rect 38612 26234 38668 26236
rect 38612 26182 38614 26234
rect 38614 26182 38666 26234
rect 38666 26182 38668 26234
rect 38612 26180 38668 26182
rect 38716 26234 38772 26236
rect 38716 26182 38718 26234
rect 38718 26182 38770 26234
rect 38770 26182 38772 26234
rect 38716 26180 38772 26182
rect 34524 25564 34580 25620
rect 5874 25226 5930 25228
rect 5874 25174 5876 25226
rect 5876 25174 5928 25226
rect 5928 25174 5930 25226
rect 5874 25172 5930 25174
rect 5978 25226 6034 25228
rect 5978 25174 5980 25226
rect 5980 25174 6032 25226
rect 6032 25174 6034 25226
rect 5978 25172 6034 25174
rect 6082 25226 6138 25228
rect 6082 25174 6084 25226
rect 6084 25174 6136 25226
rect 6136 25174 6138 25226
rect 6082 25172 6138 25174
rect 15198 25226 15254 25228
rect 15198 25174 15200 25226
rect 15200 25174 15252 25226
rect 15252 25174 15254 25226
rect 15198 25172 15254 25174
rect 15302 25226 15358 25228
rect 15302 25174 15304 25226
rect 15304 25174 15356 25226
rect 15356 25174 15358 25226
rect 15302 25172 15358 25174
rect 15406 25226 15462 25228
rect 15406 25174 15408 25226
rect 15408 25174 15460 25226
rect 15460 25174 15462 25226
rect 15406 25172 15462 25174
rect 24522 25226 24578 25228
rect 24522 25174 24524 25226
rect 24524 25174 24576 25226
rect 24576 25174 24578 25226
rect 24522 25172 24578 25174
rect 24626 25226 24682 25228
rect 24626 25174 24628 25226
rect 24628 25174 24680 25226
rect 24680 25174 24682 25226
rect 24626 25172 24682 25174
rect 24730 25226 24786 25228
rect 24730 25174 24732 25226
rect 24732 25174 24784 25226
rect 24784 25174 24786 25226
rect 24730 25172 24786 25174
rect 33846 25226 33902 25228
rect 33846 25174 33848 25226
rect 33848 25174 33900 25226
rect 33900 25174 33902 25226
rect 33846 25172 33902 25174
rect 33950 25226 34006 25228
rect 33950 25174 33952 25226
rect 33952 25174 34004 25226
rect 34004 25174 34006 25226
rect 33950 25172 34006 25174
rect 34054 25226 34110 25228
rect 34054 25174 34056 25226
rect 34056 25174 34108 25226
rect 34108 25174 34110 25226
rect 34054 25172 34110 25174
rect 4172 24220 4228 24276
rect 4060 23548 4116 23604
rect 10536 24218 10592 24220
rect 10536 24166 10538 24218
rect 10538 24166 10590 24218
rect 10590 24166 10592 24218
rect 10536 24164 10592 24166
rect 10640 24218 10696 24220
rect 10640 24166 10642 24218
rect 10642 24166 10694 24218
rect 10694 24166 10696 24218
rect 10640 24164 10696 24166
rect 10744 24218 10800 24220
rect 10744 24166 10746 24218
rect 10746 24166 10798 24218
rect 10798 24166 10800 24218
rect 10744 24164 10800 24166
rect 19860 24218 19916 24220
rect 19860 24166 19862 24218
rect 19862 24166 19914 24218
rect 19914 24166 19916 24218
rect 19860 24164 19916 24166
rect 19964 24218 20020 24220
rect 19964 24166 19966 24218
rect 19966 24166 20018 24218
rect 20018 24166 20020 24218
rect 19964 24164 20020 24166
rect 20068 24218 20124 24220
rect 20068 24166 20070 24218
rect 20070 24166 20122 24218
rect 20122 24166 20124 24218
rect 20068 24164 20124 24166
rect 29184 24218 29240 24220
rect 29184 24166 29186 24218
rect 29186 24166 29238 24218
rect 29238 24166 29240 24218
rect 29184 24164 29240 24166
rect 29288 24218 29344 24220
rect 29288 24166 29290 24218
rect 29290 24166 29342 24218
rect 29342 24166 29344 24218
rect 29288 24164 29344 24166
rect 29392 24218 29448 24220
rect 29392 24166 29394 24218
rect 29394 24166 29446 24218
rect 29446 24166 29448 24218
rect 29392 24164 29448 24166
rect 5874 23210 5930 23212
rect 5874 23158 5876 23210
rect 5876 23158 5928 23210
rect 5928 23158 5930 23210
rect 5874 23156 5930 23158
rect 5978 23210 6034 23212
rect 5978 23158 5980 23210
rect 5980 23158 6032 23210
rect 6032 23158 6034 23210
rect 5978 23156 6034 23158
rect 6082 23210 6138 23212
rect 6082 23158 6084 23210
rect 6084 23158 6136 23210
rect 6136 23158 6138 23210
rect 6082 23156 6138 23158
rect 15198 23210 15254 23212
rect 15198 23158 15200 23210
rect 15200 23158 15252 23210
rect 15252 23158 15254 23210
rect 15198 23156 15254 23158
rect 15302 23210 15358 23212
rect 15302 23158 15304 23210
rect 15304 23158 15356 23210
rect 15356 23158 15358 23210
rect 15302 23156 15358 23158
rect 15406 23210 15462 23212
rect 15406 23158 15408 23210
rect 15408 23158 15460 23210
rect 15460 23158 15462 23210
rect 15406 23156 15462 23158
rect 24522 23210 24578 23212
rect 24522 23158 24524 23210
rect 24524 23158 24576 23210
rect 24576 23158 24578 23210
rect 24522 23156 24578 23158
rect 24626 23210 24682 23212
rect 24626 23158 24628 23210
rect 24628 23158 24680 23210
rect 24680 23158 24682 23210
rect 24626 23156 24682 23158
rect 24730 23210 24786 23212
rect 24730 23158 24732 23210
rect 24732 23158 24784 23210
rect 24784 23158 24786 23210
rect 24730 23156 24786 23158
rect 33846 23210 33902 23212
rect 33846 23158 33848 23210
rect 33848 23158 33900 23210
rect 33900 23158 33902 23210
rect 33846 23156 33902 23158
rect 33950 23210 34006 23212
rect 33950 23158 33952 23210
rect 33952 23158 34004 23210
rect 34004 23158 34006 23210
rect 33950 23156 34006 23158
rect 34054 23210 34110 23212
rect 34054 23158 34056 23210
rect 34056 23158 34108 23210
rect 34108 23158 34110 23210
rect 34054 23156 34110 23158
rect 4172 22652 4228 22708
rect 4284 22876 4340 22932
rect 13580 22652 13636 22708
rect 10536 22202 10592 22204
rect 10536 22150 10538 22202
rect 10538 22150 10590 22202
rect 10590 22150 10592 22202
rect 10536 22148 10592 22150
rect 10640 22202 10696 22204
rect 10640 22150 10642 22202
rect 10642 22150 10694 22202
rect 10694 22150 10696 22202
rect 10640 22148 10696 22150
rect 10744 22202 10800 22204
rect 10744 22150 10746 22202
rect 10746 22150 10798 22202
rect 10798 22150 10800 22202
rect 10744 22148 10800 22150
rect 5874 21194 5930 21196
rect 5874 21142 5876 21194
rect 5876 21142 5928 21194
rect 5928 21142 5930 21194
rect 5874 21140 5930 21142
rect 5978 21194 6034 21196
rect 5978 21142 5980 21194
rect 5980 21142 6032 21194
rect 6032 21142 6034 21194
rect 5978 21140 6034 21142
rect 6082 21194 6138 21196
rect 6082 21142 6084 21194
rect 6084 21142 6136 21194
rect 6136 21142 6138 21194
rect 6082 21140 6138 21142
rect 4284 20636 4340 20692
rect 4060 20524 4116 20580
rect 12460 20466 12516 20468
rect 12460 20414 12462 20466
rect 12462 20414 12514 20466
rect 12514 20414 12516 20466
rect 12460 20412 12516 20414
rect 4620 20300 4676 20356
rect 4060 18732 4116 18788
rect 4284 18620 4340 18676
rect 4172 18508 4228 18564
rect 4172 17500 4228 17556
rect 12908 20300 12964 20356
rect 10536 20186 10592 20188
rect 10536 20134 10538 20186
rect 10538 20134 10590 20186
rect 10590 20134 10592 20186
rect 10536 20132 10592 20134
rect 10640 20186 10696 20188
rect 10640 20134 10642 20186
rect 10642 20134 10694 20186
rect 10694 20134 10696 20186
rect 10640 20132 10696 20134
rect 10744 20186 10800 20188
rect 10744 20134 10746 20186
rect 10746 20134 10798 20186
rect 10798 20134 10800 20186
rect 10744 20132 10800 20134
rect 19860 22202 19916 22204
rect 19860 22150 19862 22202
rect 19862 22150 19914 22202
rect 19914 22150 19916 22202
rect 19860 22148 19916 22150
rect 19964 22202 20020 22204
rect 19964 22150 19966 22202
rect 19966 22150 20018 22202
rect 20018 22150 20020 22202
rect 19964 22148 20020 22150
rect 20068 22202 20124 22204
rect 20068 22150 20070 22202
rect 20070 22150 20122 22202
rect 20122 22150 20124 22202
rect 20068 22148 20124 22150
rect 29184 22202 29240 22204
rect 29184 22150 29186 22202
rect 29186 22150 29238 22202
rect 29238 22150 29240 22202
rect 29184 22148 29240 22150
rect 29288 22202 29344 22204
rect 29288 22150 29290 22202
rect 29290 22150 29342 22202
rect 29342 22150 29344 22202
rect 29288 22148 29344 22150
rect 29392 22202 29448 22204
rect 29392 22150 29394 22202
rect 29394 22150 29446 22202
rect 29446 22150 29448 22202
rect 29392 22148 29448 22150
rect 17948 21868 18004 21924
rect 15198 21194 15254 21196
rect 15198 21142 15200 21194
rect 15200 21142 15252 21194
rect 15252 21142 15254 21194
rect 15198 21140 15254 21142
rect 15302 21194 15358 21196
rect 15302 21142 15304 21194
rect 15304 21142 15356 21194
rect 15356 21142 15358 21194
rect 15302 21140 15358 21142
rect 15406 21194 15462 21196
rect 15406 21142 15408 21194
rect 15408 21142 15460 21194
rect 15460 21142 15462 21194
rect 15406 21140 15462 21142
rect 13692 20412 13748 20468
rect 13804 20300 13860 20356
rect 14924 20690 14980 20692
rect 14924 20638 14926 20690
rect 14926 20638 14978 20690
rect 14978 20638 14980 20690
rect 14924 20636 14980 20638
rect 5874 19178 5930 19180
rect 5874 19126 5876 19178
rect 5876 19126 5928 19178
rect 5928 19126 5930 19178
rect 5874 19124 5930 19126
rect 5978 19178 6034 19180
rect 5978 19126 5980 19178
rect 5980 19126 6032 19178
rect 6032 19126 6034 19178
rect 5978 19124 6034 19126
rect 6082 19178 6138 19180
rect 6082 19126 6084 19178
rect 6084 19126 6136 19178
rect 6136 19126 6138 19178
rect 6082 19124 6138 19126
rect 13468 19516 13524 19572
rect 11564 18674 11620 18676
rect 11564 18622 11566 18674
rect 11566 18622 11618 18674
rect 11618 18622 11620 18674
rect 11564 18620 11620 18622
rect 11116 18562 11172 18564
rect 11116 18510 11118 18562
rect 11118 18510 11170 18562
rect 11170 18510 11172 18562
rect 11116 18508 11172 18510
rect 12124 18674 12180 18676
rect 12124 18622 12126 18674
rect 12126 18622 12178 18674
rect 12178 18622 12180 18674
rect 12124 18620 12180 18622
rect 12012 18508 12068 18564
rect 4620 18172 4676 18228
rect 10536 18170 10592 18172
rect 10536 18118 10538 18170
rect 10538 18118 10590 18170
rect 10590 18118 10592 18170
rect 10536 18116 10592 18118
rect 10640 18170 10696 18172
rect 10640 18118 10642 18170
rect 10642 18118 10694 18170
rect 10694 18118 10696 18170
rect 10640 18116 10696 18118
rect 10744 18170 10800 18172
rect 10744 18118 10746 18170
rect 10746 18118 10798 18170
rect 10798 18118 10800 18170
rect 10744 18116 10800 18118
rect 17612 20524 17668 20580
rect 16716 19906 16772 19908
rect 16716 19854 16718 19906
rect 16718 19854 16770 19906
rect 16770 19854 16772 19906
rect 16716 19852 16772 19854
rect 31052 21868 31108 21924
rect 22092 21756 22148 21812
rect 19292 21532 19348 21588
rect 18060 20914 18116 20916
rect 18060 20862 18062 20914
rect 18062 20862 18114 20914
rect 18114 20862 18116 20914
rect 18060 20860 18116 20862
rect 18284 20524 18340 20580
rect 14028 19516 14084 19572
rect 15198 19178 15254 19180
rect 15198 19126 15200 19178
rect 15200 19126 15252 19178
rect 15252 19126 15254 19178
rect 15198 19124 15254 19126
rect 15302 19178 15358 19180
rect 15302 19126 15304 19178
rect 15304 19126 15356 19178
rect 15356 19126 15358 19178
rect 15302 19124 15358 19126
rect 15406 19178 15462 19180
rect 15406 19126 15408 19178
rect 15408 19126 15460 19178
rect 15460 19126 15462 19178
rect 15406 19124 15462 19126
rect 15932 18844 15988 18900
rect 16268 18786 16324 18788
rect 16268 18734 16270 18786
rect 16270 18734 16322 18786
rect 16322 18734 16324 18786
rect 16268 18732 16324 18734
rect 20860 20524 20916 20580
rect 20748 20354 20804 20356
rect 20748 20302 20750 20354
rect 20750 20302 20802 20354
rect 20802 20302 20804 20354
rect 20748 20300 20804 20302
rect 18844 19852 18900 19908
rect 19860 20186 19916 20188
rect 19860 20134 19862 20186
rect 19862 20134 19914 20186
rect 19914 20134 19916 20186
rect 19860 20132 19916 20134
rect 19964 20186 20020 20188
rect 19964 20134 19966 20186
rect 19966 20134 20018 20186
rect 20018 20134 20020 20186
rect 19964 20132 20020 20134
rect 20068 20186 20124 20188
rect 20068 20134 20070 20186
rect 20070 20134 20122 20186
rect 20122 20134 20124 20186
rect 20068 20132 20124 20134
rect 16828 18844 16884 18900
rect 16940 18732 16996 18788
rect 27356 21532 27412 21588
rect 24522 21194 24578 21196
rect 24522 21142 24524 21194
rect 24524 21142 24576 21194
rect 24576 21142 24578 21194
rect 24522 21140 24578 21142
rect 24626 21194 24682 21196
rect 24626 21142 24628 21194
rect 24628 21142 24680 21194
rect 24680 21142 24682 21194
rect 24626 21140 24682 21142
rect 24730 21194 24786 21196
rect 24730 21142 24732 21194
rect 24732 21142 24784 21194
rect 24784 21142 24786 21194
rect 24730 21140 24786 21142
rect 25116 20860 25172 20916
rect 21980 20412 22036 20468
rect 21532 20300 21588 20356
rect 22316 20690 22372 20692
rect 22316 20638 22318 20690
rect 22318 20638 22370 20690
rect 22370 20638 22372 20690
rect 22316 20636 22372 20638
rect 23436 20578 23492 20580
rect 23436 20526 23438 20578
rect 23438 20526 23490 20578
rect 23490 20526 23492 20578
rect 23436 20524 23492 20526
rect 24332 20578 24388 20580
rect 24332 20526 24334 20578
rect 24334 20526 24386 20578
rect 24386 20526 24388 20578
rect 24332 20524 24388 20526
rect 22876 20466 22932 20468
rect 22876 20414 22878 20466
rect 22878 20414 22930 20466
rect 22930 20414 22932 20466
rect 22876 20412 22932 20414
rect 23660 20188 23716 20244
rect 22876 19852 22932 19908
rect 25116 20188 25172 20244
rect 24332 19516 24388 19572
rect 19860 18170 19916 18172
rect 19860 18118 19862 18170
rect 19862 18118 19914 18170
rect 19914 18118 19916 18170
rect 19860 18116 19916 18118
rect 19964 18170 20020 18172
rect 19964 18118 19966 18170
rect 19966 18118 20018 18170
rect 20018 18118 20020 18170
rect 19964 18116 20020 18118
rect 20068 18170 20124 18172
rect 20068 18118 20070 18170
rect 20070 18118 20122 18170
rect 20122 18118 20124 18170
rect 20068 18116 20124 18118
rect 24522 19178 24578 19180
rect 24522 19126 24524 19178
rect 24524 19126 24576 19178
rect 24576 19126 24578 19178
rect 24522 19124 24578 19126
rect 24626 19178 24682 19180
rect 24626 19126 24628 19178
rect 24628 19126 24680 19178
rect 24680 19126 24682 19178
rect 24626 19124 24682 19126
rect 24730 19178 24786 19180
rect 24730 19126 24732 19178
rect 24732 19126 24784 19178
rect 24784 19126 24786 19178
rect 24730 19124 24786 19126
rect 23436 17500 23492 17556
rect 5874 17162 5930 17164
rect 5874 17110 5876 17162
rect 5876 17110 5928 17162
rect 5928 17110 5930 17162
rect 5874 17108 5930 17110
rect 5978 17162 6034 17164
rect 5978 17110 5980 17162
rect 5980 17110 6032 17162
rect 6032 17110 6034 17162
rect 5978 17108 6034 17110
rect 6082 17162 6138 17164
rect 6082 17110 6084 17162
rect 6084 17110 6136 17162
rect 6136 17110 6138 17162
rect 6082 17108 6138 17110
rect 15198 17162 15254 17164
rect 15198 17110 15200 17162
rect 15200 17110 15252 17162
rect 15252 17110 15254 17162
rect 15198 17108 15254 17110
rect 15302 17162 15358 17164
rect 15302 17110 15304 17162
rect 15304 17110 15356 17162
rect 15356 17110 15358 17162
rect 15302 17108 15358 17110
rect 15406 17162 15462 17164
rect 15406 17110 15408 17162
rect 15408 17110 15460 17162
rect 15460 17110 15462 17162
rect 15406 17108 15462 17110
rect 24522 17162 24578 17164
rect 24522 17110 24524 17162
rect 24524 17110 24576 17162
rect 24576 17110 24578 17162
rect 24522 17108 24578 17110
rect 24626 17162 24682 17164
rect 24626 17110 24628 17162
rect 24628 17110 24680 17162
rect 24680 17110 24682 17162
rect 24626 17108 24682 17110
rect 24730 17162 24786 17164
rect 24730 17110 24732 17162
rect 24732 17110 24784 17162
rect 24784 17110 24786 17162
rect 24730 17108 24786 17110
rect 4284 16828 4340 16884
rect 4060 16156 4116 16212
rect 10536 16154 10592 16156
rect 10536 16102 10538 16154
rect 10538 16102 10590 16154
rect 10590 16102 10592 16154
rect 10536 16100 10592 16102
rect 10640 16154 10696 16156
rect 10640 16102 10642 16154
rect 10642 16102 10694 16154
rect 10694 16102 10696 16154
rect 10640 16100 10696 16102
rect 10744 16154 10800 16156
rect 10744 16102 10746 16154
rect 10746 16102 10798 16154
rect 10798 16102 10800 16154
rect 10744 16100 10800 16102
rect 19860 16154 19916 16156
rect 19860 16102 19862 16154
rect 19862 16102 19914 16154
rect 19914 16102 19916 16154
rect 19860 16100 19916 16102
rect 19964 16154 20020 16156
rect 19964 16102 19966 16154
rect 19966 16102 20018 16154
rect 20018 16102 20020 16154
rect 19964 16100 20020 16102
rect 20068 16154 20124 16156
rect 20068 16102 20070 16154
rect 20070 16102 20122 16154
rect 20122 16102 20124 16154
rect 20068 16100 20124 16102
rect 26460 20188 26516 20244
rect 27244 20188 27300 20244
rect 25340 19906 25396 19908
rect 25340 19854 25342 19906
rect 25342 19854 25394 19906
rect 25394 19854 25396 19906
rect 25340 19852 25396 19854
rect 25788 19570 25844 19572
rect 25788 19518 25790 19570
rect 25790 19518 25842 19570
rect 25842 19518 25844 19570
rect 25788 19516 25844 19518
rect 26348 19570 26404 19572
rect 26348 19518 26350 19570
rect 26350 19518 26402 19570
rect 26402 19518 26404 19570
rect 26348 19516 26404 19518
rect 26012 18786 26068 18788
rect 26012 18734 26014 18786
rect 26014 18734 26066 18786
rect 26066 18734 26068 18786
rect 26012 18732 26068 18734
rect 33846 21194 33902 21196
rect 33846 21142 33848 21194
rect 33848 21142 33900 21194
rect 33900 21142 33902 21194
rect 33846 21140 33902 21142
rect 33950 21194 34006 21196
rect 33950 21142 33952 21194
rect 33952 21142 34004 21194
rect 34004 21142 34006 21194
rect 33950 21140 34006 21142
rect 34054 21194 34110 21196
rect 34054 21142 34056 21194
rect 34056 21142 34108 21194
rect 34108 21142 34110 21194
rect 34054 21140 34110 21142
rect 28140 20748 28196 20804
rect 28140 20188 28196 20244
rect 28924 20300 28980 20356
rect 29596 20300 29652 20356
rect 29184 20186 29240 20188
rect 29184 20134 29186 20186
rect 29186 20134 29238 20186
rect 29238 20134 29240 20186
rect 29184 20132 29240 20134
rect 29288 20186 29344 20188
rect 29288 20134 29290 20186
rect 29290 20134 29342 20186
rect 29342 20134 29344 20186
rect 29288 20132 29344 20134
rect 29392 20186 29448 20188
rect 29392 20134 29394 20186
rect 29394 20134 29446 20186
rect 29446 20134 29448 20186
rect 29392 20132 29448 20134
rect 30716 20412 30772 20468
rect 34300 20524 34356 20580
rect 30940 19964 30996 20020
rect 30044 19516 30100 19572
rect 30044 18844 30100 18900
rect 30716 19516 30772 19572
rect 29708 18674 29764 18676
rect 29708 18622 29710 18674
rect 29710 18622 29762 18674
rect 29762 18622 29764 18674
rect 29708 18620 29764 18622
rect 31948 19964 32004 20020
rect 31500 19570 31556 19572
rect 31500 19518 31502 19570
rect 31502 19518 31554 19570
rect 31554 19518 31556 19570
rect 31500 19516 31556 19518
rect 33846 19178 33902 19180
rect 33846 19126 33848 19178
rect 33848 19126 33900 19178
rect 33900 19126 33902 19178
rect 33846 19124 33902 19126
rect 33950 19178 34006 19180
rect 33950 19126 33952 19178
rect 33952 19126 34004 19178
rect 34004 19126 34006 19178
rect 33950 19124 34006 19126
rect 34054 19178 34110 19180
rect 34054 19126 34056 19178
rect 34056 19126 34108 19178
rect 34108 19126 34110 19178
rect 34054 19124 34110 19126
rect 30604 18674 30660 18676
rect 30604 18622 30606 18674
rect 30606 18622 30658 18674
rect 30658 18622 30660 18674
rect 30604 18620 30660 18622
rect 26908 18508 26964 18564
rect 27916 18562 27972 18564
rect 27916 18510 27918 18562
rect 27918 18510 27970 18562
rect 27970 18510 27972 18562
rect 27916 18508 27972 18510
rect 28588 18562 28644 18564
rect 28588 18510 28590 18562
rect 28590 18510 28642 18562
rect 28642 18510 28644 18562
rect 28588 18508 28644 18510
rect 30044 18450 30100 18452
rect 30044 18398 30046 18450
rect 30046 18398 30098 18450
rect 30098 18398 30100 18450
rect 30044 18396 30100 18398
rect 29184 18170 29240 18172
rect 29184 18118 29186 18170
rect 29186 18118 29238 18170
rect 29238 18118 29240 18170
rect 29184 18116 29240 18118
rect 29288 18170 29344 18172
rect 29288 18118 29290 18170
rect 29290 18118 29342 18170
rect 29342 18118 29344 18170
rect 29288 18116 29344 18118
rect 29392 18170 29448 18172
rect 29392 18118 29394 18170
rect 29394 18118 29446 18170
rect 29446 18118 29448 18170
rect 29392 18116 29448 18118
rect 26012 17554 26068 17556
rect 26012 17502 26014 17554
rect 26014 17502 26066 17554
rect 26066 17502 26068 17554
rect 26012 17500 26068 17502
rect 33846 17162 33902 17164
rect 33846 17110 33848 17162
rect 33848 17110 33900 17162
rect 33900 17110 33902 17162
rect 33846 17108 33902 17110
rect 33950 17162 34006 17164
rect 33950 17110 33952 17162
rect 33952 17110 34004 17162
rect 34004 17110 34006 17162
rect 33950 17108 34006 17110
rect 34054 17162 34110 17164
rect 34054 17110 34056 17162
rect 34056 17110 34108 17162
rect 34108 17110 34110 17162
rect 34054 17108 34110 17110
rect 29184 16154 29240 16156
rect 29184 16102 29186 16154
rect 29186 16102 29238 16154
rect 29238 16102 29240 16154
rect 29184 16100 29240 16102
rect 29288 16154 29344 16156
rect 29288 16102 29290 16154
rect 29290 16102 29342 16154
rect 29342 16102 29344 16154
rect 29288 16100 29344 16102
rect 29392 16154 29448 16156
rect 29392 16102 29394 16154
rect 29394 16102 29446 16154
rect 29446 16102 29448 16154
rect 29392 16100 29448 16102
rect 24892 15484 24948 15540
rect 5874 15146 5930 15148
rect 5874 15094 5876 15146
rect 5876 15094 5928 15146
rect 5928 15094 5930 15146
rect 5874 15092 5930 15094
rect 5978 15146 6034 15148
rect 5978 15094 5980 15146
rect 5980 15094 6032 15146
rect 6032 15094 6034 15146
rect 5978 15092 6034 15094
rect 6082 15146 6138 15148
rect 6082 15094 6084 15146
rect 6084 15094 6136 15146
rect 6136 15094 6138 15146
rect 6082 15092 6138 15094
rect 15198 15146 15254 15148
rect 15198 15094 15200 15146
rect 15200 15094 15252 15146
rect 15252 15094 15254 15146
rect 15198 15092 15254 15094
rect 15302 15146 15358 15148
rect 15302 15094 15304 15146
rect 15304 15094 15356 15146
rect 15356 15094 15358 15146
rect 15302 15092 15358 15094
rect 15406 15146 15462 15148
rect 15406 15094 15408 15146
rect 15408 15094 15460 15146
rect 15460 15094 15462 15146
rect 15406 15092 15462 15094
rect 24522 15146 24578 15148
rect 24522 15094 24524 15146
rect 24524 15094 24576 15146
rect 24576 15094 24578 15146
rect 24522 15092 24578 15094
rect 24626 15146 24682 15148
rect 24626 15094 24628 15146
rect 24628 15094 24680 15146
rect 24680 15094 24682 15146
rect 24626 15092 24682 15094
rect 24730 15146 24786 15148
rect 24730 15094 24732 15146
rect 24732 15094 24784 15146
rect 24784 15094 24786 15146
rect 24730 15092 24786 15094
rect 33846 15146 33902 15148
rect 33846 15094 33848 15146
rect 33848 15094 33900 15146
rect 33900 15094 33902 15146
rect 33846 15092 33902 15094
rect 33950 15146 34006 15148
rect 33950 15094 33952 15146
rect 33952 15094 34004 15146
rect 34004 15094 34006 15146
rect 33950 15092 34006 15094
rect 34054 15146 34110 15148
rect 34054 15094 34056 15146
rect 34056 15094 34108 15146
rect 34108 15094 34110 15146
rect 34054 15092 34110 15094
rect 34748 24892 34804 24948
rect 38508 24218 38564 24220
rect 38508 24166 38510 24218
rect 38510 24166 38562 24218
rect 38562 24166 38564 24218
rect 38508 24164 38564 24166
rect 38612 24218 38668 24220
rect 38612 24166 38614 24218
rect 38614 24166 38666 24218
rect 38666 24166 38668 24218
rect 38612 24164 38668 24166
rect 38716 24218 38772 24220
rect 38716 24166 38718 24218
rect 38718 24166 38770 24218
rect 38770 24166 38772 24218
rect 38716 24164 38772 24166
rect 35084 23996 35140 24052
rect 34972 22876 35028 22932
rect 34748 20748 34804 20804
rect 34860 21980 34916 22036
rect 35196 23548 35252 23604
rect 38508 22202 38564 22204
rect 38508 22150 38510 22202
rect 38510 22150 38562 22202
rect 38562 22150 38564 22202
rect 38508 22148 38564 22150
rect 38612 22202 38668 22204
rect 38612 22150 38614 22202
rect 38614 22150 38666 22202
rect 38666 22150 38668 22202
rect 38612 22148 38668 22150
rect 38716 22202 38772 22204
rect 38716 22150 38718 22202
rect 38718 22150 38770 22202
rect 38770 22150 38772 22202
rect 38716 22148 38772 22150
rect 35196 21868 35252 21924
rect 35084 21756 35140 21812
rect 34972 20860 35028 20916
rect 34860 20636 34916 20692
rect 34636 20300 34692 20356
rect 38508 20186 38564 20188
rect 38508 20134 38510 20186
rect 38510 20134 38562 20186
rect 38562 20134 38564 20186
rect 38508 20132 38564 20134
rect 38612 20186 38668 20188
rect 38612 20134 38614 20186
rect 38614 20134 38666 20186
rect 38666 20134 38668 20186
rect 38612 20132 38668 20134
rect 38716 20186 38772 20188
rect 38716 20134 38718 20186
rect 38718 20134 38770 20186
rect 38770 20134 38772 20186
rect 38716 20132 38772 20134
rect 34636 19964 34692 20020
rect 34524 19852 34580 19908
rect 35084 18844 35140 18900
rect 35196 18732 35252 18788
rect 38508 18170 38564 18172
rect 38508 18118 38510 18170
rect 38510 18118 38562 18170
rect 38562 18118 38564 18170
rect 38508 18116 38564 18118
rect 38612 18170 38668 18172
rect 38612 18118 38614 18170
rect 38614 18118 38666 18170
rect 38666 18118 38668 18170
rect 38612 18116 38668 18118
rect 38716 18170 38772 18172
rect 38716 18118 38718 18170
rect 38718 18118 38770 18170
rect 38770 18118 38772 18170
rect 38716 18116 38772 18118
rect 35196 16828 35252 16884
rect 35084 16268 35140 16324
rect 38508 16154 38564 16156
rect 38508 16102 38510 16154
rect 38510 16102 38562 16154
rect 38562 16102 38564 16154
rect 38508 16100 38564 16102
rect 38612 16154 38668 16156
rect 38612 16102 38614 16154
rect 38614 16102 38666 16154
rect 38666 16102 38668 16154
rect 38612 16100 38668 16102
rect 38716 16154 38772 16156
rect 38716 16102 38718 16154
rect 38718 16102 38770 16154
rect 38770 16102 38772 16154
rect 38716 16100 38772 16102
rect 34300 14812 34356 14868
rect 10536 14138 10592 14140
rect 10536 14086 10538 14138
rect 10538 14086 10590 14138
rect 10590 14086 10592 14138
rect 10536 14084 10592 14086
rect 10640 14138 10696 14140
rect 10640 14086 10642 14138
rect 10642 14086 10694 14138
rect 10694 14086 10696 14138
rect 10640 14084 10696 14086
rect 10744 14138 10800 14140
rect 10744 14086 10746 14138
rect 10746 14086 10798 14138
rect 10798 14086 10800 14138
rect 10744 14084 10800 14086
rect 19860 14138 19916 14140
rect 19860 14086 19862 14138
rect 19862 14086 19914 14138
rect 19914 14086 19916 14138
rect 19860 14084 19916 14086
rect 19964 14138 20020 14140
rect 19964 14086 19966 14138
rect 19966 14086 20018 14138
rect 20018 14086 20020 14138
rect 19964 14084 20020 14086
rect 20068 14138 20124 14140
rect 20068 14086 20070 14138
rect 20070 14086 20122 14138
rect 20122 14086 20124 14138
rect 20068 14084 20124 14086
rect 29184 14138 29240 14140
rect 29184 14086 29186 14138
rect 29186 14086 29238 14138
rect 29238 14086 29240 14138
rect 29184 14084 29240 14086
rect 29288 14138 29344 14140
rect 29288 14086 29290 14138
rect 29290 14086 29342 14138
rect 29342 14086 29344 14138
rect 29288 14084 29344 14086
rect 29392 14138 29448 14140
rect 29392 14086 29394 14138
rect 29394 14086 29446 14138
rect 29446 14086 29448 14138
rect 29392 14084 29448 14086
rect 38508 14138 38564 14140
rect 38508 14086 38510 14138
rect 38510 14086 38562 14138
rect 38562 14086 38564 14138
rect 38508 14084 38564 14086
rect 38612 14138 38668 14140
rect 38612 14086 38614 14138
rect 38614 14086 38666 14138
rect 38666 14086 38668 14138
rect 38612 14084 38668 14086
rect 38716 14138 38772 14140
rect 38716 14086 38718 14138
rect 38718 14086 38770 14138
rect 38770 14086 38772 14138
rect 38716 14084 38772 14086
rect 5874 13130 5930 13132
rect 5874 13078 5876 13130
rect 5876 13078 5928 13130
rect 5928 13078 5930 13130
rect 5874 13076 5930 13078
rect 5978 13130 6034 13132
rect 5978 13078 5980 13130
rect 5980 13078 6032 13130
rect 6032 13078 6034 13130
rect 5978 13076 6034 13078
rect 6082 13130 6138 13132
rect 6082 13078 6084 13130
rect 6084 13078 6136 13130
rect 6136 13078 6138 13130
rect 6082 13076 6138 13078
rect 15198 13130 15254 13132
rect 15198 13078 15200 13130
rect 15200 13078 15252 13130
rect 15252 13078 15254 13130
rect 15198 13076 15254 13078
rect 15302 13130 15358 13132
rect 15302 13078 15304 13130
rect 15304 13078 15356 13130
rect 15356 13078 15358 13130
rect 15302 13076 15358 13078
rect 15406 13130 15462 13132
rect 15406 13078 15408 13130
rect 15408 13078 15460 13130
rect 15460 13078 15462 13130
rect 15406 13076 15462 13078
rect 24522 13130 24578 13132
rect 24522 13078 24524 13130
rect 24524 13078 24576 13130
rect 24576 13078 24578 13130
rect 24522 13076 24578 13078
rect 24626 13130 24682 13132
rect 24626 13078 24628 13130
rect 24628 13078 24680 13130
rect 24680 13078 24682 13130
rect 24626 13076 24682 13078
rect 24730 13130 24786 13132
rect 24730 13078 24732 13130
rect 24732 13078 24784 13130
rect 24784 13078 24786 13130
rect 24730 13076 24786 13078
rect 33846 13130 33902 13132
rect 33846 13078 33848 13130
rect 33848 13078 33900 13130
rect 33900 13078 33902 13130
rect 33846 13076 33902 13078
rect 33950 13130 34006 13132
rect 33950 13078 33952 13130
rect 33952 13078 34004 13130
rect 34004 13078 34006 13130
rect 33950 13076 34006 13078
rect 34054 13130 34110 13132
rect 34054 13078 34056 13130
rect 34056 13078 34108 13130
rect 34108 13078 34110 13130
rect 34054 13076 34110 13078
rect 10536 12122 10592 12124
rect 10536 12070 10538 12122
rect 10538 12070 10590 12122
rect 10590 12070 10592 12122
rect 10536 12068 10592 12070
rect 10640 12122 10696 12124
rect 10640 12070 10642 12122
rect 10642 12070 10694 12122
rect 10694 12070 10696 12122
rect 10640 12068 10696 12070
rect 10744 12122 10800 12124
rect 10744 12070 10746 12122
rect 10746 12070 10798 12122
rect 10798 12070 10800 12122
rect 10744 12068 10800 12070
rect 19860 12122 19916 12124
rect 19860 12070 19862 12122
rect 19862 12070 19914 12122
rect 19914 12070 19916 12122
rect 19860 12068 19916 12070
rect 19964 12122 20020 12124
rect 19964 12070 19966 12122
rect 19966 12070 20018 12122
rect 20018 12070 20020 12122
rect 19964 12068 20020 12070
rect 20068 12122 20124 12124
rect 20068 12070 20070 12122
rect 20070 12070 20122 12122
rect 20122 12070 20124 12122
rect 20068 12068 20124 12070
rect 29184 12122 29240 12124
rect 29184 12070 29186 12122
rect 29186 12070 29238 12122
rect 29238 12070 29240 12122
rect 29184 12068 29240 12070
rect 29288 12122 29344 12124
rect 29288 12070 29290 12122
rect 29290 12070 29342 12122
rect 29342 12070 29344 12122
rect 29288 12068 29344 12070
rect 29392 12122 29448 12124
rect 29392 12070 29394 12122
rect 29394 12070 29446 12122
rect 29446 12070 29448 12122
rect 29392 12068 29448 12070
rect 38508 12122 38564 12124
rect 38508 12070 38510 12122
rect 38510 12070 38562 12122
rect 38562 12070 38564 12122
rect 38508 12068 38564 12070
rect 38612 12122 38668 12124
rect 38612 12070 38614 12122
rect 38614 12070 38666 12122
rect 38666 12070 38668 12122
rect 38612 12068 38668 12070
rect 38716 12122 38772 12124
rect 38716 12070 38718 12122
rect 38718 12070 38770 12122
rect 38770 12070 38772 12122
rect 38716 12068 38772 12070
rect 5874 11114 5930 11116
rect 5874 11062 5876 11114
rect 5876 11062 5928 11114
rect 5928 11062 5930 11114
rect 5874 11060 5930 11062
rect 5978 11114 6034 11116
rect 5978 11062 5980 11114
rect 5980 11062 6032 11114
rect 6032 11062 6034 11114
rect 5978 11060 6034 11062
rect 6082 11114 6138 11116
rect 6082 11062 6084 11114
rect 6084 11062 6136 11114
rect 6136 11062 6138 11114
rect 6082 11060 6138 11062
rect 15198 11114 15254 11116
rect 15198 11062 15200 11114
rect 15200 11062 15252 11114
rect 15252 11062 15254 11114
rect 15198 11060 15254 11062
rect 15302 11114 15358 11116
rect 15302 11062 15304 11114
rect 15304 11062 15356 11114
rect 15356 11062 15358 11114
rect 15302 11060 15358 11062
rect 15406 11114 15462 11116
rect 15406 11062 15408 11114
rect 15408 11062 15460 11114
rect 15460 11062 15462 11114
rect 15406 11060 15462 11062
rect 24522 11114 24578 11116
rect 24522 11062 24524 11114
rect 24524 11062 24576 11114
rect 24576 11062 24578 11114
rect 24522 11060 24578 11062
rect 24626 11114 24682 11116
rect 24626 11062 24628 11114
rect 24628 11062 24680 11114
rect 24680 11062 24682 11114
rect 24626 11060 24682 11062
rect 24730 11114 24786 11116
rect 24730 11062 24732 11114
rect 24732 11062 24784 11114
rect 24784 11062 24786 11114
rect 24730 11060 24786 11062
rect 33846 11114 33902 11116
rect 33846 11062 33848 11114
rect 33848 11062 33900 11114
rect 33900 11062 33902 11114
rect 33846 11060 33902 11062
rect 33950 11114 34006 11116
rect 33950 11062 33952 11114
rect 33952 11062 34004 11114
rect 34004 11062 34006 11114
rect 33950 11060 34006 11062
rect 34054 11114 34110 11116
rect 34054 11062 34056 11114
rect 34056 11062 34108 11114
rect 34108 11062 34110 11114
rect 34054 11060 34110 11062
rect 10536 10106 10592 10108
rect 10536 10054 10538 10106
rect 10538 10054 10590 10106
rect 10590 10054 10592 10106
rect 10536 10052 10592 10054
rect 10640 10106 10696 10108
rect 10640 10054 10642 10106
rect 10642 10054 10694 10106
rect 10694 10054 10696 10106
rect 10640 10052 10696 10054
rect 10744 10106 10800 10108
rect 10744 10054 10746 10106
rect 10746 10054 10798 10106
rect 10798 10054 10800 10106
rect 10744 10052 10800 10054
rect 19860 10106 19916 10108
rect 19860 10054 19862 10106
rect 19862 10054 19914 10106
rect 19914 10054 19916 10106
rect 19860 10052 19916 10054
rect 19964 10106 20020 10108
rect 19964 10054 19966 10106
rect 19966 10054 20018 10106
rect 20018 10054 20020 10106
rect 19964 10052 20020 10054
rect 20068 10106 20124 10108
rect 20068 10054 20070 10106
rect 20070 10054 20122 10106
rect 20122 10054 20124 10106
rect 20068 10052 20124 10054
rect 29184 10106 29240 10108
rect 29184 10054 29186 10106
rect 29186 10054 29238 10106
rect 29238 10054 29240 10106
rect 29184 10052 29240 10054
rect 29288 10106 29344 10108
rect 29288 10054 29290 10106
rect 29290 10054 29342 10106
rect 29342 10054 29344 10106
rect 29288 10052 29344 10054
rect 29392 10106 29448 10108
rect 29392 10054 29394 10106
rect 29394 10054 29446 10106
rect 29446 10054 29448 10106
rect 29392 10052 29448 10054
rect 38508 10106 38564 10108
rect 38508 10054 38510 10106
rect 38510 10054 38562 10106
rect 38562 10054 38564 10106
rect 38508 10052 38564 10054
rect 38612 10106 38668 10108
rect 38612 10054 38614 10106
rect 38614 10054 38666 10106
rect 38666 10054 38668 10106
rect 38612 10052 38668 10054
rect 38716 10106 38772 10108
rect 38716 10054 38718 10106
rect 38718 10054 38770 10106
rect 38770 10054 38772 10106
rect 38716 10052 38772 10054
rect 5874 9098 5930 9100
rect 5874 9046 5876 9098
rect 5876 9046 5928 9098
rect 5928 9046 5930 9098
rect 5874 9044 5930 9046
rect 5978 9098 6034 9100
rect 5978 9046 5980 9098
rect 5980 9046 6032 9098
rect 6032 9046 6034 9098
rect 5978 9044 6034 9046
rect 6082 9098 6138 9100
rect 6082 9046 6084 9098
rect 6084 9046 6136 9098
rect 6136 9046 6138 9098
rect 6082 9044 6138 9046
rect 15198 9098 15254 9100
rect 15198 9046 15200 9098
rect 15200 9046 15252 9098
rect 15252 9046 15254 9098
rect 15198 9044 15254 9046
rect 15302 9098 15358 9100
rect 15302 9046 15304 9098
rect 15304 9046 15356 9098
rect 15356 9046 15358 9098
rect 15302 9044 15358 9046
rect 15406 9098 15462 9100
rect 15406 9046 15408 9098
rect 15408 9046 15460 9098
rect 15460 9046 15462 9098
rect 15406 9044 15462 9046
rect 24522 9098 24578 9100
rect 24522 9046 24524 9098
rect 24524 9046 24576 9098
rect 24576 9046 24578 9098
rect 24522 9044 24578 9046
rect 24626 9098 24682 9100
rect 24626 9046 24628 9098
rect 24628 9046 24680 9098
rect 24680 9046 24682 9098
rect 24626 9044 24682 9046
rect 24730 9098 24786 9100
rect 24730 9046 24732 9098
rect 24732 9046 24784 9098
rect 24784 9046 24786 9098
rect 24730 9044 24786 9046
rect 33846 9098 33902 9100
rect 33846 9046 33848 9098
rect 33848 9046 33900 9098
rect 33900 9046 33902 9098
rect 33846 9044 33902 9046
rect 33950 9098 34006 9100
rect 33950 9046 33952 9098
rect 33952 9046 34004 9098
rect 34004 9046 34006 9098
rect 33950 9044 34006 9046
rect 34054 9098 34110 9100
rect 34054 9046 34056 9098
rect 34056 9046 34108 9098
rect 34108 9046 34110 9098
rect 34054 9044 34110 9046
rect 10536 8090 10592 8092
rect 10536 8038 10538 8090
rect 10538 8038 10590 8090
rect 10590 8038 10592 8090
rect 10536 8036 10592 8038
rect 10640 8090 10696 8092
rect 10640 8038 10642 8090
rect 10642 8038 10694 8090
rect 10694 8038 10696 8090
rect 10640 8036 10696 8038
rect 10744 8090 10800 8092
rect 10744 8038 10746 8090
rect 10746 8038 10798 8090
rect 10798 8038 10800 8090
rect 10744 8036 10800 8038
rect 19860 8090 19916 8092
rect 19860 8038 19862 8090
rect 19862 8038 19914 8090
rect 19914 8038 19916 8090
rect 19860 8036 19916 8038
rect 19964 8090 20020 8092
rect 19964 8038 19966 8090
rect 19966 8038 20018 8090
rect 20018 8038 20020 8090
rect 19964 8036 20020 8038
rect 20068 8090 20124 8092
rect 20068 8038 20070 8090
rect 20070 8038 20122 8090
rect 20122 8038 20124 8090
rect 20068 8036 20124 8038
rect 29184 8090 29240 8092
rect 29184 8038 29186 8090
rect 29186 8038 29238 8090
rect 29238 8038 29240 8090
rect 29184 8036 29240 8038
rect 29288 8090 29344 8092
rect 29288 8038 29290 8090
rect 29290 8038 29342 8090
rect 29342 8038 29344 8090
rect 29288 8036 29344 8038
rect 29392 8090 29448 8092
rect 29392 8038 29394 8090
rect 29394 8038 29446 8090
rect 29446 8038 29448 8090
rect 29392 8036 29448 8038
rect 38508 8090 38564 8092
rect 38508 8038 38510 8090
rect 38510 8038 38562 8090
rect 38562 8038 38564 8090
rect 38508 8036 38564 8038
rect 38612 8090 38668 8092
rect 38612 8038 38614 8090
rect 38614 8038 38666 8090
rect 38666 8038 38668 8090
rect 38612 8036 38668 8038
rect 38716 8090 38772 8092
rect 38716 8038 38718 8090
rect 38718 8038 38770 8090
rect 38770 8038 38772 8090
rect 38716 8036 38772 8038
rect 5874 7082 5930 7084
rect 5874 7030 5876 7082
rect 5876 7030 5928 7082
rect 5928 7030 5930 7082
rect 5874 7028 5930 7030
rect 5978 7082 6034 7084
rect 5978 7030 5980 7082
rect 5980 7030 6032 7082
rect 6032 7030 6034 7082
rect 5978 7028 6034 7030
rect 6082 7082 6138 7084
rect 6082 7030 6084 7082
rect 6084 7030 6136 7082
rect 6136 7030 6138 7082
rect 6082 7028 6138 7030
rect 15198 7082 15254 7084
rect 15198 7030 15200 7082
rect 15200 7030 15252 7082
rect 15252 7030 15254 7082
rect 15198 7028 15254 7030
rect 15302 7082 15358 7084
rect 15302 7030 15304 7082
rect 15304 7030 15356 7082
rect 15356 7030 15358 7082
rect 15302 7028 15358 7030
rect 15406 7082 15462 7084
rect 15406 7030 15408 7082
rect 15408 7030 15460 7082
rect 15460 7030 15462 7082
rect 15406 7028 15462 7030
rect 24522 7082 24578 7084
rect 24522 7030 24524 7082
rect 24524 7030 24576 7082
rect 24576 7030 24578 7082
rect 24522 7028 24578 7030
rect 24626 7082 24682 7084
rect 24626 7030 24628 7082
rect 24628 7030 24680 7082
rect 24680 7030 24682 7082
rect 24626 7028 24682 7030
rect 24730 7082 24786 7084
rect 24730 7030 24732 7082
rect 24732 7030 24784 7082
rect 24784 7030 24786 7082
rect 24730 7028 24786 7030
rect 33846 7082 33902 7084
rect 33846 7030 33848 7082
rect 33848 7030 33900 7082
rect 33900 7030 33902 7082
rect 33846 7028 33902 7030
rect 33950 7082 34006 7084
rect 33950 7030 33952 7082
rect 33952 7030 34004 7082
rect 34004 7030 34006 7082
rect 33950 7028 34006 7030
rect 34054 7082 34110 7084
rect 34054 7030 34056 7082
rect 34056 7030 34108 7082
rect 34108 7030 34110 7082
rect 34054 7028 34110 7030
rect 10536 6074 10592 6076
rect 10536 6022 10538 6074
rect 10538 6022 10590 6074
rect 10590 6022 10592 6074
rect 10536 6020 10592 6022
rect 10640 6074 10696 6076
rect 10640 6022 10642 6074
rect 10642 6022 10694 6074
rect 10694 6022 10696 6074
rect 10640 6020 10696 6022
rect 10744 6074 10800 6076
rect 10744 6022 10746 6074
rect 10746 6022 10798 6074
rect 10798 6022 10800 6074
rect 10744 6020 10800 6022
rect 19860 6074 19916 6076
rect 19860 6022 19862 6074
rect 19862 6022 19914 6074
rect 19914 6022 19916 6074
rect 19860 6020 19916 6022
rect 19964 6074 20020 6076
rect 19964 6022 19966 6074
rect 19966 6022 20018 6074
rect 20018 6022 20020 6074
rect 19964 6020 20020 6022
rect 20068 6074 20124 6076
rect 20068 6022 20070 6074
rect 20070 6022 20122 6074
rect 20122 6022 20124 6074
rect 20068 6020 20124 6022
rect 29184 6074 29240 6076
rect 29184 6022 29186 6074
rect 29186 6022 29238 6074
rect 29238 6022 29240 6074
rect 29184 6020 29240 6022
rect 29288 6074 29344 6076
rect 29288 6022 29290 6074
rect 29290 6022 29342 6074
rect 29342 6022 29344 6074
rect 29288 6020 29344 6022
rect 29392 6074 29448 6076
rect 29392 6022 29394 6074
rect 29394 6022 29446 6074
rect 29446 6022 29448 6074
rect 29392 6020 29448 6022
rect 38508 6074 38564 6076
rect 38508 6022 38510 6074
rect 38510 6022 38562 6074
rect 38562 6022 38564 6074
rect 38508 6020 38564 6022
rect 38612 6074 38668 6076
rect 38612 6022 38614 6074
rect 38614 6022 38666 6074
rect 38666 6022 38668 6074
rect 38612 6020 38668 6022
rect 38716 6074 38772 6076
rect 38716 6022 38718 6074
rect 38718 6022 38770 6074
rect 38770 6022 38772 6074
rect 38716 6020 38772 6022
rect 5874 5066 5930 5068
rect 5874 5014 5876 5066
rect 5876 5014 5928 5066
rect 5928 5014 5930 5066
rect 5874 5012 5930 5014
rect 5978 5066 6034 5068
rect 5978 5014 5980 5066
rect 5980 5014 6032 5066
rect 6032 5014 6034 5066
rect 5978 5012 6034 5014
rect 6082 5066 6138 5068
rect 6082 5014 6084 5066
rect 6084 5014 6136 5066
rect 6136 5014 6138 5066
rect 6082 5012 6138 5014
rect 15198 5066 15254 5068
rect 15198 5014 15200 5066
rect 15200 5014 15252 5066
rect 15252 5014 15254 5066
rect 15198 5012 15254 5014
rect 15302 5066 15358 5068
rect 15302 5014 15304 5066
rect 15304 5014 15356 5066
rect 15356 5014 15358 5066
rect 15302 5012 15358 5014
rect 15406 5066 15462 5068
rect 15406 5014 15408 5066
rect 15408 5014 15460 5066
rect 15460 5014 15462 5066
rect 15406 5012 15462 5014
rect 24522 5066 24578 5068
rect 24522 5014 24524 5066
rect 24524 5014 24576 5066
rect 24576 5014 24578 5066
rect 24522 5012 24578 5014
rect 24626 5066 24682 5068
rect 24626 5014 24628 5066
rect 24628 5014 24680 5066
rect 24680 5014 24682 5066
rect 24626 5012 24682 5014
rect 24730 5066 24786 5068
rect 24730 5014 24732 5066
rect 24732 5014 24784 5066
rect 24784 5014 24786 5066
rect 24730 5012 24786 5014
rect 33846 5066 33902 5068
rect 33846 5014 33848 5066
rect 33848 5014 33900 5066
rect 33900 5014 33902 5066
rect 33846 5012 33902 5014
rect 33950 5066 34006 5068
rect 33950 5014 33952 5066
rect 33952 5014 34004 5066
rect 34004 5014 34006 5066
rect 33950 5012 34006 5014
rect 34054 5066 34110 5068
rect 34054 5014 34056 5066
rect 34056 5014 34108 5066
rect 34108 5014 34110 5066
rect 34054 5012 34110 5014
rect 10536 4058 10592 4060
rect 10536 4006 10538 4058
rect 10538 4006 10590 4058
rect 10590 4006 10592 4058
rect 10536 4004 10592 4006
rect 10640 4058 10696 4060
rect 10640 4006 10642 4058
rect 10642 4006 10694 4058
rect 10694 4006 10696 4058
rect 10640 4004 10696 4006
rect 10744 4058 10800 4060
rect 10744 4006 10746 4058
rect 10746 4006 10798 4058
rect 10798 4006 10800 4058
rect 10744 4004 10800 4006
rect 19860 4058 19916 4060
rect 19860 4006 19862 4058
rect 19862 4006 19914 4058
rect 19914 4006 19916 4058
rect 19860 4004 19916 4006
rect 19964 4058 20020 4060
rect 19964 4006 19966 4058
rect 19966 4006 20018 4058
rect 20018 4006 20020 4058
rect 19964 4004 20020 4006
rect 20068 4058 20124 4060
rect 20068 4006 20070 4058
rect 20070 4006 20122 4058
rect 20122 4006 20124 4058
rect 20068 4004 20124 4006
rect 29184 4058 29240 4060
rect 29184 4006 29186 4058
rect 29186 4006 29238 4058
rect 29238 4006 29240 4058
rect 29184 4004 29240 4006
rect 29288 4058 29344 4060
rect 29288 4006 29290 4058
rect 29290 4006 29342 4058
rect 29342 4006 29344 4058
rect 29288 4004 29344 4006
rect 29392 4058 29448 4060
rect 29392 4006 29394 4058
rect 29394 4006 29446 4058
rect 29446 4006 29448 4058
rect 29392 4004 29448 4006
rect 38508 4058 38564 4060
rect 38508 4006 38510 4058
rect 38510 4006 38562 4058
rect 38562 4006 38564 4058
rect 38508 4004 38564 4006
rect 38612 4058 38668 4060
rect 38612 4006 38614 4058
rect 38614 4006 38666 4058
rect 38666 4006 38668 4058
rect 38612 4004 38668 4006
rect 38716 4058 38772 4060
rect 38716 4006 38718 4058
rect 38718 4006 38770 4058
rect 38770 4006 38772 4058
rect 38716 4004 38772 4006
<< metal3 >>
rect 10526 36260 10536 36316
rect 10592 36260 10640 36316
rect 10696 36260 10744 36316
rect 10800 36260 10810 36316
rect 19850 36260 19860 36316
rect 19916 36260 19964 36316
rect 20020 36260 20068 36316
rect 20124 36260 20134 36316
rect 29174 36260 29184 36316
rect 29240 36260 29288 36316
rect 29344 36260 29392 36316
rect 29448 36260 29458 36316
rect 38498 36260 38508 36316
rect 38564 36260 38612 36316
rect 38668 36260 38716 36316
rect 38772 36260 38782 36316
rect 5864 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6148 35308
rect 15188 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15472 35308
rect 24512 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24796 35308
rect 33836 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34120 35308
rect 10526 34244 10536 34300
rect 10592 34244 10640 34300
rect 10696 34244 10744 34300
rect 10800 34244 10810 34300
rect 19850 34244 19860 34300
rect 19916 34244 19964 34300
rect 20020 34244 20068 34300
rect 20124 34244 20134 34300
rect 29174 34244 29184 34300
rect 29240 34244 29288 34300
rect 29344 34244 29392 34300
rect 29448 34244 29458 34300
rect 38498 34244 38508 34300
rect 38564 34244 38612 34300
rect 38668 34244 38716 34300
rect 38772 34244 38782 34300
rect 5864 33236 5874 33292
rect 5930 33236 5978 33292
rect 6034 33236 6082 33292
rect 6138 33236 6148 33292
rect 15188 33236 15198 33292
rect 15254 33236 15302 33292
rect 15358 33236 15406 33292
rect 15462 33236 15472 33292
rect 24512 33236 24522 33292
rect 24578 33236 24626 33292
rect 24682 33236 24730 33292
rect 24786 33236 24796 33292
rect 33836 33236 33846 33292
rect 33902 33236 33950 33292
rect 34006 33236 34054 33292
rect 34110 33236 34120 33292
rect 10526 32228 10536 32284
rect 10592 32228 10640 32284
rect 10696 32228 10744 32284
rect 10800 32228 10810 32284
rect 19850 32228 19860 32284
rect 19916 32228 19964 32284
rect 20020 32228 20068 32284
rect 20124 32228 20134 32284
rect 29174 32228 29184 32284
rect 29240 32228 29288 32284
rect 29344 32228 29392 32284
rect 29448 32228 29458 32284
rect 38498 32228 38508 32284
rect 38564 32228 38612 32284
rect 38668 32228 38716 32284
rect 38772 32228 38782 32284
rect 5864 31220 5874 31276
rect 5930 31220 5978 31276
rect 6034 31220 6082 31276
rect 6138 31220 6148 31276
rect 15188 31220 15198 31276
rect 15254 31220 15302 31276
rect 15358 31220 15406 31276
rect 15462 31220 15472 31276
rect 24512 31220 24522 31276
rect 24578 31220 24626 31276
rect 24682 31220 24730 31276
rect 24786 31220 24796 31276
rect 33836 31220 33846 31276
rect 33902 31220 33950 31276
rect 34006 31220 34054 31276
rect 34110 31220 34120 31276
rect 10526 30212 10536 30268
rect 10592 30212 10640 30268
rect 10696 30212 10744 30268
rect 10800 30212 10810 30268
rect 19850 30212 19860 30268
rect 19916 30212 19964 30268
rect 20020 30212 20068 30268
rect 20124 30212 20134 30268
rect 29174 30212 29184 30268
rect 29240 30212 29288 30268
rect 29344 30212 29392 30268
rect 29448 30212 29458 30268
rect 38498 30212 38508 30268
rect 38564 30212 38612 30268
rect 38668 30212 38716 30268
rect 38772 30212 38782 30268
rect 5864 29204 5874 29260
rect 5930 29204 5978 29260
rect 6034 29204 6082 29260
rect 6138 29204 6148 29260
rect 15188 29204 15198 29260
rect 15254 29204 15302 29260
rect 15358 29204 15406 29260
rect 15462 29204 15472 29260
rect 24512 29204 24522 29260
rect 24578 29204 24626 29260
rect 24682 29204 24730 29260
rect 24786 29204 24796 29260
rect 33836 29204 33846 29260
rect 33902 29204 33950 29260
rect 34006 29204 34054 29260
rect 34110 29204 34120 29260
rect 10526 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10810 28252
rect 19850 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20134 28252
rect 29174 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29458 28252
rect 38498 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38782 28252
rect 5864 27188 5874 27244
rect 5930 27188 5978 27244
rect 6034 27188 6082 27244
rect 6138 27188 6148 27244
rect 15188 27188 15198 27244
rect 15254 27188 15302 27244
rect 15358 27188 15406 27244
rect 15462 27188 15472 27244
rect 24512 27188 24522 27244
rect 24578 27188 24626 27244
rect 24682 27188 24730 27244
rect 24786 27188 24796 27244
rect 33836 27188 33846 27244
rect 33902 27188 33950 27244
rect 34006 27188 34054 27244
rect 34110 27188 34120 27244
rect 10526 26180 10536 26236
rect 10592 26180 10640 26236
rect 10696 26180 10744 26236
rect 10800 26180 10810 26236
rect 19850 26180 19860 26236
rect 19916 26180 19964 26236
rect 20020 26180 20068 26236
rect 20124 26180 20134 26236
rect 29174 26180 29184 26236
rect 29240 26180 29288 26236
rect 29344 26180 29392 26236
rect 29448 26180 29458 26236
rect 38498 26180 38508 26236
rect 38564 26180 38612 26236
rect 38668 26180 38716 26236
rect 38772 26180 38782 26236
rect 39200 25620 40000 25648
rect 34514 25564 34524 25620
rect 34580 25564 40000 25620
rect 39200 25536 40000 25564
rect 5864 25172 5874 25228
rect 5930 25172 5978 25228
rect 6034 25172 6082 25228
rect 6138 25172 6148 25228
rect 15188 25172 15198 25228
rect 15254 25172 15302 25228
rect 15358 25172 15406 25228
rect 15462 25172 15472 25228
rect 24512 25172 24522 25228
rect 24578 25172 24626 25228
rect 24682 25172 24730 25228
rect 24786 25172 24796 25228
rect 33836 25172 33846 25228
rect 33902 25172 33950 25228
rect 34006 25172 34054 25228
rect 34110 25172 34120 25228
rect 39200 24948 40000 24976
rect 34738 24892 34748 24948
rect 34804 24892 40000 24948
rect 39200 24864 40000 24892
rect 0 24276 800 24304
rect 39200 24276 40000 24304
rect 0 24220 4172 24276
rect 4228 24220 4238 24276
rect 38892 24220 40000 24276
rect 0 24192 800 24220
rect 10526 24164 10536 24220
rect 10592 24164 10640 24220
rect 10696 24164 10744 24220
rect 10800 24164 10810 24220
rect 19850 24164 19860 24220
rect 19916 24164 19964 24220
rect 20020 24164 20068 24220
rect 20124 24164 20134 24220
rect 29174 24164 29184 24220
rect 29240 24164 29288 24220
rect 29344 24164 29392 24220
rect 29448 24164 29458 24220
rect 38498 24164 38508 24220
rect 38564 24164 38612 24220
rect 38668 24164 38716 24220
rect 38772 24164 38782 24220
rect 38892 24052 38948 24220
rect 39200 24192 40000 24220
rect 35074 23996 35084 24052
rect 35140 23996 38948 24052
rect 0 23604 800 23632
rect 39200 23604 40000 23632
rect 0 23548 4060 23604
rect 4116 23548 4126 23604
rect 35186 23548 35196 23604
rect 35252 23548 40000 23604
rect 0 23520 800 23548
rect 39200 23520 40000 23548
rect 5864 23156 5874 23212
rect 5930 23156 5978 23212
rect 6034 23156 6082 23212
rect 6138 23156 6148 23212
rect 15188 23156 15198 23212
rect 15254 23156 15302 23212
rect 15358 23156 15406 23212
rect 15462 23156 15472 23212
rect 24512 23156 24522 23212
rect 24578 23156 24626 23212
rect 24682 23156 24730 23212
rect 24786 23156 24796 23212
rect 33836 23156 33846 23212
rect 33902 23156 33950 23212
rect 34006 23156 34054 23212
rect 34110 23156 34120 23212
rect 0 22932 800 22960
rect 39200 22932 40000 22960
rect 0 22876 4284 22932
rect 4340 22876 4350 22932
rect 34962 22876 34972 22932
rect 35028 22876 40000 22932
rect 0 22848 800 22876
rect 39200 22848 40000 22876
rect 4162 22652 4172 22708
rect 4228 22652 13580 22708
rect 13636 22652 13646 22708
rect 0 22260 800 22288
rect 39200 22260 40000 22288
rect 0 22204 8428 22260
rect 38892 22204 40000 22260
rect 0 22176 800 22204
rect 8372 21924 8428 22204
rect 10526 22148 10536 22204
rect 10592 22148 10640 22204
rect 10696 22148 10744 22204
rect 10800 22148 10810 22204
rect 19850 22148 19860 22204
rect 19916 22148 19964 22204
rect 20020 22148 20068 22204
rect 20124 22148 20134 22204
rect 29174 22148 29184 22204
rect 29240 22148 29288 22204
rect 29344 22148 29392 22204
rect 29448 22148 29458 22204
rect 38498 22148 38508 22204
rect 38564 22148 38612 22204
rect 38668 22148 38716 22204
rect 38772 22148 38782 22204
rect 38892 22036 38948 22204
rect 39200 22176 40000 22204
rect 34850 21980 34860 22036
rect 34916 21980 38948 22036
rect 8372 21868 17948 21924
rect 18004 21868 18014 21924
rect 31042 21868 31052 21924
rect 31108 21868 35196 21924
rect 35252 21868 35262 21924
rect 22082 21756 22092 21812
rect 22148 21756 35084 21812
rect 35140 21756 35150 21812
rect 0 21588 800 21616
rect 39200 21588 40000 21616
rect 0 21532 19292 21588
rect 19348 21532 19358 21588
rect 27346 21532 27356 21588
rect 27412 21532 40000 21588
rect 0 21504 800 21532
rect 39200 21504 40000 21532
rect 5864 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6148 21196
rect 15188 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15472 21196
rect 24512 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24796 21196
rect 33836 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34120 21196
rect 0 20916 800 20944
rect 39200 20916 40000 20944
rect 0 20860 18060 20916
rect 18116 20860 18126 20916
rect 25106 20860 25116 20916
rect 25172 20860 34972 20916
rect 35028 20860 35038 20916
rect 35644 20860 40000 20916
rect 0 20832 800 20860
rect 28130 20748 28140 20804
rect 28196 20748 34748 20804
rect 34804 20748 34814 20804
rect 4274 20636 4284 20692
rect 4340 20636 14924 20692
rect 14980 20636 14990 20692
rect 22306 20636 22316 20692
rect 22372 20636 34860 20692
rect 34916 20636 34926 20692
rect 4050 20524 4060 20580
rect 4116 20524 17612 20580
rect 17668 20524 18284 20580
rect 18340 20524 18350 20580
rect 20850 20524 20860 20580
rect 20916 20524 23436 20580
rect 23492 20524 23502 20580
rect 24322 20524 24332 20580
rect 24388 20524 34300 20580
rect 34356 20524 34366 20580
rect 24332 20468 24388 20524
rect 35644 20468 35700 20860
rect 39200 20832 40000 20860
rect 4284 20412 12460 20468
rect 12516 20412 13692 20468
rect 13748 20412 13758 20468
rect 21970 20412 21980 20468
rect 22036 20412 22876 20468
rect 22932 20412 24388 20468
rect 28924 20412 30716 20468
rect 30772 20412 30782 20468
rect 31892 20412 35700 20468
rect 0 20244 800 20272
rect 4284 20244 4340 20412
rect 28924 20356 28980 20412
rect 31892 20356 31948 20412
rect 4610 20300 4620 20356
rect 4676 20300 12908 20356
rect 12964 20300 13804 20356
rect 13860 20300 13870 20356
rect 20738 20300 20748 20356
rect 20804 20300 21532 20356
rect 21588 20300 21598 20356
rect 28914 20300 28924 20356
rect 28980 20300 28990 20356
rect 29586 20300 29596 20356
rect 29652 20300 31948 20356
rect 34626 20300 34636 20356
rect 34692 20300 38948 20356
rect 38892 20244 38948 20300
rect 39200 20244 40000 20272
rect 0 20188 4340 20244
rect 23650 20188 23660 20244
rect 23716 20188 25116 20244
rect 25172 20188 25182 20244
rect 26450 20188 26460 20244
rect 26516 20188 27244 20244
rect 27300 20188 28140 20244
rect 28196 20188 28206 20244
rect 38892 20188 40000 20244
rect 0 20160 800 20188
rect 10526 20132 10536 20188
rect 10592 20132 10640 20188
rect 10696 20132 10744 20188
rect 10800 20132 10810 20188
rect 19850 20132 19860 20188
rect 19916 20132 19964 20188
rect 20020 20132 20068 20188
rect 20124 20132 20134 20188
rect 29174 20132 29184 20188
rect 29240 20132 29288 20188
rect 29344 20132 29392 20188
rect 29448 20132 29458 20188
rect 38498 20132 38508 20188
rect 38564 20132 38612 20188
rect 38668 20132 38716 20188
rect 38772 20132 38782 20188
rect 39200 20160 40000 20188
rect 30930 19964 30940 20020
rect 30996 19964 31948 20020
rect 32004 19964 34636 20020
rect 34692 19964 34702 20020
rect 16706 19852 16716 19908
rect 16772 19852 18844 19908
rect 18900 19852 18910 19908
rect 22866 19852 22876 19908
rect 22932 19852 25340 19908
rect 25396 19852 34524 19908
rect 34580 19852 34590 19908
rect 31500 19740 31948 19796
rect 0 19572 800 19600
rect 31500 19572 31556 19740
rect 31892 19572 31948 19740
rect 39200 19572 40000 19600
rect 0 19516 13468 19572
rect 13524 19516 14028 19572
rect 14084 19516 14094 19572
rect 24322 19516 24332 19572
rect 24388 19516 25788 19572
rect 25844 19516 25854 19572
rect 26338 19516 26348 19572
rect 26404 19516 30044 19572
rect 30100 19516 30110 19572
rect 30706 19516 30716 19572
rect 30772 19516 31500 19572
rect 31556 19516 31566 19572
rect 31892 19516 40000 19572
rect 0 19488 800 19516
rect 39200 19488 40000 19516
rect 5864 19124 5874 19180
rect 5930 19124 5978 19180
rect 6034 19124 6082 19180
rect 6138 19124 6148 19180
rect 15188 19124 15198 19180
rect 15254 19124 15302 19180
rect 15358 19124 15406 19180
rect 15462 19124 15472 19180
rect 24512 19124 24522 19180
rect 24578 19124 24626 19180
rect 24682 19124 24730 19180
rect 24786 19124 24796 19180
rect 33836 19124 33846 19180
rect 33902 19124 33950 19180
rect 34006 19124 34054 19180
rect 34110 19124 34120 19180
rect 0 18900 800 18928
rect 39200 18900 40000 18928
rect 0 18844 15932 18900
rect 15988 18844 16828 18900
rect 16884 18844 16894 18900
rect 30034 18844 30044 18900
rect 30100 18844 35084 18900
rect 35140 18844 35150 18900
rect 35532 18844 40000 18900
rect 0 18816 800 18844
rect 4050 18732 4060 18788
rect 4116 18732 16268 18788
rect 16324 18732 16940 18788
rect 16996 18732 17006 18788
rect 26002 18732 26012 18788
rect 26068 18732 35196 18788
rect 35252 18732 35262 18788
rect 4274 18620 4284 18676
rect 4340 18620 11564 18676
rect 11620 18620 12124 18676
rect 12180 18620 12190 18676
rect 29698 18620 29708 18676
rect 29764 18620 30604 18676
rect 30660 18620 30670 18676
rect 35532 18564 35588 18844
rect 39200 18816 40000 18844
rect 4162 18508 4172 18564
rect 4228 18508 11116 18564
rect 11172 18508 12012 18564
rect 12068 18508 12078 18564
rect 26898 18508 26908 18564
rect 26964 18508 27916 18564
rect 27972 18508 28588 18564
rect 28644 18508 35588 18564
rect 30034 18396 30044 18452
rect 30100 18396 38948 18452
rect 0 18228 800 18256
rect 38892 18228 38948 18396
rect 39200 18228 40000 18256
rect 0 18172 4620 18228
rect 4676 18172 4686 18228
rect 38892 18172 40000 18228
rect 0 18144 800 18172
rect 10526 18116 10536 18172
rect 10592 18116 10640 18172
rect 10696 18116 10744 18172
rect 10800 18116 10810 18172
rect 19850 18116 19860 18172
rect 19916 18116 19964 18172
rect 20020 18116 20068 18172
rect 20124 18116 20134 18172
rect 29174 18116 29184 18172
rect 29240 18116 29288 18172
rect 29344 18116 29392 18172
rect 29448 18116 29458 18172
rect 38498 18116 38508 18172
rect 38564 18116 38612 18172
rect 38668 18116 38716 18172
rect 38772 18116 38782 18172
rect 39200 18144 40000 18172
rect 0 17556 800 17584
rect 39200 17556 40000 17584
rect 0 17500 4172 17556
rect 4228 17500 4238 17556
rect 23426 17500 23436 17556
rect 23492 17500 26012 17556
rect 26068 17500 40000 17556
rect 0 17472 800 17500
rect 39200 17472 40000 17500
rect 5864 17108 5874 17164
rect 5930 17108 5978 17164
rect 6034 17108 6082 17164
rect 6138 17108 6148 17164
rect 15188 17108 15198 17164
rect 15254 17108 15302 17164
rect 15358 17108 15406 17164
rect 15462 17108 15472 17164
rect 24512 17108 24522 17164
rect 24578 17108 24626 17164
rect 24682 17108 24730 17164
rect 24786 17108 24796 17164
rect 33836 17108 33846 17164
rect 33902 17108 33950 17164
rect 34006 17108 34054 17164
rect 34110 17108 34120 17164
rect 0 16884 800 16912
rect 39200 16884 40000 16912
rect 0 16828 4284 16884
rect 4340 16828 4350 16884
rect 35186 16828 35196 16884
rect 35252 16828 40000 16884
rect 0 16800 800 16828
rect 39200 16800 40000 16828
rect 35074 16268 35084 16324
rect 35140 16268 38948 16324
rect 0 16212 800 16240
rect 38892 16212 38948 16268
rect 39200 16212 40000 16240
rect 0 16156 4060 16212
rect 4116 16156 4126 16212
rect 38892 16156 40000 16212
rect 0 16128 800 16156
rect 10526 16100 10536 16156
rect 10592 16100 10640 16156
rect 10696 16100 10744 16156
rect 10800 16100 10810 16156
rect 19850 16100 19860 16156
rect 19916 16100 19964 16156
rect 20020 16100 20068 16156
rect 20124 16100 20134 16156
rect 29174 16100 29184 16156
rect 29240 16100 29288 16156
rect 29344 16100 29392 16156
rect 29448 16100 29458 16156
rect 38498 16100 38508 16156
rect 38564 16100 38612 16156
rect 38668 16100 38716 16156
rect 38772 16100 38782 16156
rect 39200 16128 40000 16156
rect 39200 15540 40000 15568
rect 24882 15484 24892 15540
rect 24948 15484 40000 15540
rect 39200 15456 40000 15484
rect 5864 15092 5874 15148
rect 5930 15092 5978 15148
rect 6034 15092 6082 15148
rect 6138 15092 6148 15148
rect 15188 15092 15198 15148
rect 15254 15092 15302 15148
rect 15358 15092 15406 15148
rect 15462 15092 15472 15148
rect 24512 15092 24522 15148
rect 24578 15092 24626 15148
rect 24682 15092 24730 15148
rect 24786 15092 24796 15148
rect 33836 15092 33846 15148
rect 33902 15092 33950 15148
rect 34006 15092 34054 15148
rect 34110 15092 34120 15148
rect 39200 14868 40000 14896
rect 34290 14812 34300 14868
rect 34356 14812 40000 14868
rect 39200 14784 40000 14812
rect 10526 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10810 14140
rect 19850 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20134 14140
rect 29174 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29458 14140
rect 38498 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38782 14140
rect 5864 13076 5874 13132
rect 5930 13076 5978 13132
rect 6034 13076 6082 13132
rect 6138 13076 6148 13132
rect 15188 13076 15198 13132
rect 15254 13076 15302 13132
rect 15358 13076 15406 13132
rect 15462 13076 15472 13132
rect 24512 13076 24522 13132
rect 24578 13076 24626 13132
rect 24682 13076 24730 13132
rect 24786 13076 24796 13132
rect 33836 13076 33846 13132
rect 33902 13076 33950 13132
rect 34006 13076 34054 13132
rect 34110 13076 34120 13132
rect 10526 12068 10536 12124
rect 10592 12068 10640 12124
rect 10696 12068 10744 12124
rect 10800 12068 10810 12124
rect 19850 12068 19860 12124
rect 19916 12068 19964 12124
rect 20020 12068 20068 12124
rect 20124 12068 20134 12124
rect 29174 12068 29184 12124
rect 29240 12068 29288 12124
rect 29344 12068 29392 12124
rect 29448 12068 29458 12124
rect 38498 12068 38508 12124
rect 38564 12068 38612 12124
rect 38668 12068 38716 12124
rect 38772 12068 38782 12124
rect 5864 11060 5874 11116
rect 5930 11060 5978 11116
rect 6034 11060 6082 11116
rect 6138 11060 6148 11116
rect 15188 11060 15198 11116
rect 15254 11060 15302 11116
rect 15358 11060 15406 11116
rect 15462 11060 15472 11116
rect 24512 11060 24522 11116
rect 24578 11060 24626 11116
rect 24682 11060 24730 11116
rect 24786 11060 24796 11116
rect 33836 11060 33846 11116
rect 33902 11060 33950 11116
rect 34006 11060 34054 11116
rect 34110 11060 34120 11116
rect 10526 10052 10536 10108
rect 10592 10052 10640 10108
rect 10696 10052 10744 10108
rect 10800 10052 10810 10108
rect 19850 10052 19860 10108
rect 19916 10052 19964 10108
rect 20020 10052 20068 10108
rect 20124 10052 20134 10108
rect 29174 10052 29184 10108
rect 29240 10052 29288 10108
rect 29344 10052 29392 10108
rect 29448 10052 29458 10108
rect 38498 10052 38508 10108
rect 38564 10052 38612 10108
rect 38668 10052 38716 10108
rect 38772 10052 38782 10108
rect 5864 9044 5874 9100
rect 5930 9044 5978 9100
rect 6034 9044 6082 9100
rect 6138 9044 6148 9100
rect 15188 9044 15198 9100
rect 15254 9044 15302 9100
rect 15358 9044 15406 9100
rect 15462 9044 15472 9100
rect 24512 9044 24522 9100
rect 24578 9044 24626 9100
rect 24682 9044 24730 9100
rect 24786 9044 24796 9100
rect 33836 9044 33846 9100
rect 33902 9044 33950 9100
rect 34006 9044 34054 9100
rect 34110 9044 34120 9100
rect 10526 8036 10536 8092
rect 10592 8036 10640 8092
rect 10696 8036 10744 8092
rect 10800 8036 10810 8092
rect 19850 8036 19860 8092
rect 19916 8036 19964 8092
rect 20020 8036 20068 8092
rect 20124 8036 20134 8092
rect 29174 8036 29184 8092
rect 29240 8036 29288 8092
rect 29344 8036 29392 8092
rect 29448 8036 29458 8092
rect 38498 8036 38508 8092
rect 38564 8036 38612 8092
rect 38668 8036 38716 8092
rect 38772 8036 38782 8092
rect 5864 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6148 7084
rect 15188 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15472 7084
rect 24512 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24796 7084
rect 33836 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34120 7084
rect 10526 6020 10536 6076
rect 10592 6020 10640 6076
rect 10696 6020 10744 6076
rect 10800 6020 10810 6076
rect 19850 6020 19860 6076
rect 19916 6020 19964 6076
rect 20020 6020 20068 6076
rect 20124 6020 20134 6076
rect 29174 6020 29184 6076
rect 29240 6020 29288 6076
rect 29344 6020 29392 6076
rect 29448 6020 29458 6076
rect 38498 6020 38508 6076
rect 38564 6020 38612 6076
rect 38668 6020 38716 6076
rect 38772 6020 38782 6076
rect 5864 5012 5874 5068
rect 5930 5012 5978 5068
rect 6034 5012 6082 5068
rect 6138 5012 6148 5068
rect 15188 5012 15198 5068
rect 15254 5012 15302 5068
rect 15358 5012 15406 5068
rect 15462 5012 15472 5068
rect 24512 5012 24522 5068
rect 24578 5012 24626 5068
rect 24682 5012 24730 5068
rect 24786 5012 24796 5068
rect 33836 5012 33846 5068
rect 33902 5012 33950 5068
rect 34006 5012 34054 5068
rect 34110 5012 34120 5068
rect 10526 4004 10536 4060
rect 10592 4004 10640 4060
rect 10696 4004 10744 4060
rect 10800 4004 10810 4060
rect 19850 4004 19860 4060
rect 19916 4004 19964 4060
rect 20020 4004 20068 4060
rect 20124 4004 20134 4060
rect 29174 4004 29184 4060
rect 29240 4004 29288 4060
rect 29344 4004 29392 4060
rect 29448 4004 29458 4060
rect 38498 4004 38508 4060
rect 38564 4004 38612 4060
rect 38668 4004 38716 4060
rect 38772 4004 38782 4060
<< via3 >>
rect 10536 36260 10592 36316
rect 10640 36260 10696 36316
rect 10744 36260 10800 36316
rect 19860 36260 19916 36316
rect 19964 36260 20020 36316
rect 20068 36260 20124 36316
rect 29184 36260 29240 36316
rect 29288 36260 29344 36316
rect 29392 36260 29448 36316
rect 38508 36260 38564 36316
rect 38612 36260 38668 36316
rect 38716 36260 38772 36316
rect 5874 35252 5930 35308
rect 5978 35252 6034 35308
rect 6082 35252 6138 35308
rect 15198 35252 15254 35308
rect 15302 35252 15358 35308
rect 15406 35252 15462 35308
rect 24522 35252 24578 35308
rect 24626 35252 24682 35308
rect 24730 35252 24786 35308
rect 33846 35252 33902 35308
rect 33950 35252 34006 35308
rect 34054 35252 34110 35308
rect 10536 34244 10592 34300
rect 10640 34244 10696 34300
rect 10744 34244 10800 34300
rect 19860 34244 19916 34300
rect 19964 34244 20020 34300
rect 20068 34244 20124 34300
rect 29184 34244 29240 34300
rect 29288 34244 29344 34300
rect 29392 34244 29448 34300
rect 38508 34244 38564 34300
rect 38612 34244 38668 34300
rect 38716 34244 38772 34300
rect 5874 33236 5930 33292
rect 5978 33236 6034 33292
rect 6082 33236 6138 33292
rect 15198 33236 15254 33292
rect 15302 33236 15358 33292
rect 15406 33236 15462 33292
rect 24522 33236 24578 33292
rect 24626 33236 24682 33292
rect 24730 33236 24786 33292
rect 33846 33236 33902 33292
rect 33950 33236 34006 33292
rect 34054 33236 34110 33292
rect 10536 32228 10592 32284
rect 10640 32228 10696 32284
rect 10744 32228 10800 32284
rect 19860 32228 19916 32284
rect 19964 32228 20020 32284
rect 20068 32228 20124 32284
rect 29184 32228 29240 32284
rect 29288 32228 29344 32284
rect 29392 32228 29448 32284
rect 38508 32228 38564 32284
rect 38612 32228 38668 32284
rect 38716 32228 38772 32284
rect 5874 31220 5930 31276
rect 5978 31220 6034 31276
rect 6082 31220 6138 31276
rect 15198 31220 15254 31276
rect 15302 31220 15358 31276
rect 15406 31220 15462 31276
rect 24522 31220 24578 31276
rect 24626 31220 24682 31276
rect 24730 31220 24786 31276
rect 33846 31220 33902 31276
rect 33950 31220 34006 31276
rect 34054 31220 34110 31276
rect 10536 30212 10592 30268
rect 10640 30212 10696 30268
rect 10744 30212 10800 30268
rect 19860 30212 19916 30268
rect 19964 30212 20020 30268
rect 20068 30212 20124 30268
rect 29184 30212 29240 30268
rect 29288 30212 29344 30268
rect 29392 30212 29448 30268
rect 38508 30212 38564 30268
rect 38612 30212 38668 30268
rect 38716 30212 38772 30268
rect 5874 29204 5930 29260
rect 5978 29204 6034 29260
rect 6082 29204 6138 29260
rect 15198 29204 15254 29260
rect 15302 29204 15358 29260
rect 15406 29204 15462 29260
rect 24522 29204 24578 29260
rect 24626 29204 24682 29260
rect 24730 29204 24786 29260
rect 33846 29204 33902 29260
rect 33950 29204 34006 29260
rect 34054 29204 34110 29260
rect 10536 28196 10592 28252
rect 10640 28196 10696 28252
rect 10744 28196 10800 28252
rect 19860 28196 19916 28252
rect 19964 28196 20020 28252
rect 20068 28196 20124 28252
rect 29184 28196 29240 28252
rect 29288 28196 29344 28252
rect 29392 28196 29448 28252
rect 38508 28196 38564 28252
rect 38612 28196 38668 28252
rect 38716 28196 38772 28252
rect 5874 27188 5930 27244
rect 5978 27188 6034 27244
rect 6082 27188 6138 27244
rect 15198 27188 15254 27244
rect 15302 27188 15358 27244
rect 15406 27188 15462 27244
rect 24522 27188 24578 27244
rect 24626 27188 24682 27244
rect 24730 27188 24786 27244
rect 33846 27188 33902 27244
rect 33950 27188 34006 27244
rect 34054 27188 34110 27244
rect 10536 26180 10592 26236
rect 10640 26180 10696 26236
rect 10744 26180 10800 26236
rect 19860 26180 19916 26236
rect 19964 26180 20020 26236
rect 20068 26180 20124 26236
rect 29184 26180 29240 26236
rect 29288 26180 29344 26236
rect 29392 26180 29448 26236
rect 38508 26180 38564 26236
rect 38612 26180 38668 26236
rect 38716 26180 38772 26236
rect 5874 25172 5930 25228
rect 5978 25172 6034 25228
rect 6082 25172 6138 25228
rect 15198 25172 15254 25228
rect 15302 25172 15358 25228
rect 15406 25172 15462 25228
rect 24522 25172 24578 25228
rect 24626 25172 24682 25228
rect 24730 25172 24786 25228
rect 33846 25172 33902 25228
rect 33950 25172 34006 25228
rect 34054 25172 34110 25228
rect 10536 24164 10592 24220
rect 10640 24164 10696 24220
rect 10744 24164 10800 24220
rect 19860 24164 19916 24220
rect 19964 24164 20020 24220
rect 20068 24164 20124 24220
rect 29184 24164 29240 24220
rect 29288 24164 29344 24220
rect 29392 24164 29448 24220
rect 38508 24164 38564 24220
rect 38612 24164 38668 24220
rect 38716 24164 38772 24220
rect 5874 23156 5930 23212
rect 5978 23156 6034 23212
rect 6082 23156 6138 23212
rect 15198 23156 15254 23212
rect 15302 23156 15358 23212
rect 15406 23156 15462 23212
rect 24522 23156 24578 23212
rect 24626 23156 24682 23212
rect 24730 23156 24786 23212
rect 33846 23156 33902 23212
rect 33950 23156 34006 23212
rect 34054 23156 34110 23212
rect 10536 22148 10592 22204
rect 10640 22148 10696 22204
rect 10744 22148 10800 22204
rect 19860 22148 19916 22204
rect 19964 22148 20020 22204
rect 20068 22148 20124 22204
rect 29184 22148 29240 22204
rect 29288 22148 29344 22204
rect 29392 22148 29448 22204
rect 38508 22148 38564 22204
rect 38612 22148 38668 22204
rect 38716 22148 38772 22204
rect 5874 21140 5930 21196
rect 5978 21140 6034 21196
rect 6082 21140 6138 21196
rect 15198 21140 15254 21196
rect 15302 21140 15358 21196
rect 15406 21140 15462 21196
rect 24522 21140 24578 21196
rect 24626 21140 24682 21196
rect 24730 21140 24786 21196
rect 33846 21140 33902 21196
rect 33950 21140 34006 21196
rect 34054 21140 34110 21196
rect 10536 20132 10592 20188
rect 10640 20132 10696 20188
rect 10744 20132 10800 20188
rect 19860 20132 19916 20188
rect 19964 20132 20020 20188
rect 20068 20132 20124 20188
rect 29184 20132 29240 20188
rect 29288 20132 29344 20188
rect 29392 20132 29448 20188
rect 38508 20132 38564 20188
rect 38612 20132 38668 20188
rect 38716 20132 38772 20188
rect 5874 19124 5930 19180
rect 5978 19124 6034 19180
rect 6082 19124 6138 19180
rect 15198 19124 15254 19180
rect 15302 19124 15358 19180
rect 15406 19124 15462 19180
rect 24522 19124 24578 19180
rect 24626 19124 24682 19180
rect 24730 19124 24786 19180
rect 33846 19124 33902 19180
rect 33950 19124 34006 19180
rect 34054 19124 34110 19180
rect 10536 18116 10592 18172
rect 10640 18116 10696 18172
rect 10744 18116 10800 18172
rect 19860 18116 19916 18172
rect 19964 18116 20020 18172
rect 20068 18116 20124 18172
rect 29184 18116 29240 18172
rect 29288 18116 29344 18172
rect 29392 18116 29448 18172
rect 38508 18116 38564 18172
rect 38612 18116 38668 18172
rect 38716 18116 38772 18172
rect 5874 17108 5930 17164
rect 5978 17108 6034 17164
rect 6082 17108 6138 17164
rect 15198 17108 15254 17164
rect 15302 17108 15358 17164
rect 15406 17108 15462 17164
rect 24522 17108 24578 17164
rect 24626 17108 24682 17164
rect 24730 17108 24786 17164
rect 33846 17108 33902 17164
rect 33950 17108 34006 17164
rect 34054 17108 34110 17164
rect 10536 16100 10592 16156
rect 10640 16100 10696 16156
rect 10744 16100 10800 16156
rect 19860 16100 19916 16156
rect 19964 16100 20020 16156
rect 20068 16100 20124 16156
rect 29184 16100 29240 16156
rect 29288 16100 29344 16156
rect 29392 16100 29448 16156
rect 38508 16100 38564 16156
rect 38612 16100 38668 16156
rect 38716 16100 38772 16156
rect 5874 15092 5930 15148
rect 5978 15092 6034 15148
rect 6082 15092 6138 15148
rect 15198 15092 15254 15148
rect 15302 15092 15358 15148
rect 15406 15092 15462 15148
rect 24522 15092 24578 15148
rect 24626 15092 24682 15148
rect 24730 15092 24786 15148
rect 33846 15092 33902 15148
rect 33950 15092 34006 15148
rect 34054 15092 34110 15148
rect 10536 14084 10592 14140
rect 10640 14084 10696 14140
rect 10744 14084 10800 14140
rect 19860 14084 19916 14140
rect 19964 14084 20020 14140
rect 20068 14084 20124 14140
rect 29184 14084 29240 14140
rect 29288 14084 29344 14140
rect 29392 14084 29448 14140
rect 38508 14084 38564 14140
rect 38612 14084 38668 14140
rect 38716 14084 38772 14140
rect 5874 13076 5930 13132
rect 5978 13076 6034 13132
rect 6082 13076 6138 13132
rect 15198 13076 15254 13132
rect 15302 13076 15358 13132
rect 15406 13076 15462 13132
rect 24522 13076 24578 13132
rect 24626 13076 24682 13132
rect 24730 13076 24786 13132
rect 33846 13076 33902 13132
rect 33950 13076 34006 13132
rect 34054 13076 34110 13132
rect 10536 12068 10592 12124
rect 10640 12068 10696 12124
rect 10744 12068 10800 12124
rect 19860 12068 19916 12124
rect 19964 12068 20020 12124
rect 20068 12068 20124 12124
rect 29184 12068 29240 12124
rect 29288 12068 29344 12124
rect 29392 12068 29448 12124
rect 38508 12068 38564 12124
rect 38612 12068 38668 12124
rect 38716 12068 38772 12124
rect 5874 11060 5930 11116
rect 5978 11060 6034 11116
rect 6082 11060 6138 11116
rect 15198 11060 15254 11116
rect 15302 11060 15358 11116
rect 15406 11060 15462 11116
rect 24522 11060 24578 11116
rect 24626 11060 24682 11116
rect 24730 11060 24786 11116
rect 33846 11060 33902 11116
rect 33950 11060 34006 11116
rect 34054 11060 34110 11116
rect 10536 10052 10592 10108
rect 10640 10052 10696 10108
rect 10744 10052 10800 10108
rect 19860 10052 19916 10108
rect 19964 10052 20020 10108
rect 20068 10052 20124 10108
rect 29184 10052 29240 10108
rect 29288 10052 29344 10108
rect 29392 10052 29448 10108
rect 38508 10052 38564 10108
rect 38612 10052 38668 10108
rect 38716 10052 38772 10108
rect 5874 9044 5930 9100
rect 5978 9044 6034 9100
rect 6082 9044 6138 9100
rect 15198 9044 15254 9100
rect 15302 9044 15358 9100
rect 15406 9044 15462 9100
rect 24522 9044 24578 9100
rect 24626 9044 24682 9100
rect 24730 9044 24786 9100
rect 33846 9044 33902 9100
rect 33950 9044 34006 9100
rect 34054 9044 34110 9100
rect 10536 8036 10592 8092
rect 10640 8036 10696 8092
rect 10744 8036 10800 8092
rect 19860 8036 19916 8092
rect 19964 8036 20020 8092
rect 20068 8036 20124 8092
rect 29184 8036 29240 8092
rect 29288 8036 29344 8092
rect 29392 8036 29448 8092
rect 38508 8036 38564 8092
rect 38612 8036 38668 8092
rect 38716 8036 38772 8092
rect 5874 7028 5930 7084
rect 5978 7028 6034 7084
rect 6082 7028 6138 7084
rect 15198 7028 15254 7084
rect 15302 7028 15358 7084
rect 15406 7028 15462 7084
rect 24522 7028 24578 7084
rect 24626 7028 24682 7084
rect 24730 7028 24786 7084
rect 33846 7028 33902 7084
rect 33950 7028 34006 7084
rect 34054 7028 34110 7084
rect 10536 6020 10592 6076
rect 10640 6020 10696 6076
rect 10744 6020 10800 6076
rect 19860 6020 19916 6076
rect 19964 6020 20020 6076
rect 20068 6020 20124 6076
rect 29184 6020 29240 6076
rect 29288 6020 29344 6076
rect 29392 6020 29448 6076
rect 38508 6020 38564 6076
rect 38612 6020 38668 6076
rect 38716 6020 38772 6076
rect 5874 5012 5930 5068
rect 5978 5012 6034 5068
rect 6082 5012 6138 5068
rect 15198 5012 15254 5068
rect 15302 5012 15358 5068
rect 15406 5012 15462 5068
rect 24522 5012 24578 5068
rect 24626 5012 24682 5068
rect 24730 5012 24786 5068
rect 33846 5012 33902 5068
rect 33950 5012 34006 5068
rect 34054 5012 34110 5068
rect 10536 4004 10592 4060
rect 10640 4004 10696 4060
rect 10744 4004 10800 4060
rect 19860 4004 19916 4060
rect 19964 4004 20020 4060
rect 20068 4004 20124 4060
rect 29184 4004 29240 4060
rect 29288 4004 29344 4060
rect 29392 4004 29448 4060
rect 38508 4004 38564 4060
rect 38612 4004 38668 4060
rect 38716 4004 38772 4060
<< metal4 >>
rect 5846 35308 6166 36348
rect 5846 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6166 35308
rect 5846 33292 6166 35252
rect 5846 33236 5874 33292
rect 5930 33236 5978 33292
rect 6034 33236 6082 33292
rect 6138 33236 6166 33292
rect 5846 31276 6166 33236
rect 5846 31220 5874 31276
rect 5930 31220 5978 31276
rect 6034 31220 6082 31276
rect 6138 31220 6166 31276
rect 5846 29260 6166 31220
rect 5846 29204 5874 29260
rect 5930 29204 5978 29260
rect 6034 29204 6082 29260
rect 6138 29204 6166 29260
rect 5846 27244 6166 29204
rect 5846 27188 5874 27244
rect 5930 27188 5978 27244
rect 6034 27188 6082 27244
rect 6138 27188 6166 27244
rect 5846 25228 6166 27188
rect 5846 25172 5874 25228
rect 5930 25172 5978 25228
rect 6034 25172 6082 25228
rect 6138 25172 6166 25228
rect 5846 23212 6166 25172
rect 5846 23156 5874 23212
rect 5930 23156 5978 23212
rect 6034 23156 6082 23212
rect 6138 23156 6166 23212
rect 5846 21196 6166 23156
rect 5846 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6166 21196
rect 5846 19180 6166 21140
rect 5846 19124 5874 19180
rect 5930 19124 5978 19180
rect 6034 19124 6082 19180
rect 6138 19124 6166 19180
rect 5846 17164 6166 19124
rect 5846 17108 5874 17164
rect 5930 17108 5978 17164
rect 6034 17108 6082 17164
rect 6138 17108 6166 17164
rect 5846 15148 6166 17108
rect 5846 15092 5874 15148
rect 5930 15092 5978 15148
rect 6034 15092 6082 15148
rect 6138 15092 6166 15148
rect 5846 13132 6166 15092
rect 5846 13076 5874 13132
rect 5930 13076 5978 13132
rect 6034 13076 6082 13132
rect 6138 13076 6166 13132
rect 5846 11116 6166 13076
rect 5846 11060 5874 11116
rect 5930 11060 5978 11116
rect 6034 11060 6082 11116
rect 6138 11060 6166 11116
rect 5846 9100 6166 11060
rect 5846 9044 5874 9100
rect 5930 9044 5978 9100
rect 6034 9044 6082 9100
rect 6138 9044 6166 9100
rect 5846 7084 6166 9044
rect 5846 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6166 7084
rect 5846 5068 6166 7028
rect 5846 5012 5874 5068
rect 5930 5012 5978 5068
rect 6034 5012 6082 5068
rect 6138 5012 6166 5068
rect 5846 3972 6166 5012
rect 10508 36316 10828 36348
rect 10508 36260 10536 36316
rect 10592 36260 10640 36316
rect 10696 36260 10744 36316
rect 10800 36260 10828 36316
rect 10508 34300 10828 36260
rect 10508 34244 10536 34300
rect 10592 34244 10640 34300
rect 10696 34244 10744 34300
rect 10800 34244 10828 34300
rect 10508 32284 10828 34244
rect 10508 32228 10536 32284
rect 10592 32228 10640 32284
rect 10696 32228 10744 32284
rect 10800 32228 10828 32284
rect 10508 30268 10828 32228
rect 10508 30212 10536 30268
rect 10592 30212 10640 30268
rect 10696 30212 10744 30268
rect 10800 30212 10828 30268
rect 10508 28252 10828 30212
rect 10508 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10828 28252
rect 10508 26236 10828 28196
rect 10508 26180 10536 26236
rect 10592 26180 10640 26236
rect 10696 26180 10744 26236
rect 10800 26180 10828 26236
rect 10508 24220 10828 26180
rect 10508 24164 10536 24220
rect 10592 24164 10640 24220
rect 10696 24164 10744 24220
rect 10800 24164 10828 24220
rect 10508 22204 10828 24164
rect 10508 22148 10536 22204
rect 10592 22148 10640 22204
rect 10696 22148 10744 22204
rect 10800 22148 10828 22204
rect 10508 20188 10828 22148
rect 10508 20132 10536 20188
rect 10592 20132 10640 20188
rect 10696 20132 10744 20188
rect 10800 20132 10828 20188
rect 10508 18172 10828 20132
rect 10508 18116 10536 18172
rect 10592 18116 10640 18172
rect 10696 18116 10744 18172
rect 10800 18116 10828 18172
rect 10508 16156 10828 18116
rect 10508 16100 10536 16156
rect 10592 16100 10640 16156
rect 10696 16100 10744 16156
rect 10800 16100 10828 16156
rect 10508 14140 10828 16100
rect 10508 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10828 14140
rect 10508 12124 10828 14084
rect 10508 12068 10536 12124
rect 10592 12068 10640 12124
rect 10696 12068 10744 12124
rect 10800 12068 10828 12124
rect 10508 10108 10828 12068
rect 10508 10052 10536 10108
rect 10592 10052 10640 10108
rect 10696 10052 10744 10108
rect 10800 10052 10828 10108
rect 10508 8092 10828 10052
rect 10508 8036 10536 8092
rect 10592 8036 10640 8092
rect 10696 8036 10744 8092
rect 10800 8036 10828 8092
rect 10508 6076 10828 8036
rect 10508 6020 10536 6076
rect 10592 6020 10640 6076
rect 10696 6020 10744 6076
rect 10800 6020 10828 6076
rect 10508 4060 10828 6020
rect 10508 4004 10536 4060
rect 10592 4004 10640 4060
rect 10696 4004 10744 4060
rect 10800 4004 10828 4060
rect 10508 3972 10828 4004
rect 15170 35308 15490 36348
rect 15170 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15490 35308
rect 15170 33292 15490 35252
rect 15170 33236 15198 33292
rect 15254 33236 15302 33292
rect 15358 33236 15406 33292
rect 15462 33236 15490 33292
rect 15170 31276 15490 33236
rect 15170 31220 15198 31276
rect 15254 31220 15302 31276
rect 15358 31220 15406 31276
rect 15462 31220 15490 31276
rect 15170 29260 15490 31220
rect 15170 29204 15198 29260
rect 15254 29204 15302 29260
rect 15358 29204 15406 29260
rect 15462 29204 15490 29260
rect 15170 27244 15490 29204
rect 15170 27188 15198 27244
rect 15254 27188 15302 27244
rect 15358 27188 15406 27244
rect 15462 27188 15490 27244
rect 15170 25228 15490 27188
rect 15170 25172 15198 25228
rect 15254 25172 15302 25228
rect 15358 25172 15406 25228
rect 15462 25172 15490 25228
rect 15170 23212 15490 25172
rect 15170 23156 15198 23212
rect 15254 23156 15302 23212
rect 15358 23156 15406 23212
rect 15462 23156 15490 23212
rect 15170 21196 15490 23156
rect 15170 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15490 21196
rect 15170 19180 15490 21140
rect 15170 19124 15198 19180
rect 15254 19124 15302 19180
rect 15358 19124 15406 19180
rect 15462 19124 15490 19180
rect 15170 17164 15490 19124
rect 15170 17108 15198 17164
rect 15254 17108 15302 17164
rect 15358 17108 15406 17164
rect 15462 17108 15490 17164
rect 15170 15148 15490 17108
rect 15170 15092 15198 15148
rect 15254 15092 15302 15148
rect 15358 15092 15406 15148
rect 15462 15092 15490 15148
rect 15170 13132 15490 15092
rect 15170 13076 15198 13132
rect 15254 13076 15302 13132
rect 15358 13076 15406 13132
rect 15462 13076 15490 13132
rect 15170 11116 15490 13076
rect 15170 11060 15198 11116
rect 15254 11060 15302 11116
rect 15358 11060 15406 11116
rect 15462 11060 15490 11116
rect 15170 9100 15490 11060
rect 15170 9044 15198 9100
rect 15254 9044 15302 9100
rect 15358 9044 15406 9100
rect 15462 9044 15490 9100
rect 15170 7084 15490 9044
rect 15170 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15490 7084
rect 15170 5068 15490 7028
rect 15170 5012 15198 5068
rect 15254 5012 15302 5068
rect 15358 5012 15406 5068
rect 15462 5012 15490 5068
rect 15170 3972 15490 5012
rect 19832 36316 20152 36348
rect 19832 36260 19860 36316
rect 19916 36260 19964 36316
rect 20020 36260 20068 36316
rect 20124 36260 20152 36316
rect 19832 34300 20152 36260
rect 19832 34244 19860 34300
rect 19916 34244 19964 34300
rect 20020 34244 20068 34300
rect 20124 34244 20152 34300
rect 19832 32284 20152 34244
rect 19832 32228 19860 32284
rect 19916 32228 19964 32284
rect 20020 32228 20068 32284
rect 20124 32228 20152 32284
rect 19832 30268 20152 32228
rect 19832 30212 19860 30268
rect 19916 30212 19964 30268
rect 20020 30212 20068 30268
rect 20124 30212 20152 30268
rect 19832 28252 20152 30212
rect 19832 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20152 28252
rect 19832 26236 20152 28196
rect 19832 26180 19860 26236
rect 19916 26180 19964 26236
rect 20020 26180 20068 26236
rect 20124 26180 20152 26236
rect 19832 24220 20152 26180
rect 19832 24164 19860 24220
rect 19916 24164 19964 24220
rect 20020 24164 20068 24220
rect 20124 24164 20152 24220
rect 19832 22204 20152 24164
rect 19832 22148 19860 22204
rect 19916 22148 19964 22204
rect 20020 22148 20068 22204
rect 20124 22148 20152 22204
rect 19832 20188 20152 22148
rect 19832 20132 19860 20188
rect 19916 20132 19964 20188
rect 20020 20132 20068 20188
rect 20124 20132 20152 20188
rect 19832 18172 20152 20132
rect 19832 18116 19860 18172
rect 19916 18116 19964 18172
rect 20020 18116 20068 18172
rect 20124 18116 20152 18172
rect 19832 16156 20152 18116
rect 19832 16100 19860 16156
rect 19916 16100 19964 16156
rect 20020 16100 20068 16156
rect 20124 16100 20152 16156
rect 19832 14140 20152 16100
rect 19832 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20152 14140
rect 19832 12124 20152 14084
rect 19832 12068 19860 12124
rect 19916 12068 19964 12124
rect 20020 12068 20068 12124
rect 20124 12068 20152 12124
rect 19832 10108 20152 12068
rect 19832 10052 19860 10108
rect 19916 10052 19964 10108
rect 20020 10052 20068 10108
rect 20124 10052 20152 10108
rect 19832 8092 20152 10052
rect 19832 8036 19860 8092
rect 19916 8036 19964 8092
rect 20020 8036 20068 8092
rect 20124 8036 20152 8092
rect 19832 6076 20152 8036
rect 19832 6020 19860 6076
rect 19916 6020 19964 6076
rect 20020 6020 20068 6076
rect 20124 6020 20152 6076
rect 19832 4060 20152 6020
rect 19832 4004 19860 4060
rect 19916 4004 19964 4060
rect 20020 4004 20068 4060
rect 20124 4004 20152 4060
rect 19832 3972 20152 4004
rect 24494 35308 24814 36348
rect 24494 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24814 35308
rect 24494 33292 24814 35252
rect 24494 33236 24522 33292
rect 24578 33236 24626 33292
rect 24682 33236 24730 33292
rect 24786 33236 24814 33292
rect 24494 31276 24814 33236
rect 24494 31220 24522 31276
rect 24578 31220 24626 31276
rect 24682 31220 24730 31276
rect 24786 31220 24814 31276
rect 24494 29260 24814 31220
rect 24494 29204 24522 29260
rect 24578 29204 24626 29260
rect 24682 29204 24730 29260
rect 24786 29204 24814 29260
rect 24494 27244 24814 29204
rect 24494 27188 24522 27244
rect 24578 27188 24626 27244
rect 24682 27188 24730 27244
rect 24786 27188 24814 27244
rect 24494 25228 24814 27188
rect 24494 25172 24522 25228
rect 24578 25172 24626 25228
rect 24682 25172 24730 25228
rect 24786 25172 24814 25228
rect 24494 23212 24814 25172
rect 24494 23156 24522 23212
rect 24578 23156 24626 23212
rect 24682 23156 24730 23212
rect 24786 23156 24814 23212
rect 24494 21196 24814 23156
rect 24494 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24814 21196
rect 24494 19180 24814 21140
rect 24494 19124 24522 19180
rect 24578 19124 24626 19180
rect 24682 19124 24730 19180
rect 24786 19124 24814 19180
rect 24494 17164 24814 19124
rect 24494 17108 24522 17164
rect 24578 17108 24626 17164
rect 24682 17108 24730 17164
rect 24786 17108 24814 17164
rect 24494 15148 24814 17108
rect 24494 15092 24522 15148
rect 24578 15092 24626 15148
rect 24682 15092 24730 15148
rect 24786 15092 24814 15148
rect 24494 13132 24814 15092
rect 24494 13076 24522 13132
rect 24578 13076 24626 13132
rect 24682 13076 24730 13132
rect 24786 13076 24814 13132
rect 24494 11116 24814 13076
rect 24494 11060 24522 11116
rect 24578 11060 24626 11116
rect 24682 11060 24730 11116
rect 24786 11060 24814 11116
rect 24494 9100 24814 11060
rect 24494 9044 24522 9100
rect 24578 9044 24626 9100
rect 24682 9044 24730 9100
rect 24786 9044 24814 9100
rect 24494 7084 24814 9044
rect 24494 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24814 7084
rect 24494 5068 24814 7028
rect 24494 5012 24522 5068
rect 24578 5012 24626 5068
rect 24682 5012 24730 5068
rect 24786 5012 24814 5068
rect 24494 3972 24814 5012
rect 29156 36316 29476 36348
rect 29156 36260 29184 36316
rect 29240 36260 29288 36316
rect 29344 36260 29392 36316
rect 29448 36260 29476 36316
rect 29156 34300 29476 36260
rect 29156 34244 29184 34300
rect 29240 34244 29288 34300
rect 29344 34244 29392 34300
rect 29448 34244 29476 34300
rect 29156 32284 29476 34244
rect 29156 32228 29184 32284
rect 29240 32228 29288 32284
rect 29344 32228 29392 32284
rect 29448 32228 29476 32284
rect 29156 30268 29476 32228
rect 29156 30212 29184 30268
rect 29240 30212 29288 30268
rect 29344 30212 29392 30268
rect 29448 30212 29476 30268
rect 29156 28252 29476 30212
rect 29156 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29476 28252
rect 29156 26236 29476 28196
rect 29156 26180 29184 26236
rect 29240 26180 29288 26236
rect 29344 26180 29392 26236
rect 29448 26180 29476 26236
rect 29156 24220 29476 26180
rect 29156 24164 29184 24220
rect 29240 24164 29288 24220
rect 29344 24164 29392 24220
rect 29448 24164 29476 24220
rect 29156 22204 29476 24164
rect 29156 22148 29184 22204
rect 29240 22148 29288 22204
rect 29344 22148 29392 22204
rect 29448 22148 29476 22204
rect 29156 20188 29476 22148
rect 29156 20132 29184 20188
rect 29240 20132 29288 20188
rect 29344 20132 29392 20188
rect 29448 20132 29476 20188
rect 29156 18172 29476 20132
rect 29156 18116 29184 18172
rect 29240 18116 29288 18172
rect 29344 18116 29392 18172
rect 29448 18116 29476 18172
rect 29156 16156 29476 18116
rect 29156 16100 29184 16156
rect 29240 16100 29288 16156
rect 29344 16100 29392 16156
rect 29448 16100 29476 16156
rect 29156 14140 29476 16100
rect 29156 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29476 14140
rect 29156 12124 29476 14084
rect 29156 12068 29184 12124
rect 29240 12068 29288 12124
rect 29344 12068 29392 12124
rect 29448 12068 29476 12124
rect 29156 10108 29476 12068
rect 29156 10052 29184 10108
rect 29240 10052 29288 10108
rect 29344 10052 29392 10108
rect 29448 10052 29476 10108
rect 29156 8092 29476 10052
rect 29156 8036 29184 8092
rect 29240 8036 29288 8092
rect 29344 8036 29392 8092
rect 29448 8036 29476 8092
rect 29156 6076 29476 8036
rect 29156 6020 29184 6076
rect 29240 6020 29288 6076
rect 29344 6020 29392 6076
rect 29448 6020 29476 6076
rect 29156 4060 29476 6020
rect 29156 4004 29184 4060
rect 29240 4004 29288 4060
rect 29344 4004 29392 4060
rect 29448 4004 29476 4060
rect 29156 3972 29476 4004
rect 33818 35308 34138 36348
rect 33818 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34138 35308
rect 33818 33292 34138 35252
rect 33818 33236 33846 33292
rect 33902 33236 33950 33292
rect 34006 33236 34054 33292
rect 34110 33236 34138 33292
rect 33818 31276 34138 33236
rect 33818 31220 33846 31276
rect 33902 31220 33950 31276
rect 34006 31220 34054 31276
rect 34110 31220 34138 31276
rect 33818 29260 34138 31220
rect 33818 29204 33846 29260
rect 33902 29204 33950 29260
rect 34006 29204 34054 29260
rect 34110 29204 34138 29260
rect 33818 27244 34138 29204
rect 33818 27188 33846 27244
rect 33902 27188 33950 27244
rect 34006 27188 34054 27244
rect 34110 27188 34138 27244
rect 33818 25228 34138 27188
rect 33818 25172 33846 25228
rect 33902 25172 33950 25228
rect 34006 25172 34054 25228
rect 34110 25172 34138 25228
rect 33818 23212 34138 25172
rect 33818 23156 33846 23212
rect 33902 23156 33950 23212
rect 34006 23156 34054 23212
rect 34110 23156 34138 23212
rect 33818 21196 34138 23156
rect 33818 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34138 21196
rect 33818 19180 34138 21140
rect 33818 19124 33846 19180
rect 33902 19124 33950 19180
rect 34006 19124 34054 19180
rect 34110 19124 34138 19180
rect 33818 17164 34138 19124
rect 33818 17108 33846 17164
rect 33902 17108 33950 17164
rect 34006 17108 34054 17164
rect 34110 17108 34138 17164
rect 33818 15148 34138 17108
rect 33818 15092 33846 15148
rect 33902 15092 33950 15148
rect 34006 15092 34054 15148
rect 34110 15092 34138 15148
rect 33818 13132 34138 15092
rect 33818 13076 33846 13132
rect 33902 13076 33950 13132
rect 34006 13076 34054 13132
rect 34110 13076 34138 13132
rect 33818 11116 34138 13076
rect 33818 11060 33846 11116
rect 33902 11060 33950 11116
rect 34006 11060 34054 11116
rect 34110 11060 34138 11116
rect 33818 9100 34138 11060
rect 33818 9044 33846 9100
rect 33902 9044 33950 9100
rect 34006 9044 34054 9100
rect 34110 9044 34138 9100
rect 33818 7084 34138 9044
rect 33818 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34138 7084
rect 33818 5068 34138 7028
rect 33818 5012 33846 5068
rect 33902 5012 33950 5068
rect 34006 5012 34054 5068
rect 34110 5012 34138 5068
rect 33818 3972 34138 5012
rect 38480 36316 38800 36348
rect 38480 36260 38508 36316
rect 38564 36260 38612 36316
rect 38668 36260 38716 36316
rect 38772 36260 38800 36316
rect 38480 34300 38800 36260
rect 38480 34244 38508 34300
rect 38564 34244 38612 34300
rect 38668 34244 38716 34300
rect 38772 34244 38800 34300
rect 38480 32284 38800 34244
rect 38480 32228 38508 32284
rect 38564 32228 38612 32284
rect 38668 32228 38716 32284
rect 38772 32228 38800 32284
rect 38480 30268 38800 32228
rect 38480 30212 38508 30268
rect 38564 30212 38612 30268
rect 38668 30212 38716 30268
rect 38772 30212 38800 30268
rect 38480 28252 38800 30212
rect 38480 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38800 28252
rect 38480 26236 38800 28196
rect 38480 26180 38508 26236
rect 38564 26180 38612 26236
rect 38668 26180 38716 26236
rect 38772 26180 38800 26236
rect 38480 24220 38800 26180
rect 38480 24164 38508 24220
rect 38564 24164 38612 24220
rect 38668 24164 38716 24220
rect 38772 24164 38800 24220
rect 38480 22204 38800 24164
rect 38480 22148 38508 22204
rect 38564 22148 38612 22204
rect 38668 22148 38716 22204
rect 38772 22148 38800 22204
rect 38480 20188 38800 22148
rect 38480 20132 38508 20188
rect 38564 20132 38612 20188
rect 38668 20132 38716 20188
rect 38772 20132 38800 20188
rect 38480 18172 38800 20132
rect 38480 18116 38508 18172
rect 38564 18116 38612 18172
rect 38668 18116 38716 18172
rect 38772 18116 38800 18172
rect 38480 16156 38800 18116
rect 38480 16100 38508 16156
rect 38564 16100 38612 16156
rect 38668 16100 38716 16156
rect 38772 16100 38800 16156
rect 38480 14140 38800 16100
rect 38480 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38800 14140
rect 38480 12124 38800 14084
rect 38480 12068 38508 12124
rect 38564 12068 38612 12124
rect 38668 12068 38716 12124
rect 38772 12068 38800 12124
rect 38480 10108 38800 12068
rect 38480 10052 38508 10108
rect 38564 10052 38612 10108
rect 38668 10052 38716 10108
rect 38772 10052 38800 10108
rect 38480 8092 38800 10052
rect 38480 8036 38508 8092
rect 38564 8036 38612 8092
rect 38668 8036 38716 8092
rect 38772 8036 38800 8092
rect 38480 6076 38800 8036
rect 38480 6020 38508 6076
rect 38564 6020 38612 6076
rect 38668 6020 38716 6076
rect 38772 6020 38800 6076
rect 38480 4060 38800 6020
rect 38480 4004 38508 4060
rect 38564 4004 38612 4060
rect 38668 4004 38716 4060
rect 38772 4004 38800 4060
rect 38480 3972 38800 4004
use gf180mcu_fd_sc_mcu9t5v0__xnor2_1  _11_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 11760 0 1 18144
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor2_1  _12_
timestamp 1698431365
transform -1 0 14672 0 1 20160
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__xor2_1  _13_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 14896 0 1 18144
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor3_1  _14_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 11872 0 -1 20160
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor2_1  _15_
timestamp 1698431365
transform -1 0 17808 0 1 18144
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor3_1  _16_
timestamp 1698431365
transform 1 0 14448 0 -1 20160
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  _17_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 19600 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor2_1  _18_
timestamp 1698431365
transform -1 0 19152 0 1 20160
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__xnor3_1  _19_
timestamp 1698431365
transform 1 0 17696 0 -1 20160
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _20_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 20272 0 1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__xor2_1  _21_
timestamp 1698431365
transform 1 0 21168 0 1 20160
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__xor3_1  _22_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform -1 0 23184 0 -1 20160
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _23_
timestamp 1698431365
transform 1 0 23296 0 1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__xor2_1  _24_
timestamp 1698431365
transform 1 0 23520 0 -1 20160
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__xor3_1  _25_
timestamp 1698431365
transform 1 0 23184 0 1 18144
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _26_
timestamp 1698431365
transform 1 0 25984 0 1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__xor2_1  _27_
timestamp 1698431365
transform 1 0 26320 0 1 18144
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__xor3_1  _28_
timestamp 1698431365
transform 1 0 26096 0 -1 20160
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _29_
timestamp 1698431365
transform 1 0 29008 0 1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__xor2_1  _30_
timestamp 1698431365
transform 1 0 29008 0 1 18144
box -86 -90 1430 1098
use gf180mcu_fd_sc_mcu9t5v0__xor3_1  _31_
timestamp 1698431365
transform -1 0 31248 0 -1 20160
box -86 -90 2662 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _32_
timestamp 1698431365
transform 1 0 30576 0 1 20160
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__buf_1  _33_
timestamp 1698431365
transform 1 0 15008 0 -1 32256
box -86 -90 758 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__11__A1 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 11536 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__11__A2
timestamp 1698431365
transform 1 0 11088 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__12__A1
timestamp 1698431365
transform 1 0 12880 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__12__A2
timestamp 1698431365
transform 1 0 12432 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__13__A1
timestamp 1698431365
transform -1 0 13552 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__13__A2
timestamp 1698431365
transform -1 0 14000 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__15__A1
timestamp 1698431365
transform 1 0 16240 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__15__A2
timestamp 1698431365
transform -1 0 16016 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__16__A1
timestamp 1698431365
transform 1 0 14896 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__18__A1
timestamp 1698431365
transform 1 0 17584 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__19__A1
timestamp 1698431365
transform -1 0 17696 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__19__A2
timestamp 1698431365
transform -1 0 18256 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__21__A1
timestamp 1698431365
transform -1 0 22960 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__22__A1
timestamp 1698431365
transform -1 0 24416 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__22__A2
timestamp 1698431365
transform 1 0 25312 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__24__A1
timestamp 1698431365
transform 1 0 25760 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__25__A1
timestamp 1698431365
transform 1 0 25984 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__25__A2
timestamp 1698431365
transform 1 0 25984 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__27__A1
timestamp 1698431365
transform 1 0 27888 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__28__A1
timestamp 1698431365
transform 1 0 28560 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__28__A2
timestamp 1698431365
transform -1 0 30128 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__30__A1
timestamp 1698431365
transform 1 0 30576 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__31__A1
timestamp 1698431365
transform 1 0 31472 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__31__A2
timestamp 1698431365
transform 1 0 31920 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__antenna  ANTENNA__33__I
timestamp 1698431365
transform -1 0 15008 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 4032
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_0_308 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 35840 0 1 4032
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_0_324 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 37632 0 1 4032
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_0_328 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 38080 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_0_330 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 38304 0 1 4032
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 6048
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_1_314
timestamp 1698431365
transform 1 0 36512 0 -1 6048
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_1_330
timestamp 1698431365
transform 1 0 38304 0 -1 6048
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 6048
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 6048
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 6048
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_2_317 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 6048
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_2_325
timestamp 1698431365
transform 1 0 37744 0 1 6048
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_2_329
timestamp 1698431365
transform 1 0 38192 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 8064
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_3_314
timestamp 1698431365
transform 1 0 36512 0 -1 8064
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_3_330
timestamp 1698431365
transform 1 0 38304 0 -1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 8064
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 8064
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 8064
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 8064
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_4_325
timestamp 1698431365
transform 1 0 37744 0 1 8064
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_4_329
timestamp 1698431365
transform 1 0 38192 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_5_314
timestamp 1698431365
transform 1 0 36512 0 -1 10080
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_5_330
timestamp 1698431365
transform 1 0 38304 0 -1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 10080
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 10080
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 10080
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 10080
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_6_325
timestamp 1698431365
transform 1 0 37744 0 1 10080
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_6_329
timestamp 1698431365
transform 1 0 38192 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 12096
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_7_314
timestamp 1698431365
transform 1 0 36512 0 -1 12096
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_7_330
timestamp 1698431365
transform 1 0 38304 0 -1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 12096
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 12096
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 12096
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 12096
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 12096
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_8_329
timestamp 1698431365
transform 1 0 38192 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_9_314
timestamp 1698431365
transform 1 0 36512 0 -1 14112
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_9_330
timestamp 1698431365
transform 1 0 38304 0 -1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_10_325
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_10_329
timestamp 1698431365
transform 1 0 38192 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 16128
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_11_314
timestamp 1698431365
transform 1 0 36512 0 -1 16128
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_11_330
timestamp 1698431365
transform 1 0 38304 0 -1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 16128
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 16128
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 16128
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 16128
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_12_325
timestamp 1698431365
transform 1 0 37744 0 1 16128
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_12_329
timestamp 1698431365
transform 1 0 38192 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 18144
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 18144
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_104
timestamp 1698431365
transform 1 0 12992 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_106
timestamp 1698431365
transform 1 0 13216 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_109
timestamp 1698431365
transform 1 0 13552 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_13_113
timestamp 1698431365
transform 1 0 14000 0 -1 18144
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_13_129
timestamp 1698431365
transform 1 0 15792 0 -1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_137
timestamp 1698431365
transform 1 0 16688 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 18144
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_13_222
timestamp 1698431365
transform 1 0 26208 0 -1 18144
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_13_254
timestamp 1698431365
transform 1 0 29792 0 -1 18144
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_13_270
timestamp 1698431365
transform 1 0 31584 0 -1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_13_278
timestamp 1698431365
transform 1 0 32480 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 18144
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_13_314
timestamp 1698431365
transform 1 0 36512 0 -1 18144
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_13_330
timestamp 1698431365
transform 1 0 38304 0 -1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 18144
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 18144
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_14_69
timestamp 1698431365
transform 1 0 9072 0 1 18144
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_85
timestamp 1698431365
transform 1 0 10864 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_89
timestamp 1698431365
transform 1 0 11312 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_14_121
timestamp 1698431365
transform 1 0 14896 0 1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_131
timestamp 1698431365
transform 1 0 16016 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_147
timestamp 1698431365
transform 1 0 17808 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_14_151
timestamp 1698431365
transform 1 0 18256 0 1 18144
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_14_167
timestamp 1698431365
transform 1 0 20048 0 1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 18144
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_193
timestamp 1698431365
transform 1 0 22960 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_218
timestamp 1698431365
transform 1 0 25760 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_14_222
timestamp 1698431365
transform 1 0 26208 0 1 18144
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_235
timestamp 1698431365
transform 1 0 27664 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698431365
transform 1 0 28112 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_259
timestamp 1698431365
transform 1 0 30352 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_14_263
timestamp 1698431365
transform 1 0 30800 0 1 18144
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_14_295
timestamp 1698431365
transform 1 0 34384 0 1 18144
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 18144
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_14_325
timestamp 1698431365
transform 1 0 37744 0 1 18144
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_14_329
timestamp 1698431365
transform 1 0 38192 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 20160
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 20160
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_88
timestamp 1698431365
transform 1 0 11200 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_92
timestamp 1698431365
transform 1 0 11648 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_169
timestamp 1698431365
transform 1 0 20272 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_171
timestamp 1698431365
transform 1 0 20496 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_195
timestamp 1698431365
transform 1 0 23184 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_197
timestamp 1698431365
transform 1 0 23408 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_220
timestamp 1698431365
transform 1 0 25984 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_267
timestamp 1698431365
transform 1 0 31248 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_15_271
timestamp 1698431365
transform 1 0 31696 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_15_275
timestamp 1698431365
transform 1 0 32144 0 -1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 20160
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_15_314
timestamp 1698431365
transform 1 0 36512 0 -1 20160
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_15_330
timestamp 1698431365
transform 1 0 38304 0 -1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 20160
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 20160
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_16_69
timestamp 1698431365
transform 1 0 9072 0 1 20160
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_16_85
timestamp 1698431365
transform 1 0 10864 0 1 20160
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_93
timestamp 1698431365
transform 1 0 11760 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_97
timestamp 1698431365
transform 1 0 12208 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_119
timestamp 1698431365
transform 1 0 14672 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_16_123
timestamp 1698431365
transform 1 0 15120 0 1 20160
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_139
timestamp 1698431365
transform 1 0 16912 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_143
timestamp 1698431365
transform 1 0 17360 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_163
timestamp 1698431365
transform 1 0 19600 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_167
timestamp 1698431365
transform 1 0 20048 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_189
timestamp 1698431365
transform 1 0 22512 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_193
timestamp 1698431365
transform 1 0 22960 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_195
timestamp 1698431365
transform 1 0 23184 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_202
timestamp 1698431365
transform 1 0 23968 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_16_206
timestamp 1698431365
transform 1 0 24416 0 1 20160
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_214
timestamp 1698431365
transform 1 0 25312 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_218
timestamp 1698431365
transform 1 0 25760 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_16_226
timestamp 1698431365
transform 1 0 26656 0 1 20160
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_242
timestamp 1698431365
transform 1 0 28448 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 20160
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_253
timestamp 1698431365
transform 1 0 29680 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_257
timestamp 1698431365
transform 1 0 30128 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_16_267
timestamp 1698431365
transform 1 0 31248 0 1 20160
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_16_299
timestamp 1698431365
transform 1 0 34832 0 1 20160
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 20160
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_16_325
timestamp 1698431365
transform 1 0 37744 0 1 20160
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_16_329
timestamp 1698431365
transform 1 0 38192 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 22176
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 22176
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 22176
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698431365
transform 1 0 24416 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 22176
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698431365
transform 1 0 32256 0 -1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 22176
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_17_314
timestamp 1698431365
transform 1 0 36512 0 -1 22176
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_17_330
timestamp 1698431365
transform 1 0 38304 0 -1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 22176
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 22176
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 22176
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 22176
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 22176
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698431365
transform 1 0 28336 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 22176
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 22176
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_18_325
timestamp 1698431365
transform 1 0 37744 0 1 22176
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_18_329
timestamp 1698431365
transform 1 0 38192 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 24192
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 24192
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698431365
transform 1 0 16576 0 -1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 24192
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698431365
transform 1 0 24416 0 -1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 24192
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 24192
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_19_314
timestamp 1698431365
transform 1 0 36512 0 -1 24192
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_19_330
timestamp 1698431365
transform 1 0 38304 0 -1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 24192
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 24192
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 24192
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 24192
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 24192
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 24192
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698431365
transform 1 0 36176 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 24192
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_20_325
timestamp 1698431365
transform 1 0 37744 0 1 24192
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_20_329
timestamp 1698431365
transform 1 0 38192 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 26208
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 26208
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 26208
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 26208
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 26208
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_21_314
timestamp 1698431365
transform 1 0 36512 0 -1 26208
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_21_330
timestamp 1698431365
transform 1 0 38304 0 -1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 26208
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 26208
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 26208
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 26208
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 26208
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 26208
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 26208
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_22_325
timestamp 1698431365
transform 1 0 37744 0 1 26208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_22_329
timestamp 1698431365
transform 1 0 38192 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_23_314
timestamp 1698431365
transform 1 0 36512 0 -1 28224
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_23_330
timestamp 1698431365
transform 1 0 38304 0 -1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_24_325
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_24_329
timestamp 1698431365
transform 1 0 38192 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 30240
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698431365
transform 1 0 8736 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 30240
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 30240
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698431365
transform 1 0 24416 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 30240
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 30240
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_25_314
timestamp 1698431365
transform 1 0 36512 0 -1 30240
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_25_330
timestamp 1698431365
transform 1 0 38304 0 -1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 30240
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 30240
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 30240
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 30240
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 30240
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698431365
transform 1 0 28336 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 30240
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 30240
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_26_325
timestamp 1698431365
transform 1 0 37744 0 1 30240
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_26_329
timestamp 1698431365
transform 1 0 38192 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 32256
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 32256
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_27_104
timestamp 1698431365
transform 1 0 12992 0 -1 32256
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_27_128
timestamp 1698431365
transform 1 0 15680 0 -1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 32256
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 32256
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 32256
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_27_314
timestamp 1698431365
transform 1 0 36512 0 -1 32256
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_27_330
timestamp 1698431365
transform 1 0 38304 0 -1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 32256
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 32256
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 32256
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 32256
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 32256
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 32256
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698431365
transform 1 0 36176 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 32256
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_28_325
timestamp 1698431365
transform 1 0 37744 0 1 32256
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_28_329
timestamp 1698431365
transform 1 0 38192 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 34272
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698431365
transform 1 0 8736 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 34272
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 34272
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 34272
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 34272
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_29_314
timestamp 1698431365
transform 1 0 36512 0 -1 34272
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_29_330
timestamp 1698431365
transform 1 0 38304 0 -1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 34272
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 34272
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 34272
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 34272
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 34272
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 34272
box -86 -90 7254 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 36176 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_8  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 34272
box -86 -90 982 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_30_325
timestamp 1698431365
transform 1 0 37744 0 1 34272
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_30_329
timestamp 1698431365
transform 1 0 38192 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_31_36
timestamp 1698431365
transform 1 0 5376 0 -1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_31_70
timestamp 1698431365
transform 1 0 9184 0 -1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_31_104
timestamp 1698431365
transform 1 0 12992 0 -1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_31_138
timestamp 1698431365
transform 1 0 16800 0 -1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_31_172
timestamp 1698431365
transform 1 0 20608 0 -1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_31_240
timestamp 1698431365
transform 1 0 28224 0 -1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_32  FILLER_0_31_274
timestamp 1698431365
transform 1 0 32032 0 -1 36288
box -86 -90 3670 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_16  FILLER_0_31_308
timestamp 1698431365
transform 1 0 35840 0 -1 36288
box -86 -90 1878 1098
use gf180mcu_fd_sc_mcu9t5v0__fillcap_4  FILLER_0_31_324
timestamp 1698431365
transform 1 0 37632 0 -1 36288
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_2  FILLER_0_31_328
timestamp 1698431365
transform 1 0 38080 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__fill_1  FILLER_0_31_330
timestamp 1698431365
transform 1 0 38304 0 -1 36288
box -86 -90 198 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_0_Left_32 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 4032
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 38640 0 1 4032
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_1_Left_33
timestamp 1698431365
transform 1 0 1344 0 -1 6048
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 38640 0 -1 6048
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_2_Left_34
timestamp 1698431365
transform 1 0 1344 0 1 6048
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 38640 0 1 6048
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_3_Left_35
timestamp 1698431365
transform 1 0 1344 0 -1 8064
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 38640 0 -1 8064
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_4_Left_36
timestamp 1698431365
transform 1 0 1344 0 1 8064
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 38640 0 1 8064
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_5_Left_37
timestamp 1698431365
transform 1 0 1344 0 -1 10080
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 38640 0 -1 10080
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_6_Left_38
timestamp 1698431365
transform 1 0 1344 0 1 10080
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 38640 0 1 10080
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_7_Left_39
timestamp 1698431365
transform 1 0 1344 0 -1 12096
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 38640 0 -1 12096
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_8_Left_40
timestamp 1698431365
transform 1 0 1344 0 1 12096
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 38640 0 1 12096
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_9_Left_41
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 38640 0 -1 14112
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_10_Left_42
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 38640 0 1 14112
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_11_Left_43
timestamp 1698431365
transform 1 0 1344 0 -1 16128
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 38640 0 -1 16128
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_12_Left_44
timestamp 1698431365
transform 1 0 1344 0 1 16128
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 38640 0 1 16128
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_13_Left_45
timestamp 1698431365
transform 1 0 1344 0 -1 18144
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 38640 0 -1 18144
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_14_Left_46
timestamp 1698431365
transform 1 0 1344 0 1 18144
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 38640 0 1 18144
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_15_Left_47
timestamp 1698431365
transform 1 0 1344 0 -1 20160
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 38640 0 -1 20160
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_16_Left_48
timestamp 1698431365
transform 1 0 1344 0 1 20160
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 38640 0 1 20160
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_17_Left_49
timestamp 1698431365
transform 1 0 1344 0 -1 22176
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 38640 0 -1 22176
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_18_Left_50
timestamp 1698431365
transform 1 0 1344 0 1 22176
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 38640 0 1 22176
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_19_Left_51
timestamp 1698431365
transform 1 0 1344 0 -1 24192
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 38640 0 -1 24192
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_20_Left_52
timestamp 1698431365
transform 1 0 1344 0 1 24192
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 38640 0 1 24192
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_21_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 26208
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 38640 0 -1 26208
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_22_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 26208
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 38640 0 1 26208
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_23_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 38640 0 -1 28224
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_24_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 38640 0 1 28224
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_25_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 30240
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 38640 0 -1 30240
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_26_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 30240
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 38640 0 1 30240
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_27_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 32256
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 38640 0 -1 32256
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_28_Left_60
timestamp 1698431365
transform 1 0 1344 0 1 32256
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 38640 0 1 32256
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_29_Left_61
timestamp 1698431365
transform 1 0 1344 0 -1 34272
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 38640 0 -1 34272
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_30_Left_62
timestamp 1698431365
transform 1 0 1344 0 1 34272
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 38640 0 1 34272
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_31_Left_63
timestamp 1698431365
transform 1 0 1344 0 -1 36288
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 38640 0 -1 36288
box -586 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_64 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_65
timestamp 1698431365
transform 1 0 8960 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_66
timestamp 1698431365
transform 1 0 12768 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_67
timestamp 1698431365
transform 1 0 16576 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_68
timestamp 1698431365
transform 1 0 20384 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_69
timestamp 1698431365
transform 1 0 24192 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_70
timestamp 1698431365
transform 1 0 28000 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_71
timestamp 1698431365
transform 1 0 31808 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_0_72
timestamp 1698431365
transform 1 0 35616 0 1 4032
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_73
timestamp 1698431365
transform 1 0 9184 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_74
timestamp 1698431365
transform 1 0 17024 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_75
timestamp 1698431365
transform 1 0 24864 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_1_76
timestamp 1698431365
transform 1 0 32704 0 -1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_77
timestamp 1698431365
transform 1 0 5264 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_78
timestamp 1698431365
transform 1 0 13104 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_79
timestamp 1698431365
transform 1 0 20944 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_80
timestamp 1698431365
transform 1 0 28784 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_2_81
timestamp 1698431365
transform 1 0 36624 0 1 6048
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_82
timestamp 1698431365
transform 1 0 9184 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_83
timestamp 1698431365
transform 1 0 17024 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_84
timestamp 1698431365
transform 1 0 24864 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_3_85
timestamp 1698431365
transform 1 0 32704 0 -1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_86
timestamp 1698431365
transform 1 0 5264 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_87
timestamp 1698431365
transform 1 0 13104 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_88
timestamp 1698431365
transform 1 0 20944 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_89
timestamp 1698431365
transform 1 0 28784 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_4_90
timestamp 1698431365
transform 1 0 36624 0 1 8064
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_91
timestamp 1698431365
transform 1 0 9184 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_92
timestamp 1698431365
transform 1 0 17024 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_93
timestamp 1698431365
transform 1 0 24864 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_5_94
timestamp 1698431365
transform 1 0 32704 0 -1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_95
timestamp 1698431365
transform 1 0 5264 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_96
timestamp 1698431365
transform 1 0 13104 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_97
timestamp 1698431365
transform 1 0 20944 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_98
timestamp 1698431365
transform 1 0 28784 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_6_99
timestamp 1698431365
transform 1 0 36624 0 1 10080
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_100
timestamp 1698431365
transform 1 0 9184 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_101
timestamp 1698431365
transform 1 0 17024 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_102
timestamp 1698431365
transform 1 0 24864 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_7_103
timestamp 1698431365
transform 1 0 32704 0 -1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_104
timestamp 1698431365
transform 1 0 5264 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_105
timestamp 1698431365
transform 1 0 13104 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_106
timestamp 1698431365
transform 1 0 20944 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_107
timestamp 1698431365
transform 1 0 28784 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_8_108
timestamp 1698431365
transform 1 0 36624 0 1 12096
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_109
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_110
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_111
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_9_112
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_113
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_114
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_115
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_116
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_10_117
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_118
timestamp 1698431365
transform 1 0 9184 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_119
timestamp 1698431365
transform 1 0 17024 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_120
timestamp 1698431365
transform 1 0 24864 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_11_121
timestamp 1698431365
transform 1 0 32704 0 -1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_122
timestamp 1698431365
transform 1 0 5264 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_123
timestamp 1698431365
transform 1 0 13104 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_124
timestamp 1698431365
transform 1 0 20944 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_125
timestamp 1698431365
transform 1 0 28784 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_12_126
timestamp 1698431365
transform 1 0 36624 0 1 16128
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_127
timestamp 1698431365
transform 1 0 9184 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_128
timestamp 1698431365
transform 1 0 17024 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_129
timestamp 1698431365
transform 1 0 24864 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_13_130
timestamp 1698431365
transform 1 0 32704 0 -1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_131
timestamp 1698431365
transform 1 0 5264 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_132
timestamp 1698431365
transform 1 0 13104 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_133
timestamp 1698431365
transform 1 0 20944 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_134
timestamp 1698431365
transform 1 0 28784 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_14_135
timestamp 1698431365
transform 1 0 36624 0 1 18144
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_136
timestamp 1698431365
transform 1 0 9184 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_137
timestamp 1698431365
transform 1 0 17024 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_138
timestamp 1698431365
transform 1 0 24864 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_15_139
timestamp 1698431365
transform 1 0 32704 0 -1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_140
timestamp 1698431365
transform 1 0 5264 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_141
timestamp 1698431365
transform 1 0 13104 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_142
timestamp 1698431365
transform 1 0 20944 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_143
timestamp 1698431365
transform 1 0 28784 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_16_144
timestamp 1698431365
transform 1 0 36624 0 1 20160
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_145
timestamp 1698431365
transform 1 0 9184 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_146
timestamp 1698431365
transform 1 0 17024 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_147
timestamp 1698431365
transform 1 0 24864 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_17_148
timestamp 1698431365
transform 1 0 32704 0 -1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_149
timestamp 1698431365
transform 1 0 5264 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_150
timestamp 1698431365
transform 1 0 13104 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_151
timestamp 1698431365
transform 1 0 20944 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_152
timestamp 1698431365
transform 1 0 28784 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_18_153
timestamp 1698431365
transform 1 0 36624 0 1 22176
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_154
timestamp 1698431365
transform 1 0 9184 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_155
timestamp 1698431365
transform 1 0 17024 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_156
timestamp 1698431365
transform 1 0 24864 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_19_157
timestamp 1698431365
transform 1 0 32704 0 -1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_158
timestamp 1698431365
transform 1 0 5264 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_159
timestamp 1698431365
transform 1 0 13104 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_160
timestamp 1698431365
transform 1 0 20944 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_161
timestamp 1698431365
transform 1 0 28784 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_20_162
timestamp 1698431365
transform 1 0 36624 0 1 24192
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_163
timestamp 1698431365
transform 1 0 9184 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_164
timestamp 1698431365
transform 1 0 17024 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_165
timestamp 1698431365
transform 1 0 24864 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_21_166
timestamp 1698431365
transform 1 0 32704 0 -1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_167
timestamp 1698431365
transform 1 0 5264 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_168
timestamp 1698431365
transform 1 0 13104 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_169
timestamp 1698431365
transform 1 0 20944 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_170
timestamp 1698431365
transform 1 0 28784 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_22_171
timestamp 1698431365
transform 1 0 36624 0 1 26208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_172
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_173
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_174
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_23_175
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_176
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_177
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_178
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_179
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_24_180
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_181
timestamp 1698431365
transform 1 0 9184 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_182
timestamp 1698431365
transform 1 0 17024 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_183
timestamp 1698431365
transform 1 0 24864 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_25_184
timestamp 1698431365
transform 1 0 32704 0 -1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_185
timestamp 1698431365
transform 1 0 5264 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_186
timestamp 1698431365
transform 1 0 13104 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_187
timestamp 1698431365
transform 1 0 20944 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_188
timestamp 1698431365
transform 1 0 28784 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_26_189
timestamp 1698431365
transform 1 0 36624 0 1 30240
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_190
timestamp 1698431365
transform 1 0 9184 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_191
timestamp 1698431365
transform 1 0 17024 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_192
timestamp 1698431365
transform 1 0 24864 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_27_193
timestamp 1698431365
transform 1 0 32704 0 -1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_194
timestamp 1698431365
transform 1 0 5264 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_195
timestamp 1698431365
transform 1 0 13104 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_196
timestamp 1698431365
transform 1 0 20944 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_197
timestamp 1698431365
transform 1 0 28784 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_28_198
timestamp 1698431365
transform 1 0 36624 0 1 32256
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_199
timestamp 1698431365
transform 1 0 9184 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_200
timestamp 1698431365
transform 1 0 17024 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_201
timestamp 1698431365
transform 1 0 24864 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_29_202
timestamp 1698431365
transform 1 0 32704 0 -1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_203
timestamp 1698431365
transform 1 0 5264 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_204
timestamp 1698431365
transform 1 0 13104 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_205
timestamp 1698431365
transform 1 0 20944 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_206
timestamp 1698431365
transform 1 0 28784 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_30_207
timestamp 1698431365
transform 1 0 36624 0 1 34272
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_208
timestamp 1698431365
transform 1 0 5152 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_209
timestamp 1698431365
transform 1 0 8960 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_210
timestamp 1698431365
transform 1 0 12768 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_211
timestamp 1698431365
transform 1 0 16576 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_212
timestamp 1698431365
transform 1 0 20384 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_213
timestamp 1698431365
transform 1 0 24192 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_214
timestamp 1698431365
transform 1 0 28000 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_215
timestamp 1698431365
transform 1 0 31808 0 -1 36288
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  TAP_TAPCELL_ROW_31_216
timestamp 1698431365
transform 1 0 35616 0 -1 36288
box -86 -90 310 1098
<< labels >>
flabel metal2 s 14784 39200 14896 40000 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 in[0]
port 1 nsew signal input
flabel metal3 s 39200 14784 40000 14896 0 FreeSans 448 0 0 0 in[10]
port 2 nsew signal input
flabel metal3 s 39200 25536 40000 25648 0 FreeSans 448 0 0 0 in[11]
port 3 nsew signal input
flabel metal3 s 39200 16800 40000 16912 0 FreeSans 448 0 0 0 in[12]
port 4 nsew signal input
flabel metal3 s 39200 17472 40000 17584 0 FreeSans 448 0 0 0 in[13]
port 5 nsew signal input
flabel metal3 s 39200 18816 40000 18928 0 FreeSans 448 0 0 0 in[14]
port 6 nsew signal input
flabel metal3 s 39200 16128 40000 16240 0 FreeSans 448 0 0 0 in[15]
port 7 nsew signal input
flabel metal3 s 39200 19488 40000 19600 0 FreeSans 448 0 0 0 in[16]
port 8 nsew signal input
flabel metal3 s 39200 20160 40000 20272 0 FreeSans 448 0 0 0 in[17]
port 9 nsew signal input
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 in[1]
port 10 nsew signal input
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 in[2]
port 11 nsew signal input
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 in[3]
port 12 nsew signal input
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 in[4]
port 13 nsew signal input
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 in[5]
port 14 nsew signal input
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 in[6]
port 15 nsew signal input
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 in[7]
port 16 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 in[8]
port 17 nsew signal input
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 in[9]
port 18 nsew signal input
flabel metal2 s 15456 39200 15568 40000 0 FreeSans 448 90 0 0 out[0]
port 19 nsew signal tristate
flabel metal3 s 39200 18144 40000 18256 0 FreeSans 448 0 0 0 out[10]
port 20 nsew signal tristate
flabel metal3 s 39200 23520 40000 23632 0 FreeSans 448 0 0 0 out[11]
port 21 nsew signal tristate
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 out[1]
port 22 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 out[2]
port 23 nsew signal tristate
flabel metal3 s 39200 24192 40000 24304 0 FreeSans 448 0 0 0 out[3]
port 24 nsew signal tristate
flabel metal3 s 39200 22176 40000 22288 0 FreeSans 448 0 0 0 out[4]
port 25 nsew signal tristate
flabel metal3 s 39200 22848 40000 22960 0 FreeSans 448 0 0 0 out[5]
port 26 nsew signal tristate
flabel metal3 s 39200 15456 40000 15568 0 FreeSans 448 0 0 0 out[6]
port 27 nsew signal tristate
flabel metal3 s 39200 24864 40000 24976 0 FreeSans 448 0 0 0 out[7]
port 28 nsew signal tristate
flabel metal3 s 39200 21504 40000 21616 0 FreeSans 448 0 0 0 out[8]
port 29 nsew signal tristate
flabel metal3 s 39200 20832 40000 20944 0 FreeSans 448 0 0 0 out[9]
port 30 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 rst_n
port 31 nsew signal input
flabel metal4 s 5846 3972 6166 36348 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 15170 3972 15490 36348 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 24494 3972 24814 36348 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 33818 3972 34138 36348 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 10508 3972 10828 36348 0 FreeSans 1280 90 0 0 vss
port 33 nsew ground bidirectional
flabel metal4 s 19832 3972 20152 36348 0 FreeSans 1280 90 0 0 vss
port 33 nsew ground bidirectional
flabel metal4 s 29156 3972 29476 36348 0 FreeSans 1280 90 0 0 vss
port 33 nsew ground bidirectional
flabel metal4 s 38480 3972 38800 36348 0 FreeSans 1280 90 0 0 vss
port 33 nsew ground bidirectional
rlabel metal1 19992 35280 19992 35280 0 vdd
rlabel via1 20072 36288 20072 36288 0 vss
rlabel metal2 12712 19320 12712 19320 0 _00_
rlabel metal2 13496 20300 13496 20300 0 _01_
rlabel metal2 13832 19208 13832 19208 0 _02_
rlabel metal2 14504 19656 14504 19656 0 _03_
rlabel metal2 16632 19208 16632 19208 0 _04_
rlabel metal2 19152 20552 19152 20552 0 _05_
rlabel metal2 20440 20356 20440 20356 0 _06_
rlabel metal3 22176 20552 22176 20552 0 _07_
rlabel metal2 26152 20356 26152 20356 0 _08_
rlabel metal2 28840 20552 28840 20552 0 _09_
rlabel metal3 28952 20384 28952 20384 0 _10_
rlabel metal2 15064 31864 15064 31864 0 clk
rlabel metal3 2422 16184 2422 16184 0 in[0]
rlabel metal3 23632 20440 23632 20440 0 in[10]
rlabel metal2 22904 19712 22904 19712 0 in[11]
rlabel metal2 25816 19152 25816 19152 0 in[12]
rlabel metal2 23464 18144 23464 18144 0 in[13]
rlabel metal3 28280 18536 28280 18536 0 in[14]
rlabel metal3 28224 19544 28224 19544 0 in[15]
rlabel metal3 30184 18648 30184 18648 0 in[16]
rlabel metal2 30968 19768 30968 19768 0 in[17]
rlabel metal2 14168 19096 14168 19096 0 in[1]
rlabel metal3 2478 24248 2478 24248 0 in[2]
rlabel metal3 2702 18200 2702 18200 0 in[3]
rlabel metal3 2534 16856 2534 16856 0 in[4]
rlabel metal3 2534 20216 2534 20216 0 in[5]
rlabel metal3 2478 17528 2478 17528 0 in[6]
rlabel metal3 2534 22904 2534 22904 0 in[7]
rlabel metal3 2422 23576 2422 23576 0 in[8]
rlabel metal3 4578 22232 4578 22232 0 in[9]
rlabel metal2 15568 32088 15568 32088 0 out[0]
rlabel metal3 38920 18312 38920 18312 0 out[10]
rlabel metal2 31080 21392 31080 21392 0 out[11]
rlabel metal2 19320 21280 19320 21280 0 out[1]
rlabel metal3 9422 20888 9422 20888 0 out[2]
rlabel metal2 22120 21224 22120 21224 0 out[3]
rlabel metal2 34888 21336 34888 21336 0 out[4]
rlabel metal3 24416 20216 24416 20216 0 out[5]
rlabel metal2 24920 17584 24920 17584 0 out[6]
rlabel metal3 27720 20216 27720 20216 0 out[7]
rlabel metal2 27384 20160 27384 20160 0 out[8]
rlabel metal2 29568 20328 29568 20328 0 out[9]
rlabel metal2 15960 18816 15960 18816 0 rst_n
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
