magic
tech gf180mcuD
magscale 1 5
timestamp 1702354951
<< obsm1 >>
rect 672 1538 59304 48246
<< metal2 >>
rect 29568 49600 29624 50000
rect 29904 49600 29960 50000
rect 30240 49600 30296 50000
rect 30576 49600 30632 50000
rect 30912 49600 30968 50000
rect 31248 49600 31304 50000
rect 31584 49600 31640 50000
rect 32256 49600 32312 50000
rect 32592 49600 32648 50000
rect 32928 49600 32984 50000
rect 0 0 56 400
rect 336 0 392 400
rect 672 0 728 400
rect 1008 0 1064 400
rect 1344 0 1400 400
rect 1680 0 1736 400
rect 2016 0 2072 400
rect 2352 0 2408 400
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 31920 0 31976 400
rect 32256 0 32312 400
rect 32928 0 32984 400
<< obsm2 >>
rect 238 49570 29538 49600
rect 29654 49570 29874 49600
rect 29990 49570 30210 49600
rect 30326 49570 30546 49600
rect 30662 49570 30882 49600
rect 30998 49570 31218 49600
rect 31334 49570 31554 49600
rect 31670 49570 32226 49600
rect 32342 49570 32562 49600
rect 32678 49570 32898 49600
rect 33014 49570 59178 49600
rect 238 430 59178 49570
rect 238 400 306 430
rect 422 400 642 430
rect 758 400 978 430
rect 1094 400 1314 430
rect 1430 400 1650 430
rect 1766 400 1986 430
rect 2102 400 2322 430
rect 2438 400 2658 430
rect 2774 400 2994 430
rect 3110 400 3330 430
rect 3446 400 3666 430
rect 3782 400 31890 430
rect 32006 400 32226 430
rect 32342 400 32898 430
rect 33014 400 59178 430
<< metal3 >>
rect 0 42672 400 42728
rect 59600 25200 60000 25256
rect 59600 24864 60000 24920
rect 0 24528 400 24584
rect 59600 24528 60000 24584
rect 59600 24192 60000 24248
rect 0 23856 400 23912
rect 0 23520 400 23576
<< obsm3 >>
rect 233 42758 59600 48706
rect 430 42642 59600 42758
rect 233 25286 59600 42642
rect 233 25170 59570 25286
rect 233 24950 59600 25170
rect 233 24834 59570 24950
rect 233 24614 59600 24834
rect 430 24498 59570 24614
rect 233 24278 59600 24498
rect 233 24162 59570 24278
rect 233 23942 59600 24162
rect 430 23826 59600 23942
rect 233 23606 59600 23826
rect 430 23490 59600 23606
rect 233 1302 59600 23490
<< metal4 >>
rect 2224 1538 2384 48246
rect 9904 1538 10064 48246
rect 17584 1538 17744 48246
rect 25264 1538 25424 48246
rect 32944 1538 33104 48246
rect 40624 1538 40784 48246
rect 48304 1538 48464 48246
rect 55984 1538 56144 48246
<< obsm4 >>
rect 1078 1508 2194 38127
rect 2414 1508 9874 38127
rect 10094 1508 17554 38127
rect 17774 1508 25234 38127
rect 25454 1508 32914 38127
rect 33134 1508 40594 38127
rect 40814 1508 48274 38127
rect 48494 1508 55954 38127
rect 56174 1508 58170 38127
rect 1078 1353 58170 1508
<< labels >>
rlabel metal3 s 0 42672 400 42728 6 clk
port 1 nsew signal input
rlabel metal2 s 29904 49600 29960 50000 6 in[0]
port 2 nsew signal input
rlabel metal2 s 0 0 56 400 6 in[10]
port 3 nsew signal input
rlabel metal2 s 336 0 392 400 6 in[11]
port 4 nsew signal input
rlabel metal2 s 672 0 728 400 6 in[12]
port 5 nsew signal input
rlabel metal2 s 1008 0 1064 400 6 in[13]
port 6 nsew signal input
rlabel metal2 s 1344 0 1400 400 6 in[14]
port 7 nsew signal input
rlabel metal2 s 1680 0 1736 400 6 in[15]
port 8 nsew signal input
rlabel metal2 s 2016 0 2072 400 6 in[16]
port 9 nsew signal input
rlabel metal2 s 2352 0 2408 400 6 in[17]
port 10 nsew signal input
rlabel metal2 s 2688 0 2744 400 6 in[18]
port 11 nsew signal input
rlabel metal2 s 31248 49600 31304 50000 6 in[1]
port 12 nsew signal input
rlabel metal2 s 29568 49600 29624 50000 6 in[2]
port 13 nsew signal input
rlabel metal3 s 0 23520 400 23576 6 in[3]
port 14 nsew signal input
rlabel metal3 s 0 23856 400 23912 6 in[4]
port 15 nsew signal input
rlabel metal3 s 0 24528 400 24584 6 in[5]
port 16 nsew signal input
rlabel metal2 s 32592 49600 32648 50000 6 in[6]
port 17 nsew signal input
rlabel metal2 s 3024 0 3080 400 6 in[7]
port 18 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 in[8]
port 19 nsew signal input
rlabel metal2 s 3696 0 3752 400 6 in[9]
port 20 nsew signal input
rlabel metal3 s 59600 24864 60000 24920 6 out[0]
port 21 nsew signal output
rlabel metal2 s 30912 49600 30968 50000 6 out[10]
port 22 nsew signal output
rlabel metal3 s 59600 25200 60000 25256 6 out[11]
port 23 nsew signal output
rlabel metal2 s 32928 0 32984 400 6 out[1]
port 24 nsew signal output
rlabel metal2 s 31920 0 31976 400 6 out[2]
port 25 nsew signal output
rlabel metal2 s 32256 0 32312 400 6 out[3]
port 26 nsew signal output
rlabel metal2 s 31584 49600 31640 50000 6 out[4]
port 27 nsew signal output
rlabel metal3 s 59600 24528 60000 24584 6 out[5]
port 28 nsew signal output
rlabel metal3 s 59600 24192 60000 24248 6 out[6]
port 29 nsew signal output
rlabel metal2 s 32928 49600 32984 50000 6 out[7]
port 30 nsew signal output
rlabel metal2 s 30576 49600 30632 50000 6 out[8]
port 31 nsew signal output
rlabel metal2 s 30240 49600 30296 50000 6 out[9]
port 32 nsew signal output
rlabel metal2 s 32256 49600 32312 50000 6 rst_n
port 33 nsew signal input
rlabel metal4 s 2224 1538 2384 48246 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 48246 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 48246 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 48246 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 48246 6 vss
port 35 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 48246 6 vss
port 35 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 48246 6 vss
port 35 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 48246 6 vss
port 35 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6378204
string GDS_FILE /home/htamas/progs/gfmpw1-multi/openlane/totp/runs/23_12_12_05_13/results/signoff/totp.magic.gds
string GDS_START 395712
<< end >>

