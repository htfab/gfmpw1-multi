magic
tech gf180mcuD
magscale 1 5
timestamp 1702441932
<< obsm1 >>
rect 672 1538 23296 22374
<< metal2 >>
rect 0 0 56 400
rect 336 0 392 400
rect 672 0 728 400
rect 1008 0 1064 400
rect 1344 0 1400 400
rect 1680 0 1736 400
rect 2016 0 2072 400
rect 2352 0 2408 400
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
<< obsm2 >>
rect 854 1549 23114 22363
<< metal3 >>
rect 0 21504 400 21560
rect 0 21168 400 21224
rect 23600 21168 24000 21224
rect 0 17136 400 17192
rect 0 13776 400 13832
rect 0 13440 400 13496
rect 0 13104 400 13160
rect 0 12768 400 12824
rect 0 12432 400 12488
rect 0 12096 400 12152
rect 0 11760 400 11816
rect 0 11424 400 11480
rect 0 10752 400 10808
rect 0 10416 400 10472
rect 0 10080 400 10136
rect 0 9744 400 9800
rect 0 9408 400 9464
rect 0 9072 400 9128
rect 0 8400 400 8456
rect 0 2352 400 2408
<< obsm3 >>
rect 350 21590 23600 22358
rect 430 21474 23600 21590
rect 350 21254 23600 21474
rect 430 21138 23570 21254
rect 350 17222 23600 21138
rect 430 17106 23600 17222
rect 350 13862 23600 17106
rect 430 13746 23600 13862
rect 350 13526 23600 13746
rect 430 13410 23600 13526
rect 350 13190 23600 13410
rect 430 13074 23600 13190
rect 350 12854 23600 13074
rect 430 12738 23600 12854
rect 350 12518 23600 12738
rect 430 12402 23600 12518
rect 350 12182 23600 12402
rect 430 12066 23600 12182
rect 350 11846 23600 12066
rect 430 11730 23600 11846
rect 350 11510 23600 11730
rect 430 11394 23600 11510
rect 350 10838 23600 11394
rect 430 10722 23600 10838
rect 350 10502 23600 10722
rect 430 10386 23600 10502
rect 350 10166 23600 10386
rect 430 10050 23600 10166
rect 350 9830 23600 10050
rect 430 9714 23600 9830
rect 350 9494 23600 9714
rect 430 9378 23600 9494
rect 350 9158 23600 9378
rect 430 9042 23600 9158
rect 350 8486 23600 9042
rect 430 8370 23600 8486
rect 350 2438 23600 8370
rect 430 2322 23600 2438
rect 350 1554 23600 2322
<< metal4 >>
rect 2224 1538 2384 22374
rect 9904 1538 10064 22374
rect 17584 1538 17744 22374
<< obsm4 >>
rect 7854 5833 9874 18527
rect 10094 5833 17554 18527
rect 17774 5833 17850 18527
<< labels >>
rlabel metal2 s 0 0 56 400 6 clk
port 1 nsew signal input
rlabel metal3 s 0 17136 400 17192 6 in[0]
port 2 nsew signal input
rlabel metal2 s 336 0 392 400 6 in[10]
port 3 nsew signal input
rlabel metal2 s 672 0 728 400 6 in[11]
port 4 nsew signal input
rlabel metal2 s 1008 0 1064 400 6 in[12]
port 5 nsew signal input
rlabel metal2 s 1344 0 1400 400 6 in[13]
port 6 nsew signal input
rlabel metal2 s 1680 0 1736 400 6 in[14]
port 7 nsew signal input
rlabel metal2 s 2016 0 2072 400 6 in[15]
port 8 nsew signal input
rlabel metal2 s 2352 0 2408 400 6 in[16]
port 9 nsew signal input
rlabel metal2 s 2688 0 2744 400 6 in[17]
port 10 nsew signal input
rlabel metal3 s 0 9408 400 9464 6 in[1]
port 11 nsew signal input
rlabel metal3 s 0 9072 400 9128 6 in[2]
port 12 nsew signal input
rlabel metal3 s 0 8400 400 8456 6 in[3]
port 13 nsew signal input
rlabel metal3 s 0 10752 400 10808 6 in[4]
port 14 nsew signal input
rlabel metal3 s 0 10416 400 10472 6 in[5]
port 15 nsew signal input
rlabel metal3 s 0 10080 400 10136 6 in[6]
port 16 nsew signal input
rlabel metal3 s 0 9744 400 9800 6 in[7]
port 17 nsew signal input
rlabel metal2 s 3024 0 3080 400 6 in[8]
port 18 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 in[9]
port 19 nsew signal input
rlabel metal3 s 0 13104 400 13160 6 out[0]
port 20 nsew signal output
rlabel metal3 s 23600 21168 24000 21224 6 out[10]
port 21 nsew signal output
rlabel metal3 s 0 21504 400 21560 6 out[11]
port 22 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 out[1]
port 23 nsew signal output
rlabel metal3 s 0 12432 400 12488 6 out[2]
port 24 nsew signal output
rlabel metal3 s 0 12096 400 12152 6 out[3]
port 25 nsew signal output
rlabel metal3 s 0 11760 400 11816 6 out[4]
port 26 nsew signal output
rlabel metal3 s 0 11424 400 11480 6 out[5]
port 27 nsew signal output
rlabel metal3 s 0 13776 400 13832 6 out[6]
port 28 nsew signal output
rlabel metal3 s 0 13440 400 13496 6 out[7]
port 29 nsew signal output
rlabel metal3 s 0 21168 400 21224 6 out[8]
port 30 nsew signal output
rlabel metal3 s 0 2352 400 2408 6 out[9]
port 31 nsew signal output
rlabel metal2 s 3696 0 3752 400 6 rst_n
port 32 nsew signal input
rlabel metal4 s 2224 1538 2384 22374 6 vdd
port 33 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 22374 6 vdd
port 33 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 22374 6 vss
port 34 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 24000 24000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2702372
string GDS_FILE /home/htamas/progs/gfmpw1-multi.v2/openlane/cells7/runs/23_12_13_05_28/results/signoff/cells7.magic.gds
string GDS_START 1428956
<< end >>

