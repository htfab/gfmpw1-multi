magic
tech gf180mcuD
magscale 1 5
timestamp 1702353931
<< obsm1 >>
rect 672 1538 7360 6302
<< metal2 >>
rect 4368 7600 4424 8000
rect 4704 7600 4760 8000
rect 5712 7600 5768 8000
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 4032 0 4088 400
rect 4368 0 4424 400
rect 4704 0 4760 400
<< obsm2 >>
rect 854 7570 4338 7600
rect 4454 7570 4674 7600
rect 4790 7570 5682 7600
rect 5798 7570 7346 7600
rect 854 430 7346 7570
rect 854 400 2994 430
rect 3110 400 3330 430
rect 3446 400 3666 430
rect 3782 400 4002 430
rect 4118 400 4338 430
rect 4454 400 4674 430
rect 4790 400 7346 430
<< metal3 >>
rect 7600 7056 8000 7112
rect 7600 6720 8000 6776
rect 7600 6384 8000 6440
rect 7600 6048 8000 6104
rect 7600 5712 8000 5768
rect 7600 5376 8000 5432
rect 7600 5040 8000 5096
rect 0 4704 400 4760
rect 7600 4704 8000 4760
rect 0 4368 400 4424
rect 7600 4368 8000 4424
rect 0 4032 400 4088
rect 7600 4032 8000 4088
rect 0 3696 400 3752
rect 7600 3696 8000 3752
rect 0 3360 400 3416
rect 7600 3360 8000 3416
rect 0 3024 400 3080
rect 7600 3024 8000 3080
rect 0 2688 400 2744
rect 7600 2688 8000 2744
rect 0 2352 400 2408
rect 0 2016 400 2072
rect 0 1680 400 1736
<< obsm3 >>
rect 400 7026 7570 7098
rect 400 6806 7602 7026
rect 400 6690 7570 6806
rect 400 6470 7602 6690
rect 400 6354 7570 6470
rect 400 6134 7602 6354
rect 400 6018 7570 6134
rect 400 5798 7602 6018
rect 400 5682 7570 5798
rect 400 5462 7602 5682
rect 400 5346 7570 5462
rect 400 5126 7602 5346
rect 400 5010 7570 5126
rect 400 4790 7602 5010
rect 430 4674 7570 4790
rect 400 4454 7602 4674
rect 430 4338 7570 4454
rect 400 4118 7602 4338
rect 430 4002 7570 4118
rect 400 3782 7602 4002
rect 430 3666 7570 3782
rect 400 3446 7602 3666
rect 430 3330 7570 3446
rect 400 3110 7602 3330
rect 430 2994 7570 3110
rect 400 2774 7602 2994
rect 430 2658 7570 2774
rect 400 2438 7602 2658
rect 430 2322 7602 2438
rect 400 2102 7602 2322
rect 430 1986 7602 2102
rect 400 1766 7602 1986
rect 430 1650 7602 1766
rect 400 1554 7602 1650
<< metal4 >>
rect 1418 1538 1578 6302
rect 2244 1538 2404 6302
rect 3070 1538 3230 6302
rect 3896 1538 4056 6302
rect 4722 1538 4882 6302
rect 5548 1538 5708 6302
rect 6374 1538 6534 6302
rect 7200 1538 7360 6302
<< labels >>
rlabel metal2 s 3024 0 3080 400 6 clk
port 1 nsew signal input
rlabel metal3 s 0 3360 400 3416 6 in[0]
port 2 nsew signal input
rlabel metal2 s 3696 0 3752 400 6 in[10]
port 3 nsew signal input
rlabel metal3 s 7600 2688 8000 2744 6 in[11]
port 4 nsew signal input
rlabel metal3 s 7600 3024 8000 3080 6 in[12]
port 5 nsew signal input
rlabel metal2 s 4704 7600 4760 8000 6 in[13]
port 6 nsew signal input
rlabel metal2 s 4368 7600 4424 8000 6 in[14]
port 7 nsew signal input
rlabel metal3 s 7600 7056 8000 7112 6 in[15]
port 8 nsew signal input
rlabel metal3 s 7600 5376 8000 5432 6 in[16]
port 9 nsew signal input
rlabel metal3 s 7600 5712 8000 5768 6 in[17]
port 10 nsew signal input
rlabel metal2 s 5712 7600 5768 8000 6 in[18]
port 11 nsew signal input
rlabel metal3 s 0 1680 400 1736 6 in[1]
port 12 nsew signal input
rlabel metal3 s 0 4368 400 4424 6 in[2]
port 13 nsew signal input
rlabel metal3 s 0 2352 400 2408 6 in[3]
port 14 nsew signal input
rlabel metal3 s 0 3024 400 3080 6 in[4]
port 15 nsew signal input
rlabel metal3 s 0 4704 400 4760 6 in[5]
port 16 nsew signal input
rlabel metal3 s 0 4032 400 4088 6 in[6]
port 17 nsew signal input
rlabel metal3 s 0 2016 400 2072 6 in[7]
port 18 nsew signal input
rlabel metal3 s 0 2688 400 2744 6 in[8]
port 19 nsew signal input
rlabel metal2 s 4032 0 4088 400 6 in[9]
port 20 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 out[0]
port 21 nsew signal output
rlabel metal3 s 7600 6720 8000 6776 6 out[10]
port 22 nsew signal output
rlabel metal3 s 7600 6384 8000 6440 6 out[11]
port 23 nsew signal output
rlabel metal2 s 4704 0 4760 400 6 out[1]
port 24 nsew signal output
rlabel metal2 s 4368 0 4424 400 6 out[2]
port 25 nsew signal output
rlabel metal3 s 7600 3360 8000 3416 6 out[3]
port 26 nsew signal output
rlabel metal3 s 7600 3696 8000 3752 6 out[4]
port 27 nsew signal output
rlabel metal3 s 7600 4032 8000 4088 6 out[5]
port 28 nsew signal output
rlabel metal3 s 7600 4368 8000 4424 6 out[6]
port 29 nsew signal output
rlabel metal3 s 7600 5040 8000 5096 6 out[7]
port 30 nsew signal output
rlabel metal3 s 7600 4704 8000 4760 6 out[8]
port 31 nsew signal output
rlabel metal3 s 7600 6048 8000 6104 6 out[9]
port 32 nsew signal output
rlabel metal3 s 0 3696 400 3752 6 rst_n
port 33 nsew signal input
rlabel metal4 s 1418 1538 1578 6302 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 3070 1538 3230 6302 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 4722 1538 4882 6302 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 6374 1538 6534 6302 6 vdd
port 34 nsew power bidirectional
rlabel metal4 s 2244 1538 2404 6302 6 vss
port 35 nsew ground bidirectional
rlabel metal4 s 3896 1538 4056 6302 6 vss
port 35 nsew ground bidirectional
rlabel metal4 s 5548 1538 5708 6302 6 vss
port 35 nsew ground bidirectional
rlabel metal4 s 7200 1538 7360 6302 6 vss
port 35 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 8000 8000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 176462
string GDS_FILE /home/htamas/progs/gfmpw1-multi/openlane/loopback/runs/23_12_12_05_02/results/signoff/loopback.magic.gds
string GDS_START 54574
<< end >>

