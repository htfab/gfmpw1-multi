module user_project_wrapper (user_clock2,
    vdd,
    vss,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input vdd;
 input vss;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire clk;
 wire \in[0] ;
 wire \in[10] ;
 wire \in[11] ;
 wire \in[12] ;
 wire \in[13] ;
 wire \in[14] ;
 wire \in[15] ;
 wire \in[16] ;
 wire \in[17] ;
 wire \in[1] ;
 wire \in[2] ;
 wire \in[3] ;
 wire \in[4] ;
 wire \in[5] ;
 wire \in[6] ;
 wire \in[7] ;
 wire \in[8] ;
 wire \in[9] ;
 wire \out[0] ;
 wire \out[10] ;
 wire \out[11] ;
 wire \out[1] ;
 wire \out[2] ;
 wire \out[3] ;
 wire \out[4] ;
 wire \out[5] ;
 wire \out[6] ;
 wire \out[7] ;
 wire \out[8] ;
 wire \out[9] ;
 wire \proj_clk[0] ;
 wire \proj_clk[1] ;
 wire \proj_clk[2] ;
 wire \proj_clk[3] ;
 wire \proj_clk[4] ;
 wire \proj_clk[5] ;
 wire \proj_clk[6] ;
 wire \proj_clk[7] ;
 wire \proj_in[0] ;
 wire \proj_in[100] ;
 wire \proj_in[101] ;
 wire \proj_in[102] ;
 wire \proj_in[103] ;
 wire \proj_in[104] ;
 wire \proj_in[105] ;
 wire \proj_in[106] ;
 wire \proj_in[107] ;
 wire \proj_in[108] ;
 wire \proj_in[109] ;
 wire \proj_in[10] ;
 wire \proj_in[110] ;
 wire \proj_in[111] ;
 wire \proj_in[112] ;
 wire \proj_in[113] ;
 wire \proj_in[114] ;
 wire \proj_in[115] ;
 wire \proj_in[116] ;
 wire \proj_in[117] ;
 wire \proj_in[118] ;
 wire \proj_in[119] ;
 wire \proj_in[11] ;
 wire \proj_in[120] ;
 wire \proj_in[121] ;
 wire \proj_in[122] ;
 wire \proj_in[123] ;
 wire \proj_in[124] ;
 wire \proj_in[125] ;
 wire \proj_in[126] ;
 wire \proj_in[127] ;
 wire \proj_in[128] ;
 wire \proj_in[129] ;
 wire \proj_in[12] ;
 wire \proj_in[130] ;
 wire \proj_in[131] ;
 wire \proj_in[132] ;
 wire \proj_in[133] ;
 wire \proj_in[134] ;
 wire \proj_in[135] ;
 wire \proj_in[136] ;
 wire \proj_in[137] ;
 wire \proj_in[138] ;
 wire \proj_in[139] ;
 wire \proj_in[13] ;
 wire \proj_in[140] ;
 wire \proj_in[141] ;
 wire \proj_in[142] ;
 wire \proj_in[143] ;
 wire \proj_in[14] ;
 wire \proj_in[15] ;
 wire \proj_in[16] ;
 wire \proj_in[17] ;
 wire \proj_in[18] ;
 wire \proj_in[19] ;
 wire \proj_in[1] ;
 wire \proj_in[20] ;
 wire \proj_in[21] ;
 wire \proj_in[22] ;
 wire \proj_in[23] ;
 wire \proj_in[24] ;
 wire \proj_in[25] ;
 wire \proj_in[26] ;
 wire \proj_in[27] ;
 wire \proj_in[28] ;
 wire \proj_in[29] ;
 wire \proj_in[2] ;
 wire \proj_in[30] ;
 wire \proj_in[31] ;
 wire \proj_in[32] ;
 wire \proj_in[33] ;
 wire \proj_in[34] ;
 wire \proj_in[35] ;
 wire \proj_in[36] ;
 wire \proj_in[37] ;
 wire \proj_in[38] ;
 wire \proj_in[39] ;
 wire \proj_in[3] ;
 wire \proj_in[40] ;
 wire \proj_in[41] ;
 wire \proj_in[42] ;
 wire \proj_in[43] ;
 wire \proj_in[44] ;
 wire \proj_in[45] ;
 wire \proj_in[46] ;
 wire \proj_in[47] ;
 wire \proj_in[48] ;
 wire \proj_in[49] ;
 wire \proj_in[4] ;
 wire \proj_in[50] ;
 wire \proj_in[51] ;
 wire \proj_in[52] ;
 wire \proj_in[53] ;
 wire \proj_in[54] ;
 wire \proj_in[55] ;
 wire \proj_in[56] ;
 wire \proj_in[57] ;
 wire \proj_in[58] ;
 wire \proj_in[59] ;
 wire \proj_in[5] ;
 wire \proj_in[60] ;
 wire \proj_in[61] ;
 wire \proj_in[62] ;
 wire \proj_in[63] ;
 wire \proj_in[64] ;
 wire \proj_in[65] ;
 wire \proj_in[66] ;
 wire \proj_in[67] ;
 wire \proj_in[68] ;
 wire \proj_in[69] ;
 wire \proj_in[6] ;
 wire \proj_in[70] ;
 wire \proj_in[71] ;
 wire \proj_in[72] ;
 wire \proj_in[73] ;
 wire \proj_in[74] ;
 wire \proj_in[75] ;
 wire \proj_in[76] ;
 wire \proj_in[77] ;
 wire \proj_in[78] ;
 wire \proj_in[79] ;
 wire \proj_in[7] ;
 wire \proj_in[80] ;
 wire \proj_in[81] ;
 wire \proj_in[82] ;
 wire \proj_in[83] ;
 wire \proj_in[84] ;
 wire \proj_in[85] ;
 wire \proj_in[86] ;
 wire \proj_in[87] ;
 wire \proj_in[88] ;
 wire \proj_in[89] ;
 wire \proj_in[8] ;
 wire \proj_in[90] ;
 wire \proj_in[91] ;
 wire \proj_in[92] ;
 wire \proj_in[93] ;
 wire \proj_in[94] ;
 wire \proj_in[95] ;
 wire \proj_in[96] ;
 wire \proj_in[97] ;
 wire \proj_in[98] ;
 wire \proj_in[99] ;
 wire \proj_in[9] ;
 wire \proj_out[0] ;
 wire \proj_out[10] ;
 wire \proj_out[11] ;
 wire \proj_out[12] ;
 wire \proj_out[13] ;
 wire \proj_out[14] ;
 wire \proj_out[15] ;
 wire \proj_out[16] ;
 wire \proj_out[17] ;
 wire \proj_out[18] ;
 wire \proj_out[19] ;
 wire \proj_out[1] ;
 wire \proj_out[20] ;
 wire \proj_out[21] ;
 wire \proj_out[22] ;
 wire \proj_out[23] ;
 wire \proj_out[24] ;
 wire \proj_out[25] ;
 wire \proj_out[26] ;
 wire \proj_out[27] ;
 wire \proj_out[28] ;
 wire \proj_out[29] ;
 wire \proj_out[2] ;
 wire \proj_out[30] ;
 wire \proj_out[31] ;
 wire \proj_out[32] ;
 wire \proj_out[33] ;
 wire \proj_out[34] ;
 wire \proj_out[35] ;
 wire \proj_out[36] ;
 wire \proj_out[37] ;
 wire \proj_out[38] ;
 wire \proj_out[39] ;
 wire \proj_out[3] ;
 wire \proj_out[40] ;
 wire \proj_out[41] ;
 wire \proj_out[42] ;
 wire \proj_out[43] ;
 wire \proj_out[44] ;
 wire \proj_out[45] ;
 wire \proj_out[46] ;
 wire \proj_out[47] ;
 wire \proj_out[48] ;
 wire \proj_out[49] ;
 wire \proj_out[4] ;
 wire \proj_out[50] ;
 wire \proj_out[51] ;
 wire \proj_out[52] ;
 wire \proj_out[53] ;
 wire \proj_out[54] ;
 wire \proj_out[55] ;
 wire \proj_out[56] ;
 wire \proj_out[57] ;
 wire \proj_out[58] ;
 wire \proj_out[59] ;
 wire \proj_out[5] ;
 wire \proj_out[60] ;
 wire \proj_out[61] ;
 wire \proj_out[62] ;
 wire \proj_out[63] ;
 wire \proj_out[64] ;
 wire \proj_out[65] ;
 wire \proj_out[66] ;
 wire \proj_out[67] ;
 wire \proj_out[68] ;
 wire \proj_out[69] ;
 wire \proj_out[6] ;
 wire \proj_out[70] ;
 wire \proj_out[71] ;
 wire \proj_out[72] ;
 wire \proj_out[73] ;
 wire \proj_out[74] ;
 wire \proj_out[75] ;
 wire \proj_out[76] ;
 wire \proj_out[77] ;
 wire \proj_out[78] ;
 wire \proj_out[79] ;
 wire \proj_out[7] ;
 wire \proj_out[80] ;
 wire \proj_out[81] ;
 wire \proj_out[82] ;
 wire \proj_out[83] ;
 wire \proj_out[84] ;
 wire \proj_out[85] ;
 wire \proj_out[86] ;
 wire \proj_out[87] ;
 wire \proj_out[88] ;
 wire \proj_out[89] ;
 wire \proj_out[8] ;
 wire \proj_out[90] ;
 wire \proj_out[91] ;
 wire \proj_out[92] ;
 wire \proj_out[93] ;
 wire \proj_out[94] ;
 wire \proj_out[95] ;
 wire \proj_out[9] ;
 wire \proj_rst_n[0] ;
 wire \proj_rst_n[1] ;
 wire \proj_rst_n[2] ;
 wire \proj_rst_n[3] ;
 wire \proj_rst_n[4] ;
 wire \proj_rst_n[5] ;
 wire \proj_rst_n[6] ;
 wire \proj_rst_n[7] ;
 wire rst_n;
 wire \sel[0] ;
 wire \sel[1] ;
 wire \sel[2] ;

 caravel_if ci (.clk(clk),
    .rst_n(rst_n),
    .user_clock2(user_clock2),
    .vdd(vdd),
    .vss(vss),
    .wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),
    .wbs_ack_o(wbs_ack_o),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(wbs_stb_i),
    .wbs_we_i(wbs_we_i),
    .in({\in[17] ,
    \in[16] ,
    \in[15] ,
    \in[14] ,
    \in[13] ,
    \in[12] ,
    \in[11] ,
    \in[10] ,
    \in[9] ,
    \in[8] ,
    \in[7] ,
    \in[6] ,
    \in[5] ,
    \in[4] ,
    \in[3] ,
    \in[2] ,
    \in[1] ,
    \in[0] }),
    .io_in({io_in[37],
    io_in[36],
    io_in[35],
    io_in[34],
    io_in[33],
    io_in[32],
    io_in[31],
    io_in[30],
    io_in[29],
    io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24],
    io_in[23],
    io_in[22],
    io_in[21],
    io_in[20],
    io_in[19],
    io_in[18],
    io_in[17],
    io_in[16],
    io_in[15],
    io_in[14],
    io_in[13],
    io_in[12],
    io_in[11],
    io_in[10],
    io_in[9],
    io_in[8],
    io_in[7],
    io_in[6],
    io_in[5],
    io_in[4],
    io_in[3],
    io_in[2],
    io_in[1],
    io_in[0]}),
    .io_oeb({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21],
    io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13],
    io_oeb[12],
    io_oeb[11],
    io_oeb[10],
    io_oeb[9],
    io_oeb[8],
    io_oeb[7],
    io_oeb[6],
    io_oeb[5],
    io_oeb[4],
    io_oeb[3],
    io_oeb[2],
    io_oeb[1],
    io_oeb[0]}),
    .io_out({io_out[37],
    io_out[36],
    io_out[35],
    io_out[34],
    io_out[33],
    io_out[32],
    io_out[31],
    io_out[30],
    io_out[29],
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24],
    io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16],
    io_out[15],
    io_out[14],
    io_out[13],
    io_out[12],
    io_out[11],
    io_out[10],
    io_out[9],
    io_out[8],
    io_out[7],
    io_out[6],
    io_out[5],
    io_out[4],
    io_out[3],
    io_out[2],
    io_out[1],
    io_out[0]}),
    .la_data_in({la_data_in[63],
    la_data_in[62],
    la_data_in[61],
    la_data_in[60],
    la_data_in[59],
    la_data_in[58],
    la_data_in[57],
    la_data_in[56],
    la_data_in[55],
    la_data_in[54],
    la_data_in[53],
    la_data_in[52],
    la_data_in[51],
    la_data_in[50],
    la_data_in[49],
    la_data_in[48],
    la_data_in[47],
    la_data_in[46],
    la_data_in[45],
    la_data_in[44],
    la_data_in[43],
    la_data_in[42],
    la_data_in[41],
    la_data_in[40],
    la_data_in[39],
    la_data_in[38],
    la_data_in[37],
    la_data_in[36],
    la_data_in[35],
    la_data_in[34],
    la_data_in[33],
    la_data_in[32],
    la_data_in[31],
    la_data_in[30],
    la_data_in[29],
    la_data_in[28],
    la_data_in[27],
    la_data_in[26],
    la_data_in[25],
    la_data_in[24],
    la_data_in[23],
    la_data_in[22],
    la_data_in[21],
    la_data_in[20],
    la_data_in[19],
    la_data_in[18],
    la_data_in[17],
    la_data_in[16],
    la_data_in[15],
    la_data_in[14],
    la_data_in[13],
    la_data_in[12],
    la_data_in[11],
    la_data_in[10],
    la_data_in[9],
    la_data_in[8],
    la_data_in[7],
    la_data_in[6],
    la_data_in[5],
    la_data_in[4],
    la_data_in[3],
    la_data_in[2],
    la_data_in[1],
    la_data_in[0]}),
    .la_data_out({la_data_out[63],
    la_data_out[62],
    la_data_out[61],
    la_data_out[60],
    la_data_out[59],
    la_data_out[58],
    la_data_out[57],
    la_data_out[56],
    la_data_out[55],
    la_data_out[54],
    la_data_out[53],
    la_data_out[52],
    la_data_out[51],
    la_data_out[50],
    la_data_out[49],
    la_data_out[48],
    la_data_out[47],
    la_data_out[46],
    la_data_out[45],
    la_data_out[44],
    la_data_out[43],
    la_data_out[42],
    la_data_out[41],
    la_data_out[40],
    la_data_out[39],
    la_data_out[38],
    la_data_out[37],
    la_data_out[36],
    la_data_out[35],
    la_data_out[34],
    la_data_out[33],
    la_data_out[32],
    la_data_out[31],
    la_data_out[30],
    la_data_out[29],
    la_data_out[28],
    la_data_out[27],
    la_data_out[26],
    la_data_out[25],
    la_data_out[24],
    la_data_out[23],
    la_data_out[22],
    la_data_out[21],
    la_data_out[20],
    la_data_out[19],
    la_data_out[18],
    la_data_out[17],
    la_data_out[16],
    la_data_out[15],
    la_data_out[14],
    la_data_out[13],
    la_data_out[12],
    la_data_out[11],
    la_data_out[10],
    la_data_out[9],
    la_data_out[8],
    la_data_out[7],
    la_data_out[6],
    la_data_out[5],
    la_data_out[4],
    la_data_out[3],
    la_data_out[2],
    la_data_out[1],
    la_data_out[0]}),
    .la_oenb({la_oenb[63],
    la_oenb[62],
    la_oenb[61],
    la_oenb[60],
    la_oenb[59],
    la_oenb[58],
    la_oenb[57],
    la_oenb[56],
    la_oenb[55],
    la_oenb[54],
    la_oenb[53],
    la_oenb[52],
    la_oenb[51],
    la_oenb[50],
    la_oenb[49],
    la_oenb[48],
    la_oenb[47],
    la_oenb[46],
    la_oenb[45],
    la_oenb[44],
    la_oenb[43],
    la_oenb[42],
    la_oenb[41],
    la_oenb[40],
    la_oenb[39],
    la_oenb[38],
    la_oenb[37],
    la_oenb[36],
    la_oenb[35],
    la_oenb[34],
    la_oenb[33],
    la_oenb[32],
    la_oenb[31],
    la_oenb[30],
    la_oenb[29],
    la_oenb[28],
    la_oenb[27],
    la_oenb[26],
    la_oenb[25],
    la_oenb[24],
    la_oenb[23],
    la_oenb[22],
    la_oenb[21],
    la_oenb[20],
    la_oenb[19],
    la_oenb[18],
    la_oenb[17],
    la_oenb[16],
    la_oenb[15],
    la_oenb[14],
    la_oenb[13],
    la_oenb[12],
    la_oenb[11],
    la_oenb[10],
    la_oenb[9],
    la_oenb[8],
    la_oenb[7],
    la_oenb[6],
    la_oenb[5],
    la_oenb[4],
    la_oenb[3],
    la_oenb[2],
    la_oenb[1],
    la_oenb[0]}),
    .out({\out[11] ,
    \out[10] ,
    \out[9] ,
    \out[8] ,
    \out[7] ,
    \out[6] ,
    \out[5] ,
    \out[4] ,
    \out[3] ,
    \out[2] ,
    \out[1] ,
    \out[0] }),
    .sel({\sel[2] ,
    \sel[1] ,
    \sel[0] }),
    .user_irq({user_irq[2],
    user_irq[1],
    user_irq[0]}),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({wbs_dat_o[31],
    wbs_dat_o[30],
    wbs_dat_o[29],
    wbs_dat_o[28],
    wbs_dat_o[27],
    wbs_dat_o[26],
    wbs_dat_o[25],
    wbs_dat_o[24],
    wbs_dat_o[23],
    wbs_dat_o[22],
    wbs_dat_o[21],
    wbs_dat_o[20],
    wbs_dat_o[19],
    wbs_dat_o[18],
    wbs_dat_o[17],
    wbs_dat_o[16],
    wbs_dat_o[15],
    wbs_dat_o[14],
    wbs_dat_o[13],
    wbs_dat_o[12],
    wbs_dat_o[11],
    wbs_dat_o[10],
    wbs_dat_o[9],
    wbs_dat_o[8],
    wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 input_mux im (.clk(clk),
    .rst_n(rst_n),
    .vdd(vdd),
    .vss(vss),
    .in({\in[17] ,
    \in[16] ,
    \in[15] ,
    \in[14] ,
    \in[13] ,
    \in[12] ,
    \in[11] ,
    \in[10] ,
    \in[9] ,
    \in[8] ,
    \in[7] ,
    \in[6] ,
    \in[5] ,
    \in[4] ,
    \in[3] ,
    \in[2] ,
    \in[1] ,
    \in[0] }),
    .proj_clk({\proj_clk[7] ,
    \proj_clk[6] ,
    \proj_clk[5] ,
    \proj_clk[4] ,
    \proj_clk[3] ,
    \proj_clk[2] ,
    \proj_clk[1] ,
    \proj_clk[0] }),
    .proj_in({\proj_in[143] ,
    \proj_in[142] ,
    \proj_in[141] ,
    \proj_in[140] ,
    \proj_in[139] ,
    \proj_in[138] ,
    \proj_in[137] ,
    \proj_in[136] ,
    \proj_in[135] ,
    \proj_in[134] ,
    \proj_in[133] ,
    \proj_in[132] ,
    \proj_in[131] ,
    \proj_in[130] ,
    \proj_in[129] ,
    \proj_in[128] ,
    \proj_in[127] ,
    \proj_in[126] ,
    \proj_in[125] ,
    \proj_in[124] ,
    \proj_in[123] ,
    \proj_in[122] ,
    \proj_in[121] ,
    \proj_in[120] ,
    \proj_in[119] ,
    \proj_in[118] ,
    \proj_in[117] ,
    \proj_in[116] ,
    \proj_in[115] ,
    \proj_in[114] ,
    \proj_in[113] ,
    \proj_in[112] ,
    \proj_in[111] ,
    \proj_in[110] ,
    \proj_in[109] ,
    \proj_in[108] ,
    \proj_in[107] ,
    \proj_in[106] ,
    \proj_in[105] ,
    \proj_in[104] ,
    \proj_in[103] ,
    \proj_in[102] ,
    \proj_in[101] ,
    \proj_in[100] ,
    \proj_in[99] ,
    \proj_in[98] ,
    \proj_in[97] ,
    \proj_in[96] ,
    \proj_in[95] ,
    \proj_in[94] ,
    \proj_in[93] ,
    \proj_in[92] ,
    \proj_in[91] ,
    \proj_in[90] ,
    \proj_in[89] ,
    \proj_in[88] ,
    \proj_in[87] ,
    \proj_in[86] ,
    \proj_in[85] ,
    \proj_in[84] ,
    \proj_in[83] ,
    \proj_in[82] ,
    \proj_in[81] ,
    \proj_in[80] ,
    \proj_in[79] ,
    \proj_in[78] ,
    \proj_in[77] ,
    \proj_in[76] ,
    \proj_in[75] ,
    \proj_in[74] ,
    \proj_in[73] ,
    \proj_in[72] ,
    \proj_in[71] ,
    \proj_in[70] ,
    \proj_in[69] ,
    \proj_in[68] ,
    \proj_in[67] ,
    \proj_in[66] ,
    \proj_in[65] ,
    \proj_in[64] ,
    \proj_in[63] ,
    \proj_in[62] ,
    \proj_in[61] ,
    \proj_in[60] ,
    \proj_in[59] ,
    \proj_in[58] ,
    \proj_in[57] ,
    \proj_in[56] ,
    \proj_in[55] ,
    \proj_in[54] ,
    \proj_in[53] ,
    \proj_in[52] ,
    \proj_in[51] ,
    \proj_in[50] ,
    \proj_in[49] ,
    \proj_in[48] ,
    \proj_in[47] ,
    \proj_in[46] ,
    \proj_in[45] ,
    \proj_in[44] ,
    \proj_in[43] ,
    \proj_in[42] ,
    \proj_in[41] ,
    \proj_in[40] ,
    \proj_in[39] ,
    \proj_in[38] ,
    \proj_in[37] ,
    \proj_in[36] ,
    \proj_in[35] ,
    \proj_in[34] ,
    \proj_in[33] ,
    \proj_in[32] ,
    \proj_in[31] ,
    \proj_in[30] ,
    \proj_in[29] ,
    \proj_in[28] ,
    \proj_in[27] ,
    \proj_in[26] ,
    \proj_in[25] ,
    \proj_in[24] ,
    \proj_in[23] ,
    \proj_in[22] ,
    \proj_in[21] ,
    \proj_in[20] ,
    \proj_in[19] ,
    \proj_in[18] ,
    \proj_in[17] ,
    \proj_in[16] ,
    \proj_in[15] ,
    \proj_in[14] ,
    \proj_in[13] ,
    \proj_in[12] ,
    \proj_in[11] ,
    \proj_in[10] ,
    \proj_in[9] ,
    \proj_in[8] ,
    \proj_in[7] ,
    \proj_in[6] ,
    \proj_in[5] ,
    \proj_in[4] ,
    \proj_in[3] ,
    \proj_in[2] ,
    \proj_in[1] ,
    \proj_in[0] }),
    .proj_rst_n({\proj_rst_n[7] ,
    \proj_rst_n[6] ,
    \proj_rst_n[5] ,
    \proj_rst_n[4] ,
    \proj_rst_n[3] ,
    \proj_rst_n[2] ,
    \proj_rst_n[1] ,
    \proj_rst_n[0] }),
    .sel({\sel[2] ,
    \sel[1] ,
    \sel[0] }));
 output_mux om (.vdd(vdd),
    .vss(vss),
    .out({\out[11] ,
    \out[10] ,
    \out[9] ,
    \out[8] ,
    \out[7] ,
    \out[6] ,
    \out[5] ,
    \out[4] ,
    \out[3] ,
    \out[2] ,
    \out[1] ,
    \out[0] }),
    .proj_out({\proj_out[95] ,
    \proj_out[94] ,
    \proj_out[93] ,
    \proj_out[92] ,
    \proj_out[91] ,
    \proj_out[90] ,
    \proj_out[89] ,
    \proj_out[88] ,
    \proj_out[87] ,
    \proj_out[86] ,
    \proj_out[85] ,
    \proj_out[84] ,
    \proj_out[83] ,
    \proj_out[82] ,
    \proj_out[81] ,
    \proj_out[80] ,
    \proj_out[79] ,
    \proj_out[78] ,
    \proj_out[77] ,
    \proj_out[76] ,
    \proj_out[75] ,
    \proj_out[74] ,
    \proj_out[73] ,
    \proj_out[72] ,
    \proj_out[71] ,
    \proj_out[70] ,
    \proj_out[69] ,
    \proj_out[68] ,
    \proj_out[67] ,
    \proj_out[66] ,
    \proj_out[65] ,
    \proj_out[64] ,
    \proj_out[63] ,
    \proj_out[62] ,
    \proj_out[61] ,
    \proj_out[60] ,
    \proj_out[59] ,
    \proj_out[58] ,
    \proj_out[57] ,
    \proj_out[56] ,
    \proj_out[55] ,
    \proj_out[54] ,
    \proj_out[53] ,
    \proj_out[52] ,
    \proj_out[51] ,
    \proj_out[50] ,
    \proj_out[49] ,
    \proj_out[48] ,
    \proj_out[47] ,
    \proj_out[46] ,
    \proj_out[45] ,
    \proj_out[44] ,
    \proj_out[43] ,
    \proj_out[42] ,
    \proj_out[41] ,
    \proj_out[40] ,
    \proj_out[39] ,
    \proj_out[38] ,
    \proj_out[37] ,
    \proj_out[36] ,
    \proj_out[35] ,
    \proj_out[34] ,
    \proj_out[33] ,
    \proj_out[32] ,
    \proj_out[31] ,
    \proj_out[30] ,
    \proj_out[29] ,
    \proj_out[28] ,
    \proj_out[27] ,
    \proj_out[26] ,
    \proj_out[25] ,
    \proj_out[24] ,
    \proj_out[23] ,
    \proj_out[22] ,
    \proj_out[21] ,
    \proj_out[20] ,
    \proj_out[19] ,
    \proj_out[18] ,
    \proj_out[17] ,
    \proj_out[16] ,
    \proj_out[15] ,
    \proj_out[14] ,
    \proj_out[13] ,
    \proj_out[12] ,
    \proj_out[11] ,
    \proj_out[10] ,
    \proj_out[9] ,
    \proj_out[8] ,
    \proj_out[7] ,
    \proj_out[6] ,
    \proj_out[5] ,
    \proj_out[4] ,
    \proj_out[3] ,
    \proj_out[2] ,
    \proj_out[1] ,
    \proj_out[0] }),
    .sel({\sel[2] ,
    \sel[1] ,
    \sel[0] }));
 rotfpga2a p0 (.clk(\proj_clk[0] ),
    .rst_n(\proj_rst_n[0] ),
    .vdd(vdd),
    .vss(vss),
    .in({\proj_in[17] ,
    \proj_in[16] ,
    \proj_in[15] ,
    \proj_in[14] ,
    \proj_in[13] ,
    \proj_in[12] ,
    \proj_in[11] ,
    \proj_in[10] ,
    \proj_in[9] ,
    \proj_in[8] ,
    \proj_in[7] ,
    \proj_in[6] ,
    \proj_in[5] ,
    \proj_in[4] ,
    \proj_in[3] ,
    \proj_in[2] ,
    \proj_in[1] ,
    \proj_in[0] }),
    .out({\proj_out[11] ,
    \proj_out[10] ,
    \proj_out[9] ,
    \proj_out[8] ,
    \proj_out[7] ,
    \proj_out[6] ,
    \proj_out[5] ,
    \proj_out[4] ,
    \proj_out[3] ,
    \proj_out[2] ,
    \proj_out[1] ,
    \proj_out[0] }));
 rotfpga2b p1 (.clk(\proj_clk[1] ),
    .rst_n(\proj_rst_n[1] ),
    .vdd(vdd),
    .vss(vss),
    .in({\proj_in[35] ,
    \proj_in[34] ,
    \proj_in[33] ,
    \proj_in[32] ,
    \proj_in[31] ,
    \proj_in[30] ,
    \proj_in[29] ,
    \proj_in[28] ,
    \proj_in[27] ,
    \proj_in[26] ,
    \proj_in[25] ,
    \proj_in[24] ,
    \proj_in[23] ,
    \proj_in[22] ,
    \proj_in[21] ,
    \proj_in[20] ,
    \proj_in[19] ,
    \proj_in[18] }),
    .out({\proj_out[23] ,
    \proj_out[22] ,
    \proj_out[21] ,
    \proj_out[20] ,
    \proj_out[19] ,
    \proj_out[18] ,
    \proj_out[17] ,
    \proj_out[16] ,
    \proj_out[15] ,
    \proj_out[14] ,
    \proj_out[13] ,
    \proj_out[12] }));
 totp p2 (.clk(\proj_clk[2] ),
    .rst_n(\proj_rst_n[2] ),
    .vdd(vdd),
    .vss(vss),
    .in({\proj_in[53] ,
    \proj_in[52] ,
    \proj_in[51] ,
    \proj_in[50] ,
    \proj_in[49] ,
    \proj_in[48] ,
    \proj_in[47] ,
    \proj_in[46] ,
    \proj_in[45] ,
    \proj_in[44] ,
    \proj_in[43] ,
    \proj_in[42] ,
    \proj_in[41] ,
    \proj_in[40] ,
    \proj_in[39] ,
    \proj_in[38] ,
    \proj_in[37] ,
    \proj_in[36] }),
    .out({\proj_out[35] ,
    \proj_out[34] ,
    \proj_out[33] ,
    \proj_out[32] ,
    \proj_out[31] ,
    \proj_out[30] ,
    \proj_out[29] ,
    \proj_out[28] ,
    \proj_out[27] ,
    \proj_out[26] ,
    \proj_out[25] ,
    \proj_out[24] }));
 unigate p3 (.clk(\proj_clk[3] ),
    .rst_n(\proj_rst_n[3] ),
    .vdd(vdd),
    .vss(vss),
    .in({\proj_in[71] ,
    \proj_in[70] ,
    \proj_in[69] ,
    \proj_in[68] ,
    \proj_in[67] ,
    \proj_in[66] ,
    \proj_in[65] ,
    \proj_in[64] ,
    \proj_in[63] ,
    \proj_in[62] ,
    \proj_in[61] ,
    \proj_in[60] ,
    \proj_in[59] ,
    \proj_in[58] ,
    \proj_in[57] ,
    \proj_in[56] ,
    \proj_in[55] ,
    \proj_in[54] }),
    .out({\proj_out[47] ,
    \proj_out[46] ,
    \proj_out[45] ,
    \proj_out[44] ,
    \proj_out[43] ,
    \proj_out[42] ,
    \proj_out[41] ,
    \proj_out[40] ,
    \proj_out[39] ,
    \proj_out[38] ,
    \proj_out[37] ,
    \proj_out[36] }));
 cells7 p4 (.clk(\proj_clk[4] ),
    .rst_n(\proj_rst_n[4] ),
    .vdd(vdd),
    .vss(vss),
    .in({\proj_in[89] ,
    \proj_in[88] ,
    \proj_in[87] ,
    \proj_in[86] ,
    \proj_in[85] ,
    \proj_in[84] ,
    \proj_in[83] ,
    \proj_in[82] ,
    \proj_in[81] ,
    \proj_in[80] ,
    \proj_in[79] ,
    \proj_in[78] ,
    \proj_in[77] ,
    \proj_in[76] ,
    \proj_in[75] ,
    \proj_in[74] ,
    \proj_in[73] ,
    \proj_in[72] }),
    .out({\proj_out[59] ,
    \proj_out[58] ,
    \proj_out[57] ,
    \proj_out[56] ,
    \proj_out[55] ,
    \proj_out[54] ,
    \proj_out[53] ,
    \proj_out[52] ,
    \proj_out[51] ,
    \proj_out[50] ,
    \proj_out[49] ,
    \proj_out[48] }));
 cells7 p5 (.clk(\proj_clk[3] ),
    .rst_n(\proj_rst_n[3] ),
    .vdd(vdd),
    .vss(vss),
    .in({\proj_in[107] ,
    \proj_in[106] ,
    \proj_in[105] ,
    \proj_in[104] ,
    \proj_in[103] ,
    \proj_in[102] ,
    \proj_in[101] ,
    \proj_in[100] ,
    \proj_in[99] ,
    \proj_in[98] ,
    \proj_in[97] ,
    \proj_in[96] ,
    \proj_in[95] ,
    \proj_in[94] ,
    \proj_in[93] ,
    \proj_in[92] ,
    \proj_in[91] ,
    \proj_in[90] }),
    .out({\proj_out[71] ,
    \proj_out[70] ,
    \proj_out[69] ,
    \proj_out[68] ,
    \proj_out[67] ,
    \proj_out[66] ,
    \proj_out[65] ,
    \proj_out[64] ,
    \proj_out[63] ,
    \proj_out[62] ,
    \proj_out[61] ,
    \proj_out[60] }));
 loopback7 p6 (.clk(\proj_clk[3] ),
    .rst_n(\proj_rst_n[3] ),
    .vdd(vdd),
    .vss(vss),
    .in({\proj_in[125] ,
    \proj_in[124] ,
    \proj_in[123] ,
    \proj_in[122] ,
    \proj_in[121] ,
    \proj_in[120] ,
    \proj_in[119] ,
    \proj_in[118] ,
    \proj_in[117] ,
    \proj_in[116] ,
    \proj_in[115] ,
    \proj_in[114] ,
    \proj_in[113] ,
    \proj_in[112] ,
    \proj_in[111] ,
    \proj_in[110] ,
    \proj_in[109] ,
    \proj_in[108] }),
    .out({\proj_out[83] ,
    \proj_out[82] ,
    \proj_out[81] ,
    \proj_out[80] ,
    \proj_out[79] ,
    \proj_out[78] ,
    \proj_out[77] ,
    \proj_out[76] ,
    \proj_out[75] ,
    \proj_out[74] ,
    \proj_out[73] ,
    \proj_out[72] }));
 loopback7 p7 (.clk(\proj_clk[3] ),
    .rst_n(\proj_rst_n[3] ),
    .vdd(vdd),
    .vss(vss),
    .in({\proj_in[143] ,
    \proj_in[142] ,
    \proj_in[141] ,
    \proj_in[140] ,
    \proj_in[139] ,
    \proj_in[138] ,
    \proj_in[137] ,
    \proj_in[136] ,
    \proj_in[135] ,
    \proj_in[134] ,
    \proj_in[133] ,
    \proj_in[132] ,
    \proj_in[131] ,
    \proj_in[130] ,
    \proj_in[129] ,
    \proj_in[128] ,
    \proj_in[127] ,
    \proj_in[126] }),
    .out({\proj_out[95] ,
    \proj_out[94] ,
    \proj_out[93] ,
    \proj_out[92] ,
    \proj_out[91] ,
    \proj_out[90] ,
    \proj_out[89] ,
    \proj_out[88] ,
    \proj_out[87] ,
    \proj_out[86] ,
    \proj_out[85] ,
    \proj_out[84] }));
endmodule
