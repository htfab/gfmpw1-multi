magic
tech gf180mcuD
magscale 1 10
timestamp 1702353295
<< metal1 >>
rect 1344 36874 38640 36908
rect 1344 36822 5876 36874
rect 5928 36822 5980 36874
rect 6032 36822 6084 36874
rect 6136 36822 15200 36874
rect 15252 36822 15304 36874
rect 15356 36822 15408 36874
rect 15460 36822 24524 36874
rect 24576 36822 24628 36874
rect 24680 36822 24732 36874
rect 24784 36822 33848 36874
rect 33900 36822 33952 36874
rect 34004 36822 34056 36874
rect 34108 36822 38640 36874
rect 1344 36788 38640 36822
rect 21758 36482 21810 36494
rect 35534 36482 35586 36494
rect 14802 36430 14814 36482
rect 14866 36430 14878 36482
rect 17266 36430 17278 36482
rect 17330 36430 17342 36482
rect 21298 36430 21310 36482
rect 21362 36430 21374 36482
rect 24770 36430 24782 36482
rect 24834 36430 24846 36482
rect 26114 36430 26126 36482
rect 26178 36430 26190 36482
rect 21758 36418 21810 36430
rect 35534 36418 35586 36430
rect 37550 36482 37602 36494
rect 37550 36418 37602 36430
rect 15374 36370 15426 36382
rect 15374 36306 15426 36318
rect 15710 36370 15762 36382
rect 15710 36306 15762 36318
rect 16046 36370 16098 36382
rect 16046 36306 16098 36318
rect 16382 36370 16434 36382
rect 16382 36306 16434 36318
rect 17502 36370 17554 36382
rect 17502 36306 17554 36318
rect 17838 36370 17890 36382
rect 17838 36306 17890 36318
rect 18174 36370 18226 36382
rect 18174 36306 18226 36318
rect 18510 36370 18562 36382
rect 18510 36306 18562 36318
rect 18846 36370 18898 36382
rect 18846 36306 18898 36318
rect 19182 36370 19234 36382
rect 19182 36306 19234 36318
rect 19518 36370 19570 36382
rect 19518 36306 19570 36318
rect 19854 36370 19906 36382
rect 19854 36306 19906 36318
rect 20190 36370 20242 36382
rect 20190 36306 20242 36318
rect 21086 36370 21138 36382
rect 21086 36306 21138 36318
rect 22430 36370 22482 36382
rect 22430 36306 22482 36318
rect 22766 36370 22818 36382
rect 22766 36306 22818 36318
rect 23102 36370 23154 36382
rect 23102 36306 23154 36318
rect 23438 36370 23490 36382
rect 23438 36306 23490 36318
rect 24558 36370 24610 36382
rect 24558 36306 24610 36318
rect 25230 36370 25282 36382
rect 25230 36306 25282 36318
rect 25566 36370 25618 36382
rect 25566 36306 25618 36318
rect 36542 36370 36594 36382
rect 36542 36306 36594 36318
rect 36878 36370 36930 36382
rect 36878 36306 36930 36318
rect 22094 36258 22146 36270
rect 36318 36258 36370 36270
rect 38222 36258 38274 36270
rect 15026 36206 15038 36258
rect 15090 36206 15102 36258
rect 25890 36206 25902 36258
rect 25954 36206 25966 36258
rect 37202 36206 37214 36258
rect 37266 36206 37278 36258
rect 37874 36206 37886 36258
rect 37938 36206 37950 36258
rect 22094 36194 22146 36206
rect 36318 36194 36370 36206
rect 38222 36194 38274 36206
rect 1344 36090 38800 36124
rect 1344 36038 10538 36090
rect 10590 36038 10642 36090
rect 10694 36038 10746 36090
rect 10798 36038 19862 36090
rect 19914 36038 19966 36090
rect 20018 36038 20070 36090
rect 20122 36038 29186 36090
rect 29238 36038 29290 36090
rect 29342 36038 29394 36090
rect 29446 36038 38510 36090
rect 38562 36038 38614 36090
rect 38666 36038 38718 36090
rect 38770 36038 38800 36090
rect 1344 36004 38800 36038
rect 15262 35922 15314 35934
rect 15262 35858 15314 35870
rect 16158 35922 16210 35934
rect 16158 35858 16210 35870
rect 16382 35922 16434 35934
rect 16382 35858 16434 35870
rect 21534 35922 21586 35934
rect 21534 35858 21586 35870
rect 25678 35922 25730 35934
rect 25678 35858 25730 35870
rect 37662 35922 37714 35934
rect 37662 35858 37714 35870
rect 38222 35810 38274 35822
rect 16706 35758 16718 35810
rect 16770 35758 16782 35810
rect 38222 35746 38274 35758
rect 37102 35698 37154 35710
rect 37986 35646 37998 35698
rect 38050 35646 38062 35698
rect 37102 35634 37154 35646
rect 1344 35306 38640 35340
rect 1344 35254 5876 35306
rect 5928 35254 5980 35306
rect 6032 35254 6084 35306
rect 6136 35254 15200 35306
rect 15252 35254 15304 35306
rect 15356 35254 15408 35306
rect 15460 35254 24524 35306
rect 24576 35254 24628 35306
rect 24680 35254 24732 35306
rect 24784 35254 33848 35306
rect 33900 35254 33952 35306
rect 34004 35254 34056 35306
rect 34108 35254 38640 35306
rect 1344 35220 38640 35254
rect 37886 34802 37938 34814
rect 37886 34738 37938 34750
rect 38222 34690 38274 34702
rect 38222 34626 38274 34638
rect 1344 34522 38800 34556
rect 1344 34470 10538 34522
rect 10590 34470 10642 34522
rect 10694 34470 10746 34522
rect 10798 34470 19862 34522
rect 19914 34470 19966 34522
rect 20018 34470 20070 34522
rect 20122 34470 29186 34522
rect 29238 34470 29290 34522
rect 29342 34470 29394 34522
rect 29446 34470 38510 34522
rect 38562 34470 38614 34522
rect 38666 34470 38718 34522
rect 38770 34470 38800 34522
rect 1344 34436 38800 34470
rect 38222 34242 38274 34254
rect 38222 34178 38274 34190
rect 37986 34078 37998 34130
rect 38050 34078 38062 34130
rect 37550 34018 37602 34030
rect 37550 33954 37602 33966
rect 1344 33738 38640 33772
rect 1344 33686 5876 33738
rect 5928 33686 5980 33738
rect 6032 33686 6084 33738
rect 6136 33686 15200 33738
rect 15252 33686 15304 33738
rect 15356 33686 15408 33738
rect 15460 33686 24524 33738
rect 24576 33686 24628 33738
rect 24680 33686 24732 33738
rect 24784 33686 33848 33738
rect 33900 33686 33952 33738
rect 34004 33686 34056 33738
rect 34108 33686 38640 33738
rect 1344 33652 38640 33686
rect 37886 33234 37938 33246
rect 37886 33170 37938 33182
rect 38222 33122 38274 33134
rect 38222 33058 38274 33070
rect 1344 32954 38800 32988
rect 1344 32902 10538 32954
rect 10590 32902 10642 32954
rect 10694 32902 10746 32954
rect 10798 32902 19862 32954
rect 19914 32902 19966 32954
rect 20018 32902 20070 32954
rect 20122 32902 29186 32954
rect 29238 32902 29290 32954
rect 29342 32902 29394 32954
rect 29446 32902 38510 32954
rect 38562 32902 38614 32954
rect 38666 32902 38718 32954
rect 38770 32902 38800 32954
rect 1344 32868 38800 32902
rect 37874 32622 37886 32674
rect 37938 32622 37950 32674
rect 38222 32562 38274 32574
rect 38222 32498 38274 32510
rect 37214 32450 37266 32462
rect 37214 32386 37266 32398
rect 37662 32450 37714 32462
rect 37662 32386 37714 32398
rect 1344 32170 38640 32204
rect 1344 32118 5876 32170
rect 5928 32118 5980 32170
rect 6032 32118 6084 32170
rect 6136 32118 15200 32170
rect 15252 32118 15304 32170
rect 15356 32118 15408 32170
rect 15460 32118 24524 32170
rect 24576 32118 24628 32170
rect 24680 32118 24732 32170
rect 24784 32118 33848 32170
rect 33900 32118 33952 32170
rect 34004 32118 34056 32170
rect 34108 32118 38640 32170
rect 1344 32084 38640 32118
rect 37886 31778 37938 31790
rect 37886 31714 37938 31726
rect 37214 31666 37266 31678
rect 37214 31602 37266 31614
rect 37550 31666 37602 31678
rect 37550 31602 37602 31614
rect 36542 31554 36594 31566
rect 36542 31490 36594 31502
rect 38222 31554 38274 31566
rect 38222 31490 38274 31502
rect 1344 31386 38800 31420
rect 1344 31334 10538 31386
rect 10590 31334 10642 31386
rect 10694 31334 10746 31386
rect 10798 31334 19862 31386
rect 19914 31334 19966 31386
rect 20018 31334 20070 31386
rect 20122 31334 29186 31386
rect 29238 31334 29290 31386
rect 29342 31334 29394 31386
rect 29446 31334 38510 31386
rect 38562 31334 38614 31386
rect 38666 31334 38718 31386
rect 38770 31334 38800 31386
rect 1344 31300 38800 31334
rect 38222 31106 38274 31118
rect 38222 31042 38274 31054
rect 37886 30994 37938 31006
rect 37886 30930 37938 30942
rect 37550 30882 37602 30894
rect 37550 30818 37602 30830
rect 1344 30602 38640 30636
rect 1344 30550 5876 30602
rect 5928 30550 5980 30602
rect 6032 30550 6084 30602
rect 6136 30550 15200 30602
rect 15252 30550 15304 30602
rect 15356 30550 15408 30602
rect 15460 30550 24524 30602
rect 24576 30550 24628 30602
rect 24680 30550 24732 30602
rect 24784 30550 33848 30602
rect 33900 30550 33952 30602
rect 34004 30550 34056 30602
rect 34108 30550 38640 30602
rect 1344 30516 38640 30550
rect 37886 30098 37938 30110
rect 37886 30034 37938 30046
rect 37662 29986 37714 29998
rect 37662 29922 37714 29934
rect 38222 29986 38274 29998
rect 38222 29922 38274 29934
rect 1344 29818 38800 29852
rect 1344 29766 10538 29818
rect 10590 29766 10642 29818
rect 10694 29766 10746 29818
rect 10798 29766 19862 29818
rect 19914 29766 19966 29818
rect 20018 29766 20070 29818
rect 20122 29766 29186 29818
rect 29238 29766 29290 29818
rect 29342 29766 29394 29818
rect 29446 29766 38510 29818
rect 38562 29766 38614 29818
rect 38666 29766 38718 29818
rect 38770 29766 38800 29818
rect 1344 29732 38800 29766
rect 38222 29538 38274 29550
rect 38222 29474 38274 29486
rect 37886 29426 37938 29438
rect 37886 29362 37938 29374
rect 1344 29034 38640 29068
rect 1344 28982 5876 29034
rect 5928 28982 5980 29034
rect 6032 28982 6084 29034
rect 6136 28982 15200 29034
rect 15252 28982 15304 29034
rect 15356 28982 15408 29034
rect 15460 28982 24524 29034
rect 24576 28982 24628 29034
rect 24680 28982 24732 29034
rect 24784 28982 33848 29034
rect 33900 28982 33952 29034
rect 34004 28982 34056 29034
rect 34108 28982 38640 29034
rect 1344 28948 38640 28982
rect 37886 28642 37938 28654
rect 37886 28578 37938 28590
rect 37662 28418 37714 28430
rect 37662 28354 37714 28366
rect 38222 28418 38274 28430
rect 38222 28354 38274 28366
rect 1344 28250 38800 28284
rect 1344 28198 10538 28250
rect 10590 28198 10642 28250
rect 10694 28198 10746 28250
rect 10798 28198 19862 28250
rect 19914 28198 19966 28250
rect 20018 28198 20070 28250
rect 20122 28198 29186 28250
rect 29238 28198 29290 28250
rect 29342 28198 29394 28250
rect 29446 28198 38510 28250
rect 38562 28198 38614 28250
rect 38666 28198 38718 28250
rect 38770 28198 38800 28250
rect 1344 28164 38800 28198
rect 38222 27970 38274 27982
rect 38222 27906 38274 27918
rect 37886 27858 37938 27870
rect 37886 27794 37938 27806
rect 1344 27466 38640 27500
rect 1344 27414 5876 27466
rect 5928 27414 5980 27466
rect 6032 27414 6084 27466
rect 6136 27414 15200 27466
rect 15252 27414 15304 27466
rect 15356 27414 15408 27466
rect 15460 27414 24524 27466
rect 24576 27414 24628 27466
rect 24680 27414 24732 27466
rect 24784 27414 33848 27466
rect 33900 27414 33952 27466
rect 34004 27414 34056 27466
rect 34108 27414 38640 27466
rect 1344 27380 38640 27414
rect 37214 27074 37266 27086
rect 1810 27022 1822 27074
rect 1874 27022 1886 27074
rect 37986 27022 37998 27074
rect 38050 27022 38062 27074
rect 37214 27010 37266 27022
rect 2494 26962 2546 26974
rect 2494 26898 2546 26910
rect 37550 26962 37602 26974
rect 37550 26898 37602 26910
rect 38222 26962 38274 26974
rect 38222 26898 38274 26910
rect 2034 26798 2046 26850
rect 2098 26798 2110 26850
rect 1344 26682 38800 26716
rect 1344 26630 10538 26682
rect 10590 26630 10642 26682
rect 10694 26630 10746 26682
rect 10798 26630 19862 26682
rect 19914 26630 19966 26682
rect 20018 26630 20070 26682
rect 20122 26630 29186 26682
rect 29238 26630 29290 26682
rect 29342 26630 29394 26682
rect 29446 26630 38510 26682
rect 38562 26630 38614 26682
rect 38666 26630 38718 26682
rect 38770 26630 38800 26682
rect 1344 26596 38800 26630
rect 22318 26514 22370 26526
rect 22318 26450 22370 26462
rect 1710 26402 1762 26414
rect 1710 26338 1762 26350
rect 37886 26402 37938 26414
rect 37886 26338 37938 26350
rect 2046 26290 2098 26302
rect 2046 26226 2098 26238
rect 38222 26290 38274 26302
rect 38222 26226 38274 26238
rect 2494 26178 2546 26190
rect 2494 26114 2546 26126
rect 37662 26178 37714 26190
rect 37662 26114 37714 26126
rect 2258 26014 2270 26066
rect 2322 26063 2334 26066
rect 2482 26063 2494 26066
rect 2322 26017 2494 26063
rect 2322 26014 2334 26017
rect 2482 26014 2494 26017
rect 2546 26014 2558 26066
rect 1344 25898 38640 25932
rect 1344 25846 5876 25898
rect 5928 25846 5980 25898
rect 6032 25846 6084 25898
rect 6136 25846 15200 25898
rect 15252 25846 15304 25898
rect 15356 25846 15408 25898
rect 15460 25846 24524 25898
rect 24576 25846 24628 25898
rect 24680 25846 24732 25898
rect 24784 25846 33848 25898
rect 33900 25846 33952 25898
rect 34004 25846 34056 25898
rect 34108 25846 38640 25898
rect 1344 25812 38640 25846
rect 37650 25727 37662 25730
rect 37329 25681 37662 25727
rect 21422 25506 21474 25518
rect 23102 25506 23154 25518
rect 1810 25454 1822 25506
rect 1874 25454 1886 25506
rect 19842 25454 19854 25506
rect 19906 25454 19918 25506
rect 22082 25454 22094 25506
rect 22146 25454 22158 25506
rect 25778 25454 25790 25506
rect 25842 25454 25854 25506
rect 26450 25454 26462 25506
rect 26514 25454 26526 25506
rect 28354 25454 28366 25506
rect 28418 25454 28430 25506
rect 21422 25442 21474 25454
rect 23102 25442 23154 25454
rect 17726 25394 17778 25406
rect 17726 25330 17778 25342
rect 18062 25394 18114 25406
rect 18062 25330 18114 25342
rect 19630 25394 19682 25406
rect 19630 25330 19682 25342
rect 21534 25394 21586 25406
rect 21534 25330 21586 25342
rect 21646 25394 21698 25406
rect 21646 25330 21698 25342
rect 22430 25394 22482 25406
rect 22430 25330 22482 25342
rect 22766 25394 22818 25406
rect 22766 25330 22818 25342
rect 23438 25394 23490 25406
rect 23438 25330 23490 25342
rect 26014 25394 26066 25406
rect 26014 25330 26066 25342
rect 26686 25394 26738 25406
rect 26686 25330 26738 25342
rect 28590 25394 28642 25406
rect 28590 25330 28642 25342
rect 29150 25394 29202 25406
rect 29150 25330 29202 25342
rect 29486 25394 29538 25406
rect 29486 25330 29538 25342
rect 2494 25282 2546 25294
rect 2034 25230 2046 25282
rect 2098 25230 2110 25282
rect 2494 25218 2546 25230
rect 19182 25282 19234 25294
rect 19182 25218 19234 25230
rect 27134 25282 27186 25294
rect 37329 25282 37375 25681
rect 37650 25678 37662 25681
rect 37714 25678 37726 25730
rect 37886 25394 37938 25406
rect 37886 25330 37938 25342
rect 37662 25282 37714 25294
rect 37314 25230 37326 25282
rect 37378 25230 37390 25282
rect 27134 25218 27186 25230
rect 37662 25218 37714 25230
rect 38222 25282 38274 25294
rect 38222 25218 38274 25230
rect 1344 25114 38800 25148
rect 1344 25062 10538 25114
rect 10590 25062 10642 25114
rect 10694 25062 10746 25114
rect 10798 25062 19862 25114
rect 19914 25062 19966 25114
rect 20018 25062 20070 25114
rect 20122 25062 29186 25114
rect 29238 25062 29290 25114
rect 29342 25062 29394 25114
rect 29446 25062 38510 25114
rect 38562 25062 38614 25114
rect 38666 25062 38718 25114
rect 38770 25062 38800 25114
rect 1344 25028 38800 25062
rect 17726 24946 17778 24958
rect 20190 24946 20242 24958
rect 22206 24946 22258 24958
rect 18946 24894 18958 24946
rect 19010 24894 19022 24946
rect 21746 24894 21758 24946
rect 21810 24894 21822 24946
rect 17726 24882 17778 24894
rect 20190 24882 20242 24894
rect 22206 24882 22258 24894
rect 23438 24946 23490 24958
rect 23438 24882 23490 24894
rect 24110 24946 24162 24958
rect 27134 24946 27186 24958
rect 30158 24946 30210 24958
rect 25778 24894 25790 24946
rect 25842 24894 25854 24946
rect 26674 24894 26686 24946
rect 26738 24894 26750 24946
rect 28354 24894 28366 24946
rect 28418 24894 28430 24946
rect 29250 24894 29262 24946
rect 29314 24894 29326 24946
rect 24110 24882 24162 24894
rect 27134 24882 27186 24894
rect 30158 24882 30210 24894
rect 1710 24834 1762 24846
rect 1710 24770 1762 24782
rect 21086 24834 21138 24846
rect 21086 24770 21138 24782
rect 21310 24834 21362 24846
rect 21310 24770 21362 24782
rect 38222 24834 38274 24846
rect 38222 24770 38274 24782
rect 2046 24722 2098 24734
rect 18398 24722 18450 24734
rect 17938 24670 17950 24722
rect 18002 24670 18014 24722
rect 2046 24658 2098 24670
rect 18398 24658 18450 24670
rect 19294 24722 19346 24734
rect 20526 24722 20578 24734
rect 19842 24670 19854 24722
rect 19906 24670 19918 24722
rect 19294 24658 19346 24670
rect 20526 24658 20578 24670
rect 21198 24722 21250 24734
rect 21198 24658 21250 24670
rect 23102 24722 23154 24734
rect 23102 24658 23154 24670
rect 23774 24722 23826 24734
rect 23774 24658 23826 24670
rect 26126 24722 26178 24734
rect 26126 24658 26178 24670
rect 27806 24722 27858 24734
rect 27806 24658 27858 24670
rect 28702 24722 28754 24734
rect 28702 24658 28754 24670
rect 29710 24722 29762 24734
rect 37986 24670 37998 24722
rect 38050 24670 38062 24722
rect 29710 24658 29762 24670
rect 2494 24610 2546 24622
rect 2494 24546 2546 24558
rect 25230 24610 25282 24622
rect 25230 24546 25282 24558
rect 18622 24498 18674 24510
rect 18622 24434 18674 24446
rect 19518 24498 19570 24510
rect 19518 24434 19570 24446
rect 25454 24498 25506 24510
rect 25454 24434 25506 24446
rect 26350 24498 26402 24510
rect 26350 24434 26402 24446
rect 28030 24498 28082 24510
rect 28030 24434 28082 24446
rect 28926 24498 28978 24510
rect 28926 24434 28978 24446
rect 1344 24330 38640 24364
rect 1344 24278 5876 24330
rect 5928 24278 5980 24330
rect 6032 24278 6084 24330
rect 6136 24278 15200 24330
rect 15252 24278 15304 24330
rect 15356 24278 15408 24330
rect 15460 24278 24524 24330
rect 24576 24278 24628 24330
rect 24680 24278 24732 24330
rect 24784 24278 33848 24330
rect 33900 24278 33952 24330
rect 34004 24278 34056 24330
rect 34108 24278 38640 24330
rect 1344 24244 38640 24278
rect 17614 24162 17666 24174
rect 18622 24162 18674 24174
rect 24670 24162 24722 24174
rect 17938 24110 17950 24162
rect 18002 24110 18014 24162
rect 18274 24110 18286 24162
rect 18338 24110 18350 24162
rect 22530 24110 22542 24162
rect 22594 24110 22606 24162
rect 17614 24098 17666 24110
rect 18622 24098 18674 24110
rect 24670 24098 24722 24110
rect 26014 24162 26066 24174
rect 26014 24098 26066 24110
rect 27582 24162 27634 24174
rect 27582 24098 27634 24110
rect 29374 24162 29426 24174
rect 29374 24098 29426 24110
rect 16606 24050 16658 24062
rect 16606 23986 16658 23998
rect 17054 24050 17106 24062
rect 17054 23986 17106 23998
rect 17390 24050 17442 24062
rect 17390 23986 17442 23998
rect 20078 24050 20130 24062
rect 20078 23986 20130 23998
rect 29150 24050 29202 24062
rect 29150 23986 29202 23998
rect 18846 23938 18898 23950
rect 22094 23938 22146 23950
rect 24894 23938 24946 23950
rect 19506 23886 19518 23938
rect 19570 23886 19582 23938
rect 23762 23886 23774 23938
rect 23826 23886 23838 23938
rect 18846 23874 18898 23886
rect 22094 23874 22146 23886
rect 24894 23874 24946 23886
rect 25790 23938 25842 23950
rect 25790 23874 25842 23886
rect 27358 23938 27410 23950
rect 27358 23874 27410 23886
rect 2046 23826 2098 23838
rect 2046 23762 2098 23774
rect 19294 23826 19346 23838
rect 19294 23762 19346 23774
rect 21870 23826 21922 23838
rect 21870 23762 21922 23774
rect 21982 23826 22034 23838
rect 21982 23762 22034 23774
rect 23998 23826 24050 23838
rect 23998 23762 24050 23774
rect 25342 23826 25394 23838
rect 26686 23826 26738 23838
rect 26338 23774 26350 23826
rect 26402 23774 26414 23826
rect 25342 23762 25394 23774
rect 26686 23762 26738 23774
rect 27022 23826 27074 23838
rect 28254 23826 28306 23838
rect 27906 23774 27918 23826
rect 27970 23774 27982 23826
rect 27022 23762 27074 23774
rect 28254 23762 28306 23774
rect 28590 23826 28642 23838
rect 30046 23826 30098 23838
rect 29698 23774 29710 23826
rect 29762 23774 29774 23826
rect 28590 23762 28642 23774
rect 30046 23762 30098 23774
rect 30382 23826 30434 23838
rect 30382 23762 30434 23774
rect 37886 23826 37938 23838
rect 37886 23762 37938 23774
rect 1710 23714 1762 23726
rect 1710 23650 1762 23662
rect 21422 23714 21474 23726
rect 38222 23714 38274 23726
rect 24322 23662 24334 23714
rect 24386 23662 24398 23714
rect 21422 23650 21474 23662
rect 38222 23650 38274 23662
rect 1344 23546 38800 23580
rect 1344 23494 10538 23546
rect 10590 23494 10642 23546
rect 10694 23494 10746 23546
rect 10798 23494 19862 23546
rect 19914 23494 19966 23546
rect 20018 23494 20070 23546
rect 20122 23494 29186 23546
rect 29238 23494 29290 23546
rect 29342 23494 29394 23546
rect 29446 23494 38510 23546
rect 38562 23494 38614 23546
rect 38666 23494 38718 23546
rect 38770 23494 38800 23546
rect 1344 23460 38800 23494
rect 17726 23378 17778 23390
rect 23886 23378 23938 23390
rect 22530 23326 22542 23378
rect 22594 23326 22606 23378
rect 17726 23314 17778 23326
rect 23886 23314 23938 23326
rect 25566 23378 25618 23390
rect 25566 23314 25618 23326
rect 26014 23378 26066 23390
rect 26014 23314 26066 23326
rect 28142 23378 28194 23390
rect 28142 23314 28194 23326
rect 30158 23378 30210 23390
rect 30158 23314 30210 23326
rect 1710 23266 1762 23278
rect 1710 23202 1762 23214
rect 19742 23266 19794 23278
rect 19742 23202 19794 23214
rect 20414 23266 20466 23278
rect 20414 23202 20466 23214
rect 21086 23266 21138 23278
rect 21086 23202 21138 23214
rect 22094 23266 22146 23278
rect 22094 23202 22146 23214
rect 23214 23266 23266 23278
rect 23214 23202 23266 23214
rect 28926 23266 28978 23278
rect 28926 23202 28978 23214
rect 38222 23266 38274 23278
rect 38222 23202 38274 23214
rect 2046 23154 2098 23166
rect 2046 23090 2098 23102
rect 18062 23154 18114 23166
rect 18062 23090 18114 23102
rect 19406 23154 19458 23166
rect 21982 23154 22034 23166
rect 20178 23102 20190 23154
rect 20242 23102 20254 23154
rect 20850 23102 20862 23154
rect 20914 23102 20926 23154
rect 21746 23102 21758 23154
rect 21810 23102 21822 23154
rect 19406 23090 19458 23102
rect 21982 23090 22034 23102
rect 22878 23154 22930 23166
rect 22878 23090 22930 23102
rect 23550 23154 23602 23166
rect 37886 23154 37938 23166
rect 25330 23102 25342 23154
rect 25394 23102 25406 23154
rect 28354 23102 28366 23154
rect 28418 23102 28430 23154
rect 23550 23090 23602 23102
rect 37886 23090 37938 23102
rect 1344 22762 38640 22796
rect 1344 22710 5876 22762
rect 5928 22710 5980 22762
rect 6032 22710 6084 22762
rect 6136 22710 15200 22762
rect 15252 22710 15304 22762
rect 15356 22710 15408 22762
rect 15460 22710 24524 22762
rect 24576 22710 24628 22762
rect 24680 22710 24732 22762
rect 24784 22710 33848 22762
rect 33900 22710 33952 22762
rect 34004 22710 34056 22762
rect 34108 22710 38640 22762
rect 1344 22676 38640 22710
rect 18274 22542 18286 22594
rect 18338 22542 18350 22594
rect 19282 22542 19294 22594
rect 19346 22542 19358 22594
rect 22418 22542 22430 22594
rect 22482 22542 22494 22594
rect 16718 22482 16770 22494
rect 16718 22418 16770 22430
rect 17054 22482 17106 22494
rect 17054 22418 17106 22430
rect 17390 22482 17442 22494
rect 17390 22418 17442 22430
rect 18846 22482 18898 22494
rect 18846 22418 18898 22430
rect 19854 22482 19906 22494
rect 19854 22418 19906 22430
rect 20302 22482 20354 22494
rect 20302 22418 20354 22430
rect 20750 22482 20802 22494
rect 20750 22418 20802 22430
rect 17614 22370 17666 22382
rect 17614 22306 17666 22318
rect 18622 22370 18674 22382
rect 18622 22306 18674 22318
rect 19630 22370 19682 22382
rect 25118 22370 25170 22382
rect 21634 22318 21646 22370
rect 21698 22318 21710 22370
rect 19630 22306 19682 22318
rect 25118 22306 25170 22318
rect 26238 22370 26290 22382
rect 26238 22306 26290 22318
rect 29374 22370 29426 22382
rect 29374 22306 29426 22318
rect 1710 22258 1762 22270
rect 1710 22194 1762 22206
rect 2046 22258 2098 22270
rect 2046 22194 2098 22206
rect 2718 22258 2770 22270
rect 2718 22194 2770 22206
rect 21870 22258 21922 22270
rect 21870 22194 21922 22206
rect 21982 22258 22034 22270
rect 21982 22194 22034 22206
rect 25230 22258 25282 22270
rect 25230 22194 25282 22206
rect 25342 22258 25394 22270
rect 25342 22194 25394 22206
rect 26350 22258 26402 22270
rect 26350 22194 26402 22206
rect 26462 22258 26514 22270
rect 27246 22258 27298 22270
rect 26898 22206 26910 22258
rect 26962 22206 26974 22258
rect 26462 22194 26514 22206
rect 27246 22194 27298 22206
rect 27582 22258 27634 22270
rect 27582 22194 27634 22206
rect 29262 22258 29314 22270
rect 29262 22194 29314 22206
rect 29486 22258 29538 22270
rect 30270 22258 30322 22270
rect 29922 22206 29934 22258
rect 29986 22206 29998 22258
rect 29486 22194 29538 22206
rect 30270 22194 30322 22206
rect 30606 22258 30658 22270
rect 30606 22194 30658 22206
rect 30942 22258 30994 22270
rect 30942 22194 30994 22206
rect 31278 22258 31330 22270
rect 31278 22194 31330 22206
rect 37214 22258 37266 22270
rect 37214 22194 37266 22206
rect 37886 22258 37938 22270
rect 37886 22194 37938 22206
rect 38222 22258 38274 22270
rect 38222 22194 38274 22206
rect 2382 22146 2434 22158
rect 37550 22146 37602 22158
rect 17938 22094 17950 22146
rect 18002 22094 18014 22146
rect 25778 22094 25790 22146
rect 25842 22094 25854 22146
rect 2382 22082 2434 22094
rect 37550 22082 37602 22094
rect 1344 21978 38800 22012
rect 1344 21926 10538 21978
rect 10590 21926 10642 21978
rect 10694 21926 10746 21978
rect 10798 21926 19862 21978
rect 19914 21926 19966 21978
rect 20018 21926 20070 21978
rect 20122 21926 29186 21978
rect 29238 21926 29290 21978
rect 29342 21926 29394 21978
rect 29446 21926 38510 21978
rect 38562 21926 38614 21978
rect 38666 21926 38718 21978
rect 38770 21926 38800 21978
rect 1344 21892 38800 21926
rect 14702 21810 14754 21822
rect 14702 21746 14754 21758
rect 15374 21810 15426 21822
rect 15374 21746 15426 21758
rect 17726 21810 17778 21822
rect 17726 21746 17778 21758
rect 18846 21810 18898 21822
rect 18846 21746 18898 21758
rect 20078 21810 20130 21822
rect 20078 21746 20130 21758
rect 20974 21810 21026 21822
rect 20974 21746 21026 21758
rect 21422 21810 21474 21822
rect 23102 21810 23154 21822
rect 22418 21758 22430 21810
rect 22482 21758 22494 21810
rect 21422 21746 21474 21758
rect 23102 21746 23154 21758
rect 26126 21810 26178 21822
rect 26126 21746 26178 21758
rect 28478 21810 28530 21822
rect 30270 21810 30322 21822
rect 29586 21758 29598 21810
rect 29650 21758 29662 21810
rect 28478 21746 28530 21758
rect 30270 21746 30322 21758
rect 1710 21698 1762 21710
rect 1710 21634 1762 21646
rect 12350 21698 12402 21710
rect 12350 21634 12402 21646
rect 21758 21698 21810 21710
rect 21758 21634 21810 21646
rect 21870 21698 21922 21710
rect 21870 21634 21922 21646
rect 21982 21698 22034 21710
rect 21982 21634 22034 21646
rect 24446 21698 24498 21710
rect 24446 21634 24498 21646
rect 25790 21698 25842 21710
rect 25790 21634 25842 21646
rect 26798 21698 26850 21710
rect 26798 21634 26850 21646
rect 27246 21698 27298 21710
rect 27246 21634 27298 21646
rect 27470 21698 27522 21710
rect 27470 21634 27522 21646
rect 29038 21698 29090 21710
rect 29038 21634 29090 21646
rect 29150 21698 29202 21710
rect 29150 21634 29202 21646
rect 38222 21698 38274 21710
rect 38222 21634 38274 21646
rect 2046 21586 2098 21598
rect 18510 21586 18562 21598
rect 12562 21534 12574 21586
rect 12626 21534 12638 21586
rect 14914 21534 14926 21586
rect 14978 21534 14990 21586
rect 15586 21534 15598 21586
rect 15650 21534 15662 21586
rect 17938 21534 17950 21586
rect 18002 21534 18014 21586
rect 2046 21522 2098 21534
rect 18510 21522 18562 21534
rect 19182 21586 19234 21598
rect 19182 21522 19234 21534
rect 19406 21586 19458 21598
rect 22766 21586 22818 21598
rect 20290 21534 20302 21586
rect 20354 21534 20366 21586
rect 19406 21522 19458 21534
rect 22766 21522 22818 21534
rect 24334 21586 24386 21598
rect 26462 21586 26514 21598
rect 24658 21534 24670 21586
rect 24722 21534 24734 21586
rect 24334 21522 24386 21534
rect 26462 21522 26514 21534
rect 27358 21586 27410 21598
rect 29934 21586 29986 21598
rect 28802 21534 28814 21586
rect 28866 21534 28878 21586
rect 27358 21522 27410 21534
rect 29934 21522 29986 21534
rect 37886 21586 37938 21598
rect 37886 21522 37938 21534
rect 25454 21474 25506 21486
rect 19730 21422 19742 21474
rect 19794 21422 19806 21474
rect 25454 21410 25506 21422
rect 23874 21310 23886 21362
rect 23938 21310 23950 21362
rect 27906 21310 27918 21362
rect 27970 21310 27982 21362
rect 1344 21194 38640 21228
rect 1344 21142 5876 21194
rect 5928 21142 5980 21194
rect 6032 21142 6084 21194
rect 6136 21142 15200 21194
rect 15252 21142 15304 21194
rect 15356 21142 15408 21194
rect 15460 21142 24524 21194
rect 24576 21142 24628 21194
rect 24680 21142 24732 21194
rect 24784 21142 33848 21194
rect 33900 21142 33952 21194
rect 34004 21142 34056 21194
rect 34108 21142 38640 21194
rect 1344 21108 38640 21142
rect 12338 20974 12350 21026
rect 12402 20974 12414 21026
rect 14690 20974 14702 21026
rect 14754 20974 14766 21026
rect 22194 20974 22206 21026
rect 22258 20974 22270 21026
rect 29922 20974 29934 21026
rect 29986 20974 29998 21026
rect 15822 20914 15874 20926
rect 15822 20850 15874 20862
rect 30382 20914 30434 20926
rect 30382 20850 30434 20862
rect 11790 20802 11842 20814
rect 11790 20738 11842 20750
rect 12014 20802 12066 20814
rect 21646 20802 21698 20814
rect 13906 20750 13918 20802
rect 13970 20750 13982 20802
rect 16930 20750 16942 20802
rect 16994 20750 17006 20802
rect 17490 20750 17502 20802
rect 17554 20750 17566 20802
rect 18162 20750 18174 20802
rect 18226 20750 18238 20802
rect 19058 20750 19070 20802
rect 19122 20750 19134 20802
rect 21410 20750 21422 20802
rect 21474 20750 21486 20802
rect 12014 20738 12066 20750
rect 21646 20738 21698 20750
rect 21758 20802 21810 20814
rect 24110 20802 24162 20814
rect 22754 20750 22766 20802
rect 22818 20750 22830 20802
rect 21758 20738 21810 20750
rect 24110 20738 24162 20750
rect 25454 20802 25506 20814
rect 25454 20738 25506 20750
rect 25566 20802 25618 20814
rect 29262 20802 29314 20814
rect 27906 20750 27918 20802
rect 27970 20750 27982 20802
rect 25566 20738 25618 20750
rect 29262 20738 29314 20750
rect 29374 20802 29426 20814
rect 29374 20738 29426 20750
rect 29486 20802 29538 20814
rect 37986 20750 37998 20802
rect 38050 20750 38062 20802
rect 29486 20738 29538 20750
rect 2046 20690 2098 20702
rect 2046 20626 2098 20638
rect 11118 20690 11170 20702
rect 11118 20626 11170 20638
rect 11454 20690 11506 20702
rect 11454 20626 11506 20638
rect 14142 20690 14194 20702
rect 14142 20626 14194 20638
rect 14254 20690 14306 20702
rect 14254 20626 14306 20638
rect 16270 20690 16322 20702
rect 16270 20626 16322 20638
rect 16382 20690 16434 20702
rect 16382 20626 16434 20638
rect 16494 20690 16546 20702
rect 16494 20626 16546 20638
rect 17950 20690 18002 20702
rect 17950 20626 18002 20638
rect 18846 20690 18898 20702
rect 20414 20690 20466 20702
rect 19954 20638 19966 20690
rect 20018 20638 20030 20690
rect 18846 20626 18898 20638
rect 20414 20626 20466 20638
rect 22542 20690 22594 20702
rect 22542 20626 22594 20638
rect 23214 20690 23266 20702
rect 23214 20626 23266 20638
rect 23550 20690 23602 20702
rect 23550 20626 23602 20638
rect 24446 20690 24498 20702
rect 24446 20626 24498 20638
rect 25342 20690 25394 20702
rect 26350 20690 26402 20702
rect 26002 20638 26014 20690
rect 26066 20638 26078 20690
rect 25342 20626 25394 20638
rect 26350 20626 26402 20638
rect 27022 20690 27074 20702
rect 27022 20626 27074 20638
rect 27358 20690 27410 20702
rect 27358 20626 27410 20638
rect 28142 20690 28194 20702
rect 28142 20626 28194 20638
rect 1710 20578 1762 20590
rect 1710 20514 1762 20526
rect 10782 20578 10834 20590
rect 10782 20514 10834 20526
rect 13582 20578 13634 20590
rect 13582 20514 13634 20526
rect 17278 20578 17330 20590
rect 17278 20514 17330 20526
rect 19630 20578 19682 20590
rect 19630 20514 19682 20526
rect 20750 20578 20802 20590
rect 20750 20514 20802 20526
rect 26686 20578 26738 20590
rect 26686 20514 26738 20526
rect 38222 20578 38274 20590
rect 38222 20514 38274 20526
rect 1344 20410 38800 20444
rect 1344 20358 10538 20410
rect 10590 20358 10642 20410
rect 10694 20358 10746 20410
rect 10798 20358 19862 20410
rect 19914 20358 19966 20410
rect 20018 20358 20070 20410
rect 20122 20358 29186 20410
rect 29238 20358 29290 20410
rect 29342 20358 29394 20410
rect 29446 20358 38510 20410
rect 38562 20358 38614 20410
rect 38666 20358 38718 20410
rect 38770 20358 38800 20410
rect 1344 20324 38800 20358
rect 16158 20242 16210 20254
rect 18510 20242 18562 20254
rect 11554 20190 11566 20242
rect 11618 20190 11630 20242
rect 17938 20190 17950 20242
rect 18002 20190 18014 20242
rect 16158 20178 16210 20190
rect 18510 20178 18562 20190
rect 20526 20242 20578 20254
rect 23662 20242 23714 20254
rect 22194 20190 22206 20242
rect 22258 20190 22270 20242
rect 20526 20178 20578 20190
rect 23662 20178 23714 20190
rect 24334 20242 24386 20254
rect 24334 20178 24386 20190
rect 25790 20242 25842 20254
rect 25790 20178 25842 20190
rect 1710 20130 1762 20142
rect 1710 20066 1762 20078
rect 10782 20130 10834 20142
rect 10782 20066 10834 20078
rect 14142 20130 14194 20142
rect 14142 20066 14194 20078
rect 14254 20130 14306 20142
rect 15262 20130 15314 20142
rect 14690 20078 14702 20130
rect 14754 20078 14766 20130
rect 14254 20066 14306 20078
rect 15262 20066 15314 20078
rect 15374 20130 15426 20142
rect 19966 20130 20018 20142
rect 19170 20078 19182 20130
rect 19234 20078 19246 20130
rect 15374 20066 15426 20078
rect 19966 20066 20018 20078
rect 21534 20130 21586 20142
rect 21534 20066 21586 20078
rect 21646 20130 21698 20142
rect 21646 20066 21698 20078
rect 21758 20130 21810 20142
rect 21758 20066 21810 20078
rect 23998 20130 24050 20142
rect 23998 20066 24050 20078
rect 26350 20130 26402 20142
rect 26350 20066 26402 20078
rect 26686 20130 26738 20142
rect 26686 20066 26738 20078
rect 27022 20130 27074 20142
rect 27022 20066 27074 20078
rect 28254 20130 28306 20142
rect 28254 20066 28306 20078
rect 28926 20130 28978 20142
rect 28926 20066 28978 20078
rect 30382 20130 30434 20142
rect 30382 20066 30434 20078
rect 37886 20130 37938 20142
rect 37886 20066 37938 20078
rect 38222 20130 38274 20142
rect 38222 20066 38274 20078
rect 2046 20018 2098 20030
rect 2046 19954 2098 19966
rect 12126 20018 12178 20030
rect 12126 19954 12178 19966
rect 14030 20018 14082 20030
rect 16494 20018 16546 20030
rect 19630 20018 19682 20030
rect 15026 19966 15038 20018
rect 15090 19966 15102 20018
rect 18946 19966 18958 20018
rect 19010 19966 19022 20018
rect 14030 19954 14082 19966
rect 16494 19954 16546 19966
rect 19630 19954 19682 19966
rect 22654 20018 22706 20030
rect 26014 20018 26066 20030
rect 23426 19966 23438 20018
rect 23490 19966 23502 20018
rect 22654 19954 22706 19966
rect 26014 19954 26066 19966
rect 27918 20018 27970 20030
rect 27918 19954 27970 19966
rect 28590 20018 28642 20030
rect 28590 19954 28642 19966
rect 30046 20018 30098 20030
rect 30046 19954 30098 19966
rect 11230 19906 11282 19918
rect 11230 19842 11282 19854
rect 13022 19906 13074 19918
rect 13022 19842 13074 19854
rect 13582 19906 13634 19918
rect 13582 19842 13634 19854
rect 17390 19906 17442 19918
rect 17390 19842 17442 19854
rect 18398 19906 18450 19918
rect 18398 19842 18450 19854
rect 30942 19906 30994 19918
rect 30942 19842 30994 19854
rect 11902 19794 11954 19806
rect 12798 19794 12850 19806
rect 17614 19794 17666 19806
rect 12450 19742 12462 19794
rect 12514 19742 12526 19794
rect 15810 19742 15822 19794
rect 15874 19742 15886 19794
rect 11902 19730 11954 19742
rect 12798 19730 12850 19742
rect 17614 19730 17666 19742
rect 1344 19626 38640 19660
rect 1344 19574 5876 19626
rect 5928 19574 5980 19626
rect 6032 19574 6084 19626
rect 6136 19574 15200 19626
rect 15252 19574 15304 19626
rect 15356 19574 15408 19626
rect 15460 19574 24524 19626
rect 24576 19574 24628 19626
rect 24680 19574 24732 19626
rect 24784 19574 33848 19626
rect 33900 19574 33952 19626
rect 34004 19574 34056 19626
rect 34108 19574 38640 19626
rect 1344 19540 38640 19574
rect 27906 19406 27918 19458
rect 27970 19406 27982 19458
rect 30034 19406 30046 19458
rect 30098 19406 30110 19458
rect 11566 19346 11618 19358
rect 11566 19282 11618 19294
rect 13582 19346 13634 19358
rect 13582 19282 13634 19294
rect 18958 19346 19010 19358
rect 18958 19282 19010 19294
rect 22542 19346 22594 19358
rect 22542 19282 22594 19294
rect 2046 19234 2098 19246
rect 2046 19170 2098 19182
rect 12238 19234 12290 19246
rect 15262 19234 15314 19246
rect 18510 19234 18562 19246
rect 26014 19234 26066 19246
rect 12786 19182 12798 19234
rect 12850 19182 12862 19234
rect 17154 19182 17166 19234
rect 17218 19182 17230 19234
rect 20626 19182 20638 19234
rect 20690 19182 20702 19234
rect 22866 19182 22878 19234
rect 22930 19182 22942 19234
rect 12238 19170 12290 19182
rect 15262 19170 15314 19182
rect 18510 19170 18562 19182
rect 26014 19170 26066 19182
rect 27470 19234 27522 19246
rect 27470 19170 27522 19182
rect 29374 19234 29426 19246
rect 37886 19234 37938 19246
rect 30370 19182 30382 19234
rect 30434 19182 30446 19234
rect 29374 19170 29426 19182
rect 37886 19170 37938 19182
rect 11902 19122 11954 19134
rect 11902 19058 11954 19070
rect 14926 19122 14978 19134
rect 14926 19058 14978 19070
rect 15934 19122 15986 19134
rect 15934 19058 15986 19070
rect 18174 19122 18226 19134
rect 18174 19058 18226 19070
rect 18846 19122 18898 19134
rect 18846 19058 18898 19070
rect 19742 19122 19794 19134
rect 19742 19058 19794 19070
rect 21534 19122 21586 19134
rect 21534 19058 21586 19070
rect 21870 19122 21922 19134
rect 21870 19058 21922 19070
rect 23102 19122 23154 19134
rect 23102 19058 23154 19070
rect 23214 19122 23266 19134
rect 23214 19058 23266 19070
rect 23998 19122 24050 19134
rect 23998 19058 24050 19070
rect 24334 19122 24386 19134
rect 24334 19058 24386 19070
rect 24670 19122 24722 19134
rect 24670 19058 24722 19070
rect 25342 19122 25394 19134
rect 25342 19058 25394 19070
rect 27246 19122 27298 19134
rect 27246 19058 27298 19070
rect 27358 19122 27410 19134
rect 27358 19058 27410 19070
rect 29486 19122 29538 19134
rect 29486 19058 29538 19070
rect 29598 19122 29650 19134
rect 29598 19058 29650 19070
rect 30606 19122 30658 19134
rect 30606 19058 30658 19070
rect 30718 19122 30770 19134
rect 31502 19122 31554 19134
rect 31154 19070 31166 19122
rect 31218 19070 31230 19122
rect 30718 19058 30770 19070
rect 31502 19058 31554 19070
rect 1710 19010 1762 19022
rect 1710 18946 1762 18958
rect 12574 19010 12626 19022
rect 12574 18946 12626 18958
rect 15598 19010 15650 19022
rect 15598 18946 15650 18958
rect 16942 19010 16994 19022
rect 16942 18946 16994 18958
rect 17726 19010 17778 19022
rect 17726 18946 17778 18958
rect 19070 19010 19122 19022
rect 19070 18946 19122 18958
rect 20078 19010 20130 19022
rect 20078 18946 20130 18958
rect 20414 19010 20466 19022
rect 25006 19010 25058 19022
rect 23650 18958 23662 19010
rect 23714 18958 23726 19010
rect 20414 18946 20466 18958
rect 25006 18946 25058 18958
rect 25678 19010 25730 19022
rect 25678 18946 25730 18958
rect 26350 19010 26402 19022
rect 26350 18946 26402 18958
rect 28366 19010 28418 19022
rect 28366 18946 28418 18958
rect 31838 19010 31890 19022
rect 31838 18946 31890 18958
rect 32398 19010 32450 19022
rect 32398 18946 32450 18958
rect 38222 19010 38274 19022
rect 38222 18946 38274 18958
rect 1344 18842 38800 18876
rect 1344 18790 10538 18842
rect 10590 18790 10642 18842
rect 10694 18790 10746 18842
rect 10798 18790 19862 18842
rect 19914 18790 19966 18842
rect 20018 18790 20070 18842
rect 20122 18790 29186 18842
rect 29238 18790 29290 18842
rect 29342 18790 29394 18842
rect 29446 18790 38510 18842
rect 38562 18790 38614 18842
rect 38666 18790 38718 18842
rect 38770 18790 38800 18842
rect 1344 18756 38800 18790
rect 13470 18674 13522 18686
rect 23438 18674 23490 18686
rect 12450 18622 12462 18674
rect 12514 18622 12526 18674
rect 16818 18622 16830 18674
rect 16882 18622 16894 18674
rect 19170 18622 19182 18674
rect 19234 18622 19246 18674
rect 21522 18622 21534 18674
rect 21586 18622 21598 18674
rect 13470 18610 13522 18622
rect 23438 18610 23490 18622
rect 1710 18562 1762 18574
rect 1710 18498 1762 18510
rect 10894 18562 10946 18574
rect 10894 18498 10946 18510
rect 13918 18562 13970 18574
rect 13918 18498 13970 18510
rect 15374 18562 15426 18574
rect 15374 18498 15426 18510
rect 18174 18562 18226 18574
rect 18174 18498 18226 18510
rect 19854 18562 19906 18574
rect 19854 18498 19906 18510
rect 20974 18562 21026 18574
rect 20974 18498 21026 18510
rect 24446 18562 24498 18574
rect 24446 18498 24498 18510
rect 26574 18562 26626 18574
rect 26574 18498 26626 18510
rect 27470 18562 27522 18574
rect 27470 18498 27522 18510
rect 28926 18562 28978 18574
rect 28926 18498 28978 18510
rect 29038 18562 29090 18574
rect 29038 18498 29090 18510
rect 30046 18562 30098 18574
rect 30046 18498 30098 18510
rect 30158 18562 30210 18574
rect 30158 18498 30210 18510
rect 31278 18562 31330 18574
rect 31278 18498 31330 18510
rect 38222 18562 38274 18574
rect 38222 18498 38274 18510
rect 2046 18450 2098 18462
rect 2046 18386 2098 18398
rect 10558 18450 10610 18462
rect 10558 18386 10610 18398
rect 11230 18450 11282 18462
rect 12126 18450 12178 18462
rect 11554 18398 11566 18450
rect 11618 18398 11630 18450
rect 11230 18386 11282 18398
rect 12126 18386 12178 18398
rect 13022 18450 13074 18462
rect 13022 18386 13074 18398
rect 14030 18450 14082 18462
rect 14030 18386 14082 18398
rect 14142 18450 14194 18462
rect 15710 18450 15762 18462
rect 16270 18450 16322 18462
rect 14578 18398 14590 18450
rect 14642 18398 14654 18450
rect 16034 18398 16046 18450
rect 16098 18398 16110 18450
rect 14142 18386 14194 18398
rect 15710 18386 15762 18398
rect 16270 18386 16322 18398
rect 16382 18450 16434 18462
rect 16382 18386 16434 18398
rect 17838 18450 17890 18462
rect 17838 18386 17890 18398
rect 18510 18450 18562 18462
rect 18510 18386 18562 18398
rect 18846 18450 18898 18462
rect 18846 18386 18898 18398
rect 19518 18450 19570 18462
rect 19518 18386 19570 18398
rect 20862 18450 20914 18462
rect 20862 18386 20914 18398
rect 21086 18450 21138 18462
rect 21086 18386 21138 18398
rect 23102 18450 23154 18462
rect 23102 18386 23154 18398
rect 24110 18450 24162 18462
rect 24110 18386 24162 18398
rect 26462 18450 26514 18462
rect 27358 18450 27410 18462
rect 28814 18450 28866 18462
rect 26786 18398 26798 18450
rect 26850 18398 26862 18450
rect 27122 18398 27134 18450
rect 27186 18398 27198 18450
rect 27906 18398 27918 18450
rect 27970 18398 27982 18450
rect 26462 18386 26514 18398
rect 27358 18386 27410 18398
rect 28814 18386 28866 18398
rect 29934 18450 29986 18462
rect 30942 18450 30994 18462
rect 30594 18398 30606 18450
rect 30658 18398 30670 18450
rect 29934 18386 29986 18398
rect 30942 18386 30994 18398
rect 37886 18450 37938 18462
rect 37886 18386 37938 18398
rect 15038 18338 15090 18350
rect 15038 18274 15090 18286
rect 17726 18338 17778 18350
rect 17726 18274 17778 18286
rect 21982 18338 22034 18350
rect 21982 18274 22034 18286
rect 22766 18338 22818 18350
rect 22766 18274 22818 18286
rect 28366 18338 28418 18350
rect 28366 18274 28418 18286
rect 31726 18338 31778 18350
rect 31726 18274 31778 18286
rect 11902 18226 11954 18238
rect 11902 18162 11954 18174
rect 12798 18226 12850 18238
rect 26002 18174 26014 18226
rect 26066 18174 26078 18226
rect 29474 18174 29486 18226
rect 29538 18174 29550 18226
rect 12798 18162 12850 18174
rect 1344 18058 38640 18092
rect 1344 18006 5876 18058
rect 5928 18006 5980 18058
rect 6032 18006 6084 18058
rect 6136 18006 15200 18058
rect 15252 18006 15304 18058
rect 15356 18006 15408 18058
rect 15460 18006 24524 18058
rect 24576 18006 24628 18058
rect 24680 18006 24732 18058
rect 24784 18006 33848 18058
rect 33900 18006 33952 18058
rect 34004 18006 34056 18058
rect 34108 18006 38640 18058
rect 1344 17972 38640 18006
rect 11902 17890 11954 17902
rect 11902 17826 11954 17838
rect 16830 17890 16882 17902
rect 23762 17838 23774 17890
rect 23826 17838 23838 17890
rect 16830 17826 16882 17838
rect 30606 17778 30658 17790
rect 21298 17726 21310 17778
rect 21362 17726 21374 17778
rect 30606 17714 30658 17726
rect 2718 17666 2770 17678
rect 2718 17602 2770 17614
rect 11678 17666 11730 17678
rect 14030 17666 14082 17678
rect 13794 17614 13806 17666
rect 13858 17614 13870 17666
rect 11678 17602 11730 17614
rect 14030 17602 14082 17614
rect 14142 17666 14194 17678
rect 16606 17666 16658 17678
rect 21758 17666 21810 17678
rect 23214 17666 23266 17678
rect 14578 17614 14590 17666
rect 14642 17614 14654 17666
rect 15138 17614 15150 17666
rect 15202 17614 15214 17666
rect 17154 17614 17166 17666
rect 17218 17614 17230 17666
rect 17714 17614 17726 17666
rect 17778 17614 17790 17666
rect 19954 17614 19966 17666
rect 20018 17614 20030 17666
rect 20514 17614 20526 17666
rect 20578 17614 20590 17666
rect 22082 17614 22094 17666
rect 22146 17614 22158 17666
rect 14142 17602 14194 17614
rect 16606 17602 16658 17614
rect 21758 17602 21810 17614
rect 23214 17602 23266 17614
rect 23326 17666 23378 17678
rect 23326 17602 23378 17614
rect 26462 17666 26514 17678
rect 26462 17602 26514 17614
rect 27358 17666 27410 17678
rect 27358 17602 27410 17614
rect 27470 17666 27522 17678
rect 27470 17602 27522 17614
rect 29598 17666 29650 17678
rect 29598 17602 29650 17614
rect 37886 17666 37938 17678
rect 37886 17602 37938 17614
rect 1710 17554 1762 17566
rect 1710 17490 1762 17502
rect 3166 17554 3218 17566
rect 3166 17490 3218 17502
rect 12910 17554 12962 17566
rect 12910 17490 12962 17502
rect 14926 17554 14978 17566
rect 14926 17490 14978 17502
rect 15598 17554 15650 17566
rect 15598 17490 15650 17502
rect 15934 17554 15986 17566
rect 15934 17490 15986 17502
rect 21870 17554 21922 17566
rect 21870 17490 21922 17502
rect 22654 17554 22706 17566
rect 22654 17490 22706 17502
rect 23102 17554 23154 17566
rect 23102 17490 23154 17502
rect 24334 17554 24386 17566
rect 24334 17490 24386 17502
rect 24670 17554 24722 17566
rect 24670 17490 24722 17502
rect 27246 17554 27298 17566
rect 28254 17554 28306 17566
rect 27906 17502 27918 17554
rect 27970 17502 27982 17554
rect 27246 17490 27298 17502
rect 28254 17490 28306 17502
rect 37214 17554 37266 17566
rect 37214 17490 37266 17502
rect 38222 17554 38274 17566
rect 38222 17490 38274 17502
rect 2046 17442 2098 17454
rect 2046 17378 2098 17390
rect 2382 17442 2434 17454
rect 2382 17378 2434 17390
rect 11342 17442 11394 17454
rect 12574 17442 12626 17454
rect 12226 17390 12238 17442
rect 12290 17390 12302 17442
rect 11342 17378 11394 17390
rect 12574 17378 12626 17390
rect 17502 17442 17554 17454
rect 17502 17378 17554 17390
rect 18286 17442 18338 17454
rect 18286 17378 18338 17390
rect 18958 17442 19010 17454
rect 18958 17378 19010 17390
rect 19406 17442 19458 17454
rect 19406 17378 19458 17390
rect 19742 17442 19794 17454
rect 19742 17378 19794 17390
rect 20750 17442 20802 17454
rect 20750 17378 20802 17390
rect 25006 17442 25058 17454
rect 25006 17378 25058 17390
rect 26798 17442 26850 17454
rect 26798 17378 26850 17390
rect 28590 17442 28642 17454
rect 28590 17378 28642 17390
rect 29262 17442 29314 17454
rect 29262 17378 29314 17390
rect 29934 17442 29986 17454
rect 29934 17378 29986 17390
rect 37550 17442 37602 17454
rect 37550 17378 37602 17390
rect 1344 17274 38800 17308
rect 1344 17222 10538 17274
rect 10590 17222 10642 17274
rect 10694 17222 10746 17274
rect 10798 17222 19862 17274
rect 19914 17222 19966 17274
rect 20018 17222 20070 17274
rect 20122 17222 29186 17274
rect 29238 17222 29290 17274
rect 29342 17222 29394 17274
rect 29446 17222 38510 17274
rect 38562 17222 38614 17274
rect 38666 17222 38718 17274
rect 38770 17222 38800 17274
rect 1344 17188 38800 17222
rect 13470 17106 13522 17118
rect 16494 17106 16546 17118
rect 24670 17106 24722 17118
rect 13682 17054 13694 17106
rect 13746 17054 13758 17106
rect 17938 17054 17950 17106
rect 18002 17054 18014 17106
rect 19618 17054 19630 17106
rect 19682 17054 19694 17106
rect 23986 17054 23998 17106
rect 24050 17054 24062 17106
rect 13470 17042 13522 17054
rect 16494 17042 16546 17054
rect 24670 17042 24722 17054
rect 26910 17106 26962 17118
rect 26910 17042 26962 17054
rect 1710 16994 1762 17006
rect 1710 16930 1762 16942
rect 12126 16994 12178 17006
rect 12126 16930 12178 16942
rect 12910 16994 12962 17006
rect 12910 16930 12962 16942
rect 14142 16994 14194 17006
rect 14142 16930 14194 16942
rect 14366 16994 14418 17006
rect 14366 16930 14418 16942
rect 18286 16994 18338 17006
rect 18286 16930 18338 16942
rect 18622 16994 18674 17006
rect 18622 16930 18674 16942
rect 18958 16994 19010 17006
rect 18958 16930 19010 16942
rect 20078 16994 20130 17006
rect 20078 16930 20130 16942
rect 21086 16994 21138 17006
rect 21086 16930 21138 16942
rect 21198 16994 21250 17006
rect 21198 16930 21250 16942
rect 22318 16994 22370 17006
rect 22318 16930 22370 16942
rect 23438 16994 23490 17006
rect 23438 16930 23490 16942
rect 23550 16994 23602 17006
rect 23550 16930 23602 16942
rect 25566 16994 25618 17006
rect 25566 16930 25618 16942
rect 28478 16994 28530 17006
rect 28478 16930 28530 16942
rect 28814 16994 28866 17006
rect 28814 16930 28866 16942
rect 29150 16994 29202 17006
rect 29150 16930 29202 16942
rect 31950 16994 32002 17006
rect 31950 16930 32002 16942
rect 37886 16994 37938 17006
rect 37886 16930 37938 16942
rect 38222 16994 38274 17006
rect 38222 16930 38274 16942
rect 2046 16882 2098 16894
rect 14254 16882 14306 16894
rect 17614 16882 17666 16894
rect 20190 16882 20242 16894
rect 20974 16882 21026 16894
rect 21982 16882 22034 16894
rect 12338 16830 12350 16882
rect 12402 16830 12414 16882
rect 15922 16830 15934 16882
rect 15986 16830 15998 16882
rect 16706 16830 16718 16882
rect 16770 16830 16782 16882
rect 19170 16830 19182 16882
rect 19234 16830 19246 16882
rect 20402 16830 20414 16882
rect 20466 16830 20478 16882
rect 21634 16830 21646 16882
rect 21698 16830 21710 16882
rect 2046 16818 2098 16830
rect 14254 16818 14306 16830
rect 17614 16818 17666 16830
rect 20190 16818 20242 16830
rect 20974 16818 21026 16830
rect 21982 16818 22034 16830
rect 22878 16882 22930 16894
rect 22878 16818 22930 16830
rect 23326 16882 23378 16894
rect 23326 16818 23378 16830
rect 24334 16882 24386 16894
rect 26462 16882 26514 16894
rect 28142 16882 28194 16894
rect 25330 16830 25342 16882
rect 25394 16830 25406 16882
rect 27794 16830 27806 16882
rect 27858 16830 27870 16882
rect 24334 16818 24386 16830
rect 26462 16818 26514 16830
rect 28142 16818 28194 16830
rect 29822 16882 29874 16894
rect 29822 16818 29874 16830
rect 30718 16882 30770 16894
rect 31614 16882 31666 16894
rect 31266 16830 31278 16882
rect 31330 16830 31342 16882
rect 30718 16818 30770 16830
rect 31614 16818 31666 16830
rect 32398 16882 32450 16894
rect 32398 16818 32450 16830
rect 15374 16770 15426 16782
rect 15374 16706 15426 16718
rect 26238 16770 26290 16782
rect 26238 16706 26290 16718
rect 27246 16770 27298 16782
rect 27246 16706 27298 16718
rect 27470 16770 27522 16782
rect 27470 16706 27522 16718
rect 15598 16658 15650 16670
rect 30046 16658 30098 16670
rect 30942 16658 30994 16670
rect 25890 16606 25902 16658
rect 25954 16606 25966 16658
rect 30370 16606 30382 16658
rect 30434 16606 30446 16658
rect 15598 16594 15650 16606
rect 30046 16594 30098 16606
rect 30942 16594 30994 16606
rect 1344 16490 38640 16524
rect 1344 16438 5876 16490
rect 5928 16438 5980 16490
rect 6032 16438 6084 16490
rect 6136 16438 15200 16490
rect 15252 16438 15304 16490
rect 15356 16438 15408 16490
rect 15460 16438 24524 16490
rect 24576 16438 24628 16490
rect 24680 16438 24732 16490
rect 24784 16438 33848 16490
rect 33900 16438 33952 16490
rect 34004 16438 34056 16490
rect 34108 16438 38640 16490
rect 1344 16404 38640 16438
rect 19518 16322 19570 16334
rect 19170 16270 19182 16322
rect 19234 16270 19246 16322
rect 19518 16258 19570 16270
rect 21534 16322 21586 16334
rect 23874 16270 23886 16322
rect 23938 16270 23950 16322
rect 28242 16270 28254 16322
rect 28306 16319 28318 16322
rect 28466 16319 28478 16322
rect 28306 16273 28478 16319
rect 28306 16270 28318 16273
rect 28466 16270 28478 16273
rect 28530 16270 28542 16322
rect 21534 16258 21586 16270
rect 21310 16210 21362 16222
rect 21310 16146 21362 16158
rect 24222 16210 24274 16222
rect 24222 16146 24274 16158
rect 25902 16210 25954 16222
rect 25902 16146 25954 16158
rect 19742 16098 19794 16110
rect 1922 16046 1934 16098
rect 1986 16046 1998 16098
rect 18386 16046 18398 16098
rect 18450 16046 18462 16098
rect 19742 16034 19794 16046
rect 22430 16098 22482 16110
rect 23326 16098 23378 16110
rect 23090 16046 23102 16098
rect 23154 16046 23166 16098
rect 22430 16034 22482 16046
rect 23326 16034 23378 16046
rect 23438 16098 23490 16110
rect 23438 16034 23490 16046
rect 24446 16098 24498 16110
rect 24446 16034 24498 16046
rect 26238 16098 26290 16110
rect 26238 16034 26290 16046
rect 30494 16098 30546 16110
rect 30494 16034 30546 16046
rect 37886 16098 37938 16110
rect 37886 16034 37938 16046
rect 22766 15986 22818 15998
rect 25118 15986 25170 15998
rect 16706 15934 16718 15986
rect 16770 15934 16782 15986
rect 24770 15934 24782 15986
rect 24834 15934 24846 15986
rect 22766 15922 22818 15934
rect 25118 15922 25170 15934
rect 26574 15986 26626 15998
rect 26574 15922 26626 15934
rect 27694 15986 27746 15998
rect 27694 15922 27746 15934
rect 1710 15874 1762 15886
rect 20414 15874 20466 15886
rect 25454 15874 25506 15886
rect 20066 15822 20078 15874
rect 20130 15822 20142 15874
rect 21858 15822 21870 15874
rect 21922 15822 21934 15874
rect 1710 15810 1762 15822
rect 20414 15810 20466 15822
rect 25454 15810 25506 15822
rect 28030 15874 28082 15886
rect 28030 15810 28082 15822
rect 28478 15874 28530 15886
rect 28478 15810 28530 15822
rect 30830 15874 30882 15886
rect 30830 15810 30882 15822
rect 38222 15874 38274 15886
rect 38222 15810 38274 15822
rect 1344 15706 38800 15740
rect 1344 15654 10538 15706
rect 10590 15654 10642 15706
rect 10694 15654 10746 15706
rect 10798 15654 19862 15706
rect 19914 15654 19966 15706
rect 20018 15654 20070 15706
rect 20122 15654 29186 15706
rect 29238 15654 29290 15706
rect 29342 15654 29394 15706
rect 29446 15654 38510 15706
rect 38562 15654 38614 15706
rect 38666 15654 38718 15706
rect 38770 15654 38800 15706
rect 1344 15620 38800 15654
rect 27682 15486 27694 15538
rect 27746 15486 27758 15538
rect 1710 15426 1762 15438
rect 24110 15426 24162 15438
rect 20178 15374 20190 15426
rect 20242 15374 20254 15426
rect 1710 15362 1762 15374
rect 24110 15362 24162 15374
rect 25566 15426 25618 15438
rect 25566 15362 25618 15374
rect 31054 15426 31106 15438
rect 31054 15362 31106 15374
rect 38222 15426 38274 15438
rect 38222 15362 38274 15374
rect 2046 15314 2098 15326
rect 23214 15314 23266 15326
rect 25230 15314 25282 15326
rect 14018 15262 14030 15314
rect 14082 15262 14094 15314
rect 17378 15262 17390 15314
rect 17442 15262 17454 15314
rect 23762 15262 23774 15314
rect 23826 15262 23838 15314
rect 24322 15262 24334 15314
rect 24386 15262 24398 15314
rect 2046 15250 2098 15262
rect 23214 15250 23266 15262
rect 25230 15250 25282 15262
rect 27134 15314 27186 15326
rect 27134 15250 27186 15262
rect 28030 15314 28082 15326
rect 28030 15250 28082 15262
rect 28254 15314 28306 15326
rect 28254 15250 28306 15262
rect 29150 15314 29202 15326
rect 29150 15250 29202 15262
rect 29822 15314 29874 15326
rect 29822 15250 29874 15262
rect 30046 15314 30098 15326
rect 30718 15314 30770 15326
rect 30370 15262 30382 15314
rect 30434 15262 30446 15314
rect 30046 15250 30098 15262
rect 30718 15250 30770 15262
rect 31502 15314 31554 15326
rect 31502 15250 31554 15262
rect 37886 15314 37938 15326
rect 37886 15250 37938 15262
rect 23438 15202 23490 15214
rect 14690 15150 14702 15202
rect 14754 15150 14766 15202
rect 16818 15150 16830 15202
rect 16882 15150 16894 15202
rect 23438 15138 23490 15150
rect 27358 15202 27410 15214
rect 27358 15138 27410 15150
rect 28926 15202 28978 15214
rect 28926 15138 28978 15150
rect 26786 15038 26798 15090
rect 26850 15038 26862 15090
rect 29474 15038 29486 15090
rect 29538 15038 29550 15090
rect 1344 14922 38640 14956
rect 1344 14870 5876 14922
rect 5928 14870 5980 14922
rect 6032 14870 6084 14922
rect 6136 14870 15200 14922
rect 15252 14870 15304 14922
rect 15356 14870 15408 14922
rect 15460 14870 24524 14922
rect 24576 14870 24628 14922
rect 24680 14870 24732 14922
rect 24784 14870 33848 14922
rect 33900 14870 33952 14922
rect 34004 14870 34056 14922
rect 34108 14870 38640 14922
rect 1344 14836 38640 14870
rect 18286 14754 18338 14766
rect 18286 14690 18338 14702
rect 18510 14754 18562 14766
rect 18510 14690 18562 14702
rect 18958 14754 19010 14766
rect 18958 14690 19010 14702
rect 20414 14754 20466 14766
rect 20414 14690 20466 14702
rect 28478 14642 28530 14654
rect 17042 14590 17054 14642
rect 17106 14590 17118 14642
rect 28478 14578 28530 14590
rect 18062 14530 18114 14542
rect 19742 14530 19794 14542
rect 14242 14478 14254 14530
rect 14306 14478 14318 14530
rect 19394 14478 19406 14530
rect 19458 14478 19470 14530
rect 18062 14466 18114 14478
rect 19742 14466 19794 14478
rect 20190 14530 20242 14542
rect 27134 14530 27186 14542
rect 21858 14478 21870 14530
rect 21922 14478 21934 14530
rect 20190 14466 20242 14478
rect 27134 14466 27186 14478
rect 29486 14530 29538 14542
rect 29486 14466 29538 14478
rect 1710 14418 1762 14430
rect 17614 14418 17666 14430
rect 14914 14366 14926 14418
rect 14978 14366 14990 14418
rect 1710 14354 1762 14366
rect 17614 14354 17666 14366
rect 19182 14418 19234 14430
rect 27470 14418 27522 14430
rect 23538 14366 23550 14418
rect 23602 14366 23614 14418
rect 19182 14354 19234 14366
rect 27470 14354 27522 14366
rect 37886 14418 37938 14430
rect 37886 14354 37938 14366
rect 2046 14306 2098 14318
rect 2046 14242 2098 14254
rect 2494 14306 2546 14318
rect 2494 14242 2546 14254
rect 17726 14306 17778 14318
rect 17726 14242 17778 14254
rect 19070 14306 19122 14318
rect 29822 14306 29874 14318
rect 20738 14254 20750 14306
rect 20802 14254 20814 14306
rect 19070 14242 19122 14254
rect 29822 14242 29874 14254
rect 38222 14306 38274 14318
rect 38222 14242 38274 14254
rect 1344 14138 38800 14172
rect 1344 14086 10538 14138
rect 10590 14086 10642 14138
rect 10694 14086 10746 14138
rect 10798 14086 19862 14138
rect 19914 14086 19966 14138
rect 20018 14086 20070 14138
rect 20122 14086 29186 14138
rect 29238 14086 29290 14138
rect 29342 14086 29394 14138
rect 29446 14086 38510 14138
rect 38562 14086 38614 14138
rect 38666 14086 38718 14138
rect 38770 14086 38800 14138
rect 1344 14052 38800 14086
rect 2046 13970 2098 13982
rect 2046 13906 2098 13918
rect 15822 13970 15874 13982
rect 15822 13906 15874 13918
rect 19854 13970 19906 13982
rect 19854 13906 19906 13918
rect 15486 13858 15538 13870
rect 19966 13858 20018 13870
rect 19506 13806 19518 13858
rect 19570 13806 19582 13858
rect 15486 13794 15538 13806
rect 19966 13794 20018 13806
rect 20974 13858 21026 13870
rect 20974 13794 21026 13806
rect 25566 13858 25618 13870
rect 25566 13794 25618 13806
rect 38222 13858 38274 13870
rect 38222 13794 38274 13806
rect 1710 13746 1762 13758
rect 1710 13682 1762 13694
rect 18062 13746 18114 13758
rect 18062 13682 18114 13694
rect 18510 13746 18562 13758
rect 18510 13682 18562 13694
rect 18958 13746 19010 13758
rect 18958 13682 19010 13694
rect 19182 13746 19234 13758
rect 21646 13746 21698 13758
rect 20738 13694 20750 13746
rect 20802 13694 20814 13746
rect 19182 13682 19234 13694
rect 21646 13682 21698 13694
rect 22990 13746 23042 13758
rect 22990 13682 23042 13694
rect 23886 13746 23938 13758
rect 25230 13746 25282 13758
rect 24210 13694 24222 13746
rect 24274 13694 24286 13746
rect 23886 13682 23938 13694
rect 25230 13682 25282 13694
rect 37886 13746 37938 13758
rect 37886 13682 37938 13694
rect 2494 13634 2546 13646
rect 2494 13570 2546 13582
rect 16830 13634 16882 13646
rect 16830 13570 16882 13582
rect 17614 13634 17666 13646
rect 21870 13634 21922 13646
rect 21298 13582 21310 13634
rect 21362 13582 21374 13634
rect 17614 13570 17666 13582
rect 21870 13570 21922 13582
rect 22318 13634 22370 13646
rect 22318 13570 22370 13582
rect 22766 13634 22818 13646
rect 22766 13570 22818 13582
rect 23662 13634 23714 13646
rect 23662 13570 23714 13582
rect 24670 13634 24722 13646
rect 24670 13570 24722 13582
rect 17726 13522 17778 13534
rect 17726 13458 17778 13470
rect 18286 13522 18338 13534
rect 23314 13470 23326 13522
rect 23378 13470 23390 13522
rect 18286 13458 18338 13470
rect 1344 13354 38640 13388
rect 1344 13302 5876 13354
rect 5928 13302 5980 13354
rect 6032 13302 6084 13354
rect 6136 13302 15200 13354
rect 15252 13302 15304 13354
rect 15356 13302 15408 13354
rect 15460 13302 24524 13354
rect 24576 13302 24628 13354
rect 24680 13302 24732 13354
rect 24784 13302 33848 13354
rect 33900 13302 33952 13354
rect 34004 13302 34056 13354
rect 34108 13302 38640 13354
rect 1344 13268 38640 13302
rect 37214 12962 37266 12974
rect 17714 12910 17726 12962
rect 17778 12910 17790 12962
rect 17938 12910 17950 12962
rect 18002 12910 18014 12962
rect 21970 12910 21982 12962
rect 22034 12910 22046 12962
rect 23314 12910 23326 12962
rect 23378 12910 23390 12962
rect 37214 12898 37266 12910
rect 1710 12850 1762 12862
rect 1710 12786 1762 12798
rect 2046 12850 2098 12862
rect 2046 12786 2098 12798
rect 2494 12850 2546 12862
rect 2494 12786 2546 12798
rect 37886 12850 37938 12862
rect 37886 12786 37938 12798
rect 38222 12850 38274 12862
rect 38222 12786 38274 12798
rect 17390 12738 17442 12750
rect 17390 12674 17442 12686
rect 17502 12738 17554 12750
rect 17502 12674 17554 12686
rect 21422 12738 21474 12750
rect 21422 12674 21474 12686
rect 21758 12738 21810 12750
rect 21758 12674 21810 12686
rect 23550 12738 23602 12750
rect 23550 12674 23602 12686
rect 24446 12738 24498 12750
rect 24446 12674 24498 12686
rect 37550 12738 37602 12750
rect 37550 12674 37602 12686
rect 1344 12570 38800 12604
rect 1344 12518 10538 12570
rect 10590 12518 10642 12570
rect 10694 12518 10746 12570
rect 10798 12518 19862 12570
rect 19914 12518 19966 12570
rect 20018 12518 20070 12570
rect 20122 12518 29186 12570
rect 29238 12518 29290 12570
rect 29342 12518 29394 12570
rect 29446 12518 38510 12570
rect 38562 12518 38614 12570
rect 38666 12518 38718 12570
rect 38770 12518 38800 12570
rect 1344 12484 38800 12518
rect 37886 12402 37938 12414
rect 37886 12338 37938 12350
rect 37662 12178 37714 12190
rect 37662 12114 37714 12126
rect 38222 12178 38274 12190
rect 38222 12114 38274 12126
rect 1344 11786 38640 11820
rect 1344 11734 5876 11786
rect 5928 11734 5980 11786
rect 6032 11734 6084 11786
rect 6136 11734 15200 11786
rect 15252 11734 15304 11786
rect 15356 11734 15408 11786
rect 15460 11734 24524 11786
rect 24576 11734 24628 11786
rect 24680 11734 24732 11786
rect 24784 11734 33848 11786
rect 33900 11734 33952 11786
rect 34004 11734 34056 11786
rect 34108 11734 38640 11786
rect 1344 11700 38640 11734
rect 37886 11282 37938 11294
rect 37886 11218 37938 11230
rect 38222 11170 38274 11182
rect 38222 11106 38274 11118
rect 1344 11002 38800 11036
rect 1344 10950 10538 11002
rect 10590 10950 10642 11002
rect 10694 10950 10746 11002
rect 10798 10950 19862 11002
rect 19914 10950 19966 11002
rect 20018 10950 20070 11002
rect 20122 10950 29186 11002
rect 29238 10950 29290 11002
rect 29342 10950 29394 11002
rect 29446 10950 38510 11002
rect 38562 10950 38614 11002
rect 38666 10950 38718 11002
rect 38770 10950 38800 11002
rect 1344 10916 38800 10950
rect 38222 10722 38274 10734
rect 38222 10658 38274 10670
rect 37886 10610 37938 10622
rect 37886 10546 37938 10558
rect 1344 10218 38640 10252
rect 1344 10166 5876 10218
rect 5928 10166 5980 10218
rect 6032 10166 6084 10218
rect 6136 10166 15200 10218
rect 15252 10166 15304 10218
rect 15356 10166 15408 10218
rect 15460 10166 24524 10218
rect 24576 10166 24628 10218
rect 24680 10166 24732 10218
rect 24784 10166 33848 10218
rect 33900 10166 33952 10218
rect 34004 10166 34056 10218
rect 34108 10166 38640 10218
rect 1344 10132 38640 10166
rect 37886 9714 37938 9726
rect 37886 9650 37938 9662
rect 38222 9714 38274 9726
rect 38222 9650 38274 9662
rect 37662 9602 37714 9614
rect 37662 9538 37714 9550
rect 1344 9434 38800 9468
rect 1344 9382 10538 9434
rect 10590 9382 10642 9434
rect 10694 9382 10746 9434
rect 10798 9382 19862 9434
rect 19914 9382 19966 9434
rect 20018 9382 20070 9434
rect 20122 9382 29186 9434
rect 29238 9382 29290 9434
rect 29342 9382 29394 9434
rect 29446 9382 38510 9434
rect 38562 9382 38614 9434
rect 38666 9382 38718 9434
rect 38770 9382 38800 9434
rect 1344 9348 38800 9382
rect 37886 9154 37938 9166
rect 37886 9090 37938 9102
rect 38222 9154 38274 9166
rect 38222 9090 38274 9102
rect 1344 8650 38640 8684
rect 1344 8598 5876 8650
rect 5928 8598 5980 8650
rect 6032 8598 6084 8650
rect 6136 8598 15200 8650
rect 15252 8598 15304 8650
rect 15356 8598 15408 8650
rect 15460 8598 24524 8650
rect 24576 8598 24628 8650
rect 24680 8598 24732 8650
rect 24784 8598 33848 8650
rect 33900 8598 33952 8650
rect 34004 8598 34056 8650
rect 34108 8598 38640 8650
rect 1344 8564 38640 8598
rect 37214 8146 37266 8158
rect 38222 8146 38274 8158
rect 37874 8094 37886 8146
rect 37938 8094 37950 8146
rect 37214 8082 37266 8094
rect 38222 8082 38274 8094
rect 36430 8034 36482 8046
rect 36430 7970 36482 7982
rect 37550 8034 37602 8046
rect 37550 7970 37602 7982
rect 1344 7866 38800 7900
rect 1344 7814 10538 7866
rect 10590 7814 10642 7866
rect 10694 7814 10746 7866
rect 10798 7814 19862 7866
rect 19914 7814 19966 7866
rect 20018 7814 20070 7866
rect 20122 7814 29186 7866
rect 29238 7814 29290 7866
rect 29342 7814 29394 7866
rect 29446 7814 38510 7866
rect 38562 7814 38614 7866
rect 38666 7814 38718 7866
rect 38770 7814 38800 7866
rect 1344 7780 38800 7814
rect 37662 7698 37714 7710
rect 37662 7634 37714 7646
rect 38222 7586 38274 7598
rect 38222 7522 38274 7534
rect 37886 7474 37938 7486
rect 37886 7410 37938 7422
rect 37214 7362 37266 7374
rect 37214 7298 37266 7310
rect 1344 7082 38640 7116
rect 1344 7030 5876 7082
rect 5928 7030 5980 7082
rect 6032 7030 6084 7082
rect 6136 7030 15200 7082
rect 15252 7030 15304 7082
rect 15356 7030 15408 7082
rect 15460 7030 24524 7082
rect 24576 7030 24628 7082
rect 24680 7030 24732 7082
rect 24784 7030 33848 7082
rect 33900 7030 33952 7082
rect 34004 7030 34056 7082
rect 34108 7030 38640 7082
rect 1344 6996 38640 7030
rect 37550 6578 37602 6590
rect 37550 6514 37602 6526
rect 37886 6578 37938 6590
rect 37886 6514 37938 6526
rect 38222 6466 38274 6478
rect 38222 6402 38274 6414
rect 1344 6298 38800 6332
rect 1344 6246 10538 6298
rect 10590 6246 10642 6298
rect 10694 6246 10746 6298
rect 10798 6246 19862 6298
rect 19914 6246 19966 6298
rect 20018 6246 20070 6298
rect 20122 6246 29186 6298
rect 29238 6246 29290 6298
rect 29342 6246 29394 6298
rect 29446 6246 38510 6298
rect 38562 6246 38614 6298
rect 38666 6246 38718 6298
rect 38770 6246 38800 6298
rect 1344 6212 38800 6246
rect 38222 6018 38274 6030
rect 38222 5954 38274 5966
rect 37886 5906 37938 5918
rect 37886 5842 37938 5854
rect 37662 5794 37714 5806
rect 37662 5730 37714 5742
rect 1344 5514 38640 5548
rect 1344 5462 5876 5514
rect 5928 5462 5980 5514
rect 6032 5462 6084 5514
rect 6136 5462 15200 5514
rect 15252 5462 15304 5514
rect 15356 5462 15408 5514
rect 15460 5462 24524 5514
rect 24576 5462 24628 5514
rect 24680 5462 24732 5514
rect 24784 5462 33848 5514
rect 33900 5462 33952 5514
rect 34004 5462 34056 5514
rect 34108 5462 38640 5514
rect 1344 5428 38640 5462
rect 37550 5122 37602 5134
rect 37986 5070 37998 5122
rect 38050 5070 38062 5122
rect 37550 5058 37602 5070
rect 38222 4898 38274 4910
rect 38222 4834 38274 4846
rect 1344 4730 38800 4764
rect 1344 4678 10538 4730
rect 10590 4678 10642 4730
rect 10694 4678 10746 4730
rect 10798 4678 19862 4730
rect 19914 4678 19966 4730
rect 20018 4678 20070 4730
rect 20122 4678 29186 4730
rect 29238 4678 29290 4730
rect 29342 4678 29394 4730
rect 29446 4678 38510 4730
rect 38562 4678 38614 4730
rect 38666 4678 38718 4730
rect 38770 4678 38800 4730
rect 1344 4644 38800 4678
rect 38222 4450 38274 4462
rect 16370 4398 16382 4450
rect 16434 4398 16446 4450
rect 38222 4386 38274 4398
rect 37886 4338 37938 4350
rect 16594 4286 16606 4338
rect 16658 4286 16670 4338
rect 37886 4274 37938 4286
rect 15934 4226 15986 4238
rect 15934 4162 15986 4174
rect 25678 4226 25730 4238
rect 25678 4162 25730 4174
rect 26350 4226 26402 4238
rect 26350 4162 26402 4174
rect 37662 4226 37714 4238
rect 37662 4162 37714 4174
rect 1344 3946 38640 3980
rect 1344 3894 5876 3946
rect 5928 3894 5980 3946
rect 6032 3894 6084 3946
rect 6136 3894 15200 3946
rect 15252 3894 15304 3946
rect 15356 3894 15408 3946
rect 15460 3894 24524 3946
rect 24576 3894 24628 3946
rect 24680 3894 24732 3946
rect 24784 3894 33848 3946
rect 33900 3894 33952 3946
rect 34004 3894 34056 3946
rect 34108 3894 38640 3946
rect 1344 3860 38640 3894
rect 16046 3554 16098 3566
rect 19854 3554 19906 3566
rect 15474 3502 15486 3554
rect 15538 3502 15550 3554
rect 17266 3502 17278 3554
rect 17330 3502 17342 3554
rect 17938 3502 17950 3554
rect 18002 3502 18014 3554
rect 18610 3502 18622 3554
rect 18674 3502 18686 3554
rect 19282 3502 19294 3554
rect 19346 3502 19358 3554
rect 16046 3490 16098 3502
rect 19854 3490 19906 3502
rect 21422 3554 21474 3566
rect 22766 3554 22818 3566
rect 25566 3554 25618 3566
rect 21970 3502 21982 3554
rect 22034 3502 22046 3554
rect 23314 3502 23326 3554
rect 23378 3502 23390 3554
rect 24770 3502 24782 3554
rect 24834 3502 24846 3554
rect 21422 3490 21474 3502
rect 22766 3490 22818 3502
rect 25566 3490 25618 3502
rect 26238 3554 26290 3566
rect 26786 3502 26798 3554
rect 26850 3502 26862 3554
rect 27458 3502 27470 3554
rect 27522 3502 27534 3554
rect 26238 3490 26290 3502
rect 24110 3442 24162 3454
rect 15698 3390 15710 3442
rect 15762 3390 15774 3442
rect 16370 3390 16382 3442
rect 16434 3390 16446 3442
rect 24110 3378 24162 3390
rect 24558 3442 24610 3454
rect 24558 3378 24610 3390
rect 25230 3442 25282 3454
rect 25230 3378 25282 3390
rect 25902 3442 25954 3454
rect 25902 3378 25954 3390
rect 26574 3442 26626 3454
rect 26574 3378 26626 3390
rect 27246 3442 27298 3454
rect 27246 3378 27298 3390
rect 36430 3442 36482 3454
rect 36430 3378 36482 3390
rect 36990 3442 37042 3454
rect 37550 3442 37602 3454
rect 37202 3390 37214 3442
rect 37266 3390 37278 3442
rect 36990 3378 37042 3390
rect 37550 3378 37602 3390
rect 37886 3442 37938 3454
rect 37886 3378 37938 3390
rect 38222 3442 38274 3454
rect 38222 3378 38274 3390
rect 17502 3330 17554 3342
rect 17502 3266 17554 3278
rect 18174 3330 18226 3342
rect 20190 3330 20242 3342
rect 18834 3278 18846 3330
rect 18898 3278 18910 3330
rect 19506 3278 19518 3330
rect 19570 3278 19582 3330
rect 18174 3266 18226 3278
rect 20190 3266 20242 3278
rect 21086 3330 21138 3342
rect 21086 3266 21138 3278
rect 21758 3330 21810 3342
rect 21758 3266 21810 3278
rect 22430 3330 22482 3342
rect 22430 3266 22482 3278
rect 23102 3330 23154 3342
rect 23102 3266 23154 3278
rect 1344 3162 38800 3196
rect 1344 3110 10538 3162
rect 10590 3110 10642 3162
rect 10694 3110 10746 3162
rect 10798 3110 19862 3162
rect 19914 3110 19966 3162
rect 20018 3110 20070 3162
rect 20122 3110 29186 3162
rect 29238 3110 29290 3162
rect 29342 3110 29394 3162
rect 29446 3110 38510 3162
rect 38562 3110 38614 3162
rect 38666 3110 38718 3162
rect 38770 3110 38800 3162
rect 1344 3076 38800 3110
rect 25554 2494 25566 2546
rect 25618 2543 25630 2546
rect 26338 2543 26350 2546
rect 25618 2497 26350 2543
rect 25618 2494 25630 2497
rect 26338 2494 26350 2497
rect 26402 2543 26414 2546
rect 26786 2543 26798 2546
rect 26402 2497 26798 2543
rect 26402 2494 26414 2497
rect 26786 2494 26798 2497
rect 26850 2494 26862 2546
<< via1 >>
rect 5876 36822 5928 36874
rect 5980 36822 6032 36874
rect 6084 36822 6136 36874
rect 15200 36822 15252 36874
rect 15304 36822 15356 36874
rect 15408 36822 15460 36874
rect 24524 36822 24576 36874
rect 24628 36822 24680 36874
rect 24732 36822 24784 36874
rect 33848 36822 33900 36874
rect 33952 36822 34004 36874
rect 34056 36822 34108 36874
rect 14814 36430 14866 36482
rect 17278 36430 17330 36482
rect 21310 36430 21362 36482
rect 21758 36430 21810 36482
rect 24782 36430 24834 36482
rect 26126 36430 26178 36482
rect 35534 36430 35586 36482
rect 37550 36430 37602 36482
rect 15374 36318 15426 36370
rect 15710 36318 15762 36370
rect 16046 36318 16098 36370
rect 16382 36318 16434 36370
rect 17502 36318 17554 36370
rect 17838 36318 17890 36370
rect 18174 36318 18226 36370
rect 18510 36318 18562 36370
rect 18846 36318 18898 36370
rect 19182 36318 19234 36370
rect 19518 36318 19570 36370
rect 19854 36318 19906 36370
rect 20190 36318 20242 36370
rect 21086 36318 21138 36370
rect 22430 36318 22482 36370
rect 22766 36318 22818 36370
rect 23102 36318 23154 36370
rect 23438 36318 23490 36370
rect 24558 36318 24610 36370
rect 25230 36318 25282 36370
rect 25566 36318 25618 36370
rect 36542 36318 36594 36370
rect 36878 36318 36930 36370
rect 15038 36206 15090 36258
rect 22094 36206 22146 36258
rect 25902 36206 25954 36258
rect 36318 36206 36370 36258
rect 37214 36206 37266 36258
rect 37886 36206 37938 36258
rect 38222 36206 38274 36258
rect 10538 36038 10590 36090
rect 10642 36038 10694 36090
rect 10746 36038 10798 36090
rect 19862 36038 19914 36090
rect 19966 36038 20018 36090
rect 20070 36038 20122 36090
rect 29186 36038 29238 36090
rect 29290 36038 29342 36090
rect 29394 36038 29446 36090
rect 38510 36038 38562 36090
rect 38614 36038 38666 36090
rect 38718 36038 38770 36090
rect 15262 35870 15314 35922
rect 16158 35870 16210 35922
rect 16382 35870 16434 35922
rect 21534 35870 21586 35922
rect 25678 35870 25730 35922
rect 37662 35870 37714 35922
rect 16718 35758 16770 35810
rect 38222 35758 38274 35810
rect 37102 35646 37154 35698
rect 37998 35646 38050 35698
rect 5876 35254 5928 35306
rect 5980 35254 6032 35306
rect 6084 35254 6136 35306
rect 15200 35254 15252 35306
rect 15304 35254 15356 35306
rect 15408 35254 15460 35306
rect 24524 35254 24576 35306
rect 24628 35254 24680 35306
rect 24732 35254 24784 35306
rect 33848 35254 33900 35306
rect 33952 35254 34004 35306
rect 34056 35254 34108 35306
rect 37886 34750 37938 34802
rect 38222 34638 38274 34690
rect 10538 34470 10590 34522
rect 10642 34470 10694 34522
rect 10746 34470 10798 34522
rect 19862 34470 19914 34522
rect 19966 34470 20018 34522
rect 20070 34470 20122 34522
rect 29186 34470 29238 34522
rect 29290 34470 29342 34522
rect 29394 34470 29446 34522
rect 38510 34470 38562 34522
rect 38614 34470 38666 34522
rect 38718 34470 38770 34522
rect 38222 34190 38274 34242
rect 37998 34078 38050 34130
rect 37550 33966 37602 34018
rect 5876 33686 5928 33738
rect 5980 33686 6032 33738
rect 6084 33686 6136 33738
rect 15200 33686 15252 33738
rect 15304 33686 15356 33738
rect 15408 33686 15460 33738
rect 24524 33686 24576 33738
rect 24628 33686 24680 33738
rect 24732 33686 24784 33738
rect 33848 33686 33900 33738
rect 33952 33686 34004 33738
rect 34056 33686 34108 33738
rect 37886 33182 37938 33234
rect 38222 33070 38274 33122
rect 10538 32902 10590 32954
rect 10642 32902 10694 32954
rect 10746 32902 10798 32954
rect 19862 32902 19914 32954
rect 19966 32902 20018 32954
rect 20070 32902 20122 32954
rect 29186 32902 29238 32954
rect 29290 32902 29342 32954
rect 29394 32902 29446 32954
rect 38510 32902 38562 32954
rect 38614 32902 38666 32954
rect 38718 32902 38770 32954
rect 37886 32622 37938 32674
rect 38222 32510 38274 32562
rect 37214 32398 37266 32450
rect 37662 32398 37714 32450
rect 5876 32118 5928 32170
rect 5980 32118 6032 32170
rect 6084 32118 6136 32170
rect 15200 32118 15252 32170
rect 15304 32118 15356 32170
rect 15408 32118 15460 32170
rect 24524 32118 24576 32170
rect 24628 32118 24680 32170
rect 24732 32118 24784 32170
rect 33848 32118 33900 32170
rect 33952 32118 34004 32170
rect 34056 32118 34108 32170
rect 37886 31726 37938 31778
rect 37214 31614 37266 31666
rect 37550 31614 37602 31666
rect 36542 31502 36594 31554
rect 38222 31502 38274 31554
rect 10538 31334 10590 31386
rect 10642 31334 10694 31386
rect 10746 31334 10798 31386
rect 19862 31334 19914 31386
rect 19966 31334 20018 31386
rect 20070 31334 20122 31386
rect 29186 31334 29238 31386
rect 29290 31334 29342 31386
rect 29394 31334 29446 31386
rect 38510 31334 38562 31386
rect 38614 31334 38666 31386
rect 38718 31334 38770 31386
rect 38222 31054 38274 31106
rect 37886 30942 37938 30994
rect 37550 30830 37602 30882
rect 5876 30550 5928 30602
rect 5980 30550 6032 30602
rect 6084 30550 6136 30602
rect 15200 30550 15252 30602
rect 15304 30550 15356 30602
rect 15408 30550 15460 30602
rect 24524 30550 24576 30602
rect 24628 30550 24680 30602
rect 24732 30550 24784 30602
rect 33848 30550 33900 30602
rect 33952 30550 34004 30602
rect 34056 30550 34108 30602
rect 37886 30046 37938 30098
rect 37662 29934 37714 29986
rect 38222 29934 38274 29986
rect 10538 29766 10590 29818
rect 10642 29766 10694 29818
rect 10746 29766 10798 29818
rect 19862 29766 19914 29818
rect 19966 29766 20018 29818
rect 20070 29766 20122 29818
rect 29186 29766 29238 29818
rect 29290 29766 29342 29818
rect 29394 29766 29446 29818
rect 38510 29766 38562 29818
rect 38614 29766 38666 29818
rect 38718 29766 38770 29818
rect 38222 29486 38274 29538
rect 37886 29374 37938 29426
rect 5876 28982 5928 29034
rect 5980 28982 6032 29034
rect 6084 28982 6136 29034
rect 15200 28982 15252 29034
rect 15304 28982 15356 29034
rect 15408 28982 15460 29034
rect 24524 28982 24576 29034
rect 24628 28982 24680 29034
rect 24732 28982 24784 29034
rect 33848 28982 33900 29034
rect 33952 28982 34004 29034
rect 34056 28982 34108 29034
rect 37886 28590 37938 28642
rect 37662 28366 37714 28418
rect 38222 28366 38274 28418
rect 10538 28198 10590 28250
rect 10642 28198 10694 28250
rect 10746 28198 10798 28250
rect 19862 28198 19914 28250
rect 19966 28198 20018 28250
rect 20070 28198 20122 28250
rect 29186 28198 29238 28250
rect 29290 28198 29342 28250
rect 29394 28198 29446 28250
rect 38510 28198 38562 28250
rect 38614 28198 38666 28250
rect 38718 28198 38770 28250
rect 38222 27918 38274 27970
rect 37886 27806 37938 27858
rect 5876 27414 5928 27466
rect 5980 27414 6032 27466
rect 6084 27414 6136 27466
rect 15200 27414 15252 27466
rect 15304 27414 15356 27466
rect 15408 27414 15460 27466
rect 24524 27414 24576 27466
rect 24628 27414 24680 27466
rect 24732 27414 24784 27466
rect 33848 27414 33900 27466
rect 33952 27414 34004 27466
rect 34056 27414 34108 27466
rect 1822 27022 1874 27074
rect 37214 27022 37266 27074
rect 37998 27022 38050 27074
rect 2494 26910 2546 26962
rect 37550 26910 37602 26962
rect 38222 26910 38274 26962
rect 2046 26798 2098 26850
rect 10538 26630 10590 26682
rect 10642 26630 10694 26682
rect 10746 26630 10798 26682
rect 19862 26630 19914 26682
rect 19966 26630 20018 26682
rect 20070 26630 20122 26682
rect 29186 26630 29238 26682
rect 29290 26630 29342 26682
rect 29394 26630 29446 26682
rect 38510 26630 38562 26682
rect 38614 26630 38666 26682
rect 38718 26630 38770 26682
rect 22318 26462 22370 26514
rect 1710 26350 1762 26402
rect 37886 26350 37938 26402
rect 2046 26238 2098 26290
rect 38222 26238 38274 26290
rect 2494 26126 2546 26178
rect 37662 26126 37714 26178
rect 2270 26014 2322 26066
rect 2494 26014 2546 26066
rect 5876 25846 5928 25898
rect 5980 25846 6032 25898
rect 6084 25846 6136 25898
rect 15200 25846 15252 25898
rect 15304 25846 15356 25898
rect 15408 25846 15460 25898
rect 24524 25846 24576 25898
rect 24628 25846 24680 25898
rect 24732 25846 24784 25898
rect 33848 25846 33900 25898
rect 33952 25846 34004 25898
rect 34056 25846 34108 25898
rect 1822 25454 1874 25506
rect 19854 25454 19906 25506
rect 21422 25454 21474 25506
rect 22094 25454 22146 25506
rect 23102 25454 23154 25506
rect 25790 25454 25842 25506
rect 26462 25454 26514 25506
rect 28366 25454 28418 25506
rect 17726 25342 17778 25394
rect 18062 25342 18114 25394
rect 19630 25342 19682 25394
rect 21534 25342 21586 25394
rect 21646 25342 21698 25394
rect 22430 25342 22482 25394
rect 22766 25342 22818 25394
rect 23438 25342 23490 25394
rect 26014 25342 26066 25394
rect 26686 25342 26738 25394
rect 28590 25342 28642 25394
rect 29150 25342 29202 25394
rect 29486 25342 29538 25394
rect 2046 25230 2098 25282
rect 2494 25230 2546 25282
rect 19182 25230 19234 25282
rect 37662 25678 37714 25730
rect 37886 25342 37938 25394
rect 27134 25230 27186 25282
rect 37326 25230 37378 25282
rect 37662 25230 37714 25282
rect 38222 25230 38274 25282
rect 10538 25062 10590 25114
rect 10642 25062 10694 25114
rect 10746 25062 10798 25114
rect 19862 25062 19914 25114
rect 19966 25062 20018 25114
rect 20070 25062 20122 25114
rect 29186 25062 29238 25114
rect 29290 25062 29342 25114
rect 29394 25062 29446 25114
rect 38510 25062 38562 25114
rect 38614 25062 38666 25114
rect 38718 25062 38770 25114
rect 17726 24894 17778 24946
rect 18958 24894 19010 24946
rect 20190 24894 20242 24946
rect 21758 24894 21810 24946
rect 22206 24894 22258 24946
rect 23438 24894 23490 24946
rect 24110 24894 24162 24946
rect 25790 24894 25842 24946
rect 26686 24894 26738 24946
rect 27134 24894 27186 24946
rect 28366 24894 28418 24946
rect 29262 24894 29314 24946
rect 30158 24894 30210 24946
rect 1710 24782 1762 24834
rect 21086 24782 21138 24834
rect 21310 24782 21362 24834
rect 38222 24782 38274 24834
rect 2046 24670 2098 24722
rect 17950 24670 18002 24722
rect 18398 24670 18450 24722
rect 19294 24670 19346 24722
rect 19854 24670 19906 24722
rect 20526 24670 20578 24722
rect 21198 24670 21250 24722
rect 23102 24670 23154 24722
rect 23774 24670 23826 24722
rect 26126 24670 26178 24722
rect 27806 24670 27858 24722
rect 28702 24670 28754 24722
rect 29710 24670 29762 24722
rect 37998 24670 38050 24722
rect 2494 24558 2546 24610
rect 25230 24558 25282 24610
rect 18622 24446 18674 24498
rect 19518 24446 19570 24498
rect 25454 24446 25506 24498
rect 26350 24446 26402 24498
rect 28030 24446 28082 24498
rect 28926 24446 28978 24498
rect 5876 24278 5928 24330
rect 5980 24278 6032 24330
rect 6084 24278 6136 24330
rect 15200 24278 15252 24330
rect 15304 24278 15356 24330
rect 15408 24278 15460 24330
rect 24524 24278 24576 24330
rect 24628 24278 24680 24330
rect 24732 24278 24784 24330
rect 33848 24278 33900 24330
rect 33952 24278 34004 24330
rect 34056 24278 34108 24330
rect 17614 24110 17666 24162
rect 17950 24110 18002 24162
rect 18286 24110 18338 24162
rect 18622 24110 18674 24162
rect 22542 24110 22594 24162
rect 24670 24110 24722 24162
rect 26014 24110 26066 24162
rect 27582 24110 27634 24162
rect 29374 24110 29426 24162
rect 16606 23998 16658 24050
rect 17054 23998 17106 24050
rect 17390 23998 17442 24050
rect 20078 23998 20130 24050
rect 29150 23998 29202 24050
rect 18846 23886 18898 23938
rect 19518 23886 19570 23938
rect 22094 23886 22146 23938
rect 23774 23886 23826 23938
rect 24894 23886 24946 23938
rect 25790 23886 25842 23938
rect 27358 23886 27410 23938
rect 2046 23774 2098 23826
rect 19294 23774 19346 23826
rect 21870 23774 21922 23826
rect 21982 23774 22034 23826
rect 23998 23774 24050 23826
rect 25342 23774 25394 23826
rect 26350 23774 26402 23826
rect 26686 23774 26738 23826
rect 27022 23774 27074 23826
rect 27918 23774 27970 23826
rect 28254 23774 28306 23826
rect 28590 23774 28642 23826
rect 29710 23774 29762 23826
rect 30046 23774 30098 23826
rect 30382 23774 30434 23826
rect 37886 23774 37938 23826
rect 1710 23662 1762 23714
rect 21422 23662 21474 23714
rect 24334 23662 24386 23714
rect 38222 23662 38274 23714
rect 10538 23494 10590 23546
rect 10642 23494 10694 23546
rect 10746 23494 10798 23546
rect 19862 23494 19914 23546
rect 19966 23494 20018 23546
rect 20070 23494 20122 23546
rect 29186 23494 29238 23546
rect 29290 23494 29342 23546
rect 29394 23494 29446 23546
rect 38510 23494 38562 23546
rect 38614 23494 38666 23546
rect 38718 23494 38770 23546
rect 17726 23326 17778 23378
rect 22542 23326 22594 23378
rect 23886 23326 23938 23378
rect 25566 23326 25618 23378
rect 26014 23326 26066 23378
rect 28142 23326 28194 23378
rect 30158 23326 30210 23378
rect 1710 23214 1762 23266
rect 19742 23214 19794 23266
rect 20414 23214 20466 23266
rect 21086 23214 21138 23266
rect 22094 23214 22146 23266
rect 23214 23214 23266 23266
rect 28926 23214 28978 23266
rect 38222 23214 38274 23266
rect 2046 23102 2098 23154
rect 18062 23102 18114 23154
rect 19406 23102 19458 23154
rect 20190 23102 20242 23154
rect 20862 23102 20914 23154
rect 21758 23102 21810 23154
rect 21982 23102 22034 23154
rect 22878 23102 22930 23154
rect 23550 23102 23602 23154
rect 25342 23102 25394 23154
rect 28366 23102 28418 23154
rect 37886 23102 37938 23154
rect 5876 22710 5928 22762
rect 5980 22710 6032 22762
rect 6084 22710 6136 22762
rect 15200 22710 15252 22762
rect 15304 22710 15356 22762
rect 15408 22710 15460 22762
rect 24524 22710 24576 22762
rect 24628 22710 24680 22762
rect 24732 22710 24784 22762
rect 33848 22710 33900 22762
rect 33952 22710 34004 22762
rect 34056 22710 34108 22762
rect 18286 22542 18338 22594
rect 19294 22542 19346 22594
rect 22430 22542 22482 22594
rect 16718 22430 16770 22482
rect 17054 22430 17106 22482
rect 17390 22430 17442 22482
rect 18846 22430 18898 22482
rect 19854 22430 19906 22482
rect 20302 22430 20354 22482
rect 20750 22430 20802 22482
rect 17614 22318 17666 22370
rect 18622 22318 18674 22370
rect 19630 22318 19682 22370
rect 21646 22318 21698 22370
rect 25118 22318 25170 22370
rect 26238 22318 26290 22370
rect 29374 22318 29426 22370
rect 1710 22206 1762 22258
rect 2046 22206 2098 22258
rect 2718 22206 2770 22258
rect 21870 22206 21922 22258
rect 21982 22206 22034 22258
rect 25230 22206 25282 22258
rect 25342 22206 25394 22258
rect 26350 22206 26402 22258
rect 26462 22206 26514 22258
rect 26910 22206 26962 22258
rect 27246 22206 27298 22258
rect 27582 22206 27634 22258
rect 29262 22206 29314 22258
rect 29486 22206 29538 22258
rect 29934 22206 29986 22258
rect 30270 22206 30322 22258
rect 30606 22206 30658 22258
rect 30942 22206 30994 22258
rect 31278 22206 31330 22258
rect 37214 22206 37266 22258
rect 37886 22206 37938 22258
rect 38222 22206 38274 22258
rect 2382 22094 2434 22146
rect 17950 22094 18002 22146
rect 25790 22094 25842 22146
rect 37550 22094 37602 22146
rect 10538 21926 10590 21978
rect 10642 21926 10694 21978
rect 10746 21926 10798 21978
rect 19862 21926 19914 21978
rect 19966 21926 20018 21978
rect 20070 21926 20122 21978
rect 29186 21926 29238 21978
rect 29290 21926 29342 21978
rect 29394 21926 29446 21978
rect 38510 21926 38562 21978
rect 38614 21926 38666 21978
rect 38718 21926 38770 21978
rect 14702 21758 14754 21810
rect 15374 21758 15426 21810
rect 17726 21758 17778 21810
rect 18846 21758 18898 21810
rect 20078 21758 20130 21810
rect 20974 21758 21026 21810
rect 21422 21758 21474 21810
rect 22430 21758 22482 21810
rect 23102 21758 23154 21810
rect 26126 21758 26178 21810
rect 28478 21758 28530 21810
rect 29598 21758 29650 21810
rect 30270 21758 30322 21810
rect 1710 21646 1762 21698
rect 12350 21646 12402 21698
rect 21758 21646 21810 21698
rect 21870 21646 21922 21698
rect 21982 21646 22034 21698
rect 24446 21646 24498 21698
rect 25790 21646 25842 21698
rect 26798 21646 26850 21698
rect 27246 21646 27298 21698
rect 27470 21646 27522 21698
rect 29038 21646 29090 21698
rect 29150 21646 29202 21698
rect 38222 21646 38274 21698
rect 2046 21534 2098 21586
rect 12574 21534 12626 21586
rect 14926 21534 14978 21586
rect 15598 21534 15650 21586
rect 17950 21534 18002 21586
rect 18510 21534 18562 21586
rect 19182 21534 19234 21586
rect 19406 21534 19458 21586
rect 20302 21534 20354 21586
rect 22766 21534 22818 21586
rect 24334 21534 24386 21586
rect 24670 21534 24722 21586
rect 26462 21534 26514 21586
rect 27358 21534 27410 21586
rect 28814 21534 28866 21586
rect 29934 21534 29986 21586
rect 37886 21534 37938 21586
rect 19742 21422 19794 21474
rect 25454 21422 25506 21474
rect 23886 21310 23938 21362
rect 27918 21310 27970 21362
rect 5876 21142 5928 21194
rect 5980 21142 6032 21194
rect 6084 21142 6136 21194
rect 15200 21142 15252 21194
rect 15304 21142 15356 21194
rect 15408 21142 15460 21194
rect 24524 21142 24576 21194
rect 24628 21142 24680 21194
rect 24732 21142 24784 21194
rect 33848 21142 33900 21194
rect 33952 21142 34004 21194
rect 34056 21142 34108 21194
rect 12350 20974 12402 21026
rect 14702 20974 14754 21026
rect 22206 20974 22258 21026
rect 29934 20974 29986 21026
rect 15822 20862 15874 20914
rect 30382 20862 30434 20914
rect 11790 20750 11842 20802
rect 12014 20750 12066 20802
rect 13918 20750 13970 20802
rect 16942 20750 16994 20802
rect 17502 20750 17554 20802
rect 18174 20750 18226 20802
rect 19070 20750 19122 20802
rect 21422 20750 21474 20802
rect 21646 20750 21698 20802
rect 21758 20750 21810 20802
rect 22766 20750 22818 20802
rect 24110 20750 24162 20802
rect 25454 20750 25506 20802
rect 25566 20750 25618 20802
rect 27918 20750 27970 20802
rect 29262 20750 29314 20802
rect 29374 20750 29426 20802
rect 29486 20750 29538 20802
rect 37998 20750 38050 20802
rect 2046 20638 2098 20690
rect 11118 20638 11170 20690
rect 11454 20638 11506 20690
rect 14142 20638 14194 20690
rect 14254 20638 14306 20690
rect 16270 20638 16322 20690
rect 16382 20638 16434 20690
rect 16494 20638 16546 20690
rect 17950 20638 18002 20690
rect 18846 20638 18898 20690
rect 19966 20638 20018 20690
rect 20414 20638 20466 20690
rect 22542 20638 22594 20690
rect 23214 20638 23266 20690
rect 23550 20638 23602 20690
rect 24446 20638 24498 20690
rect 25342 20638 25394 20690
rect 26014 20638 26066 20690
rect 26350 20638 26402 20690
rect 27022 20638 27074 20690
rect 27358 20638 27410 20690
rect 28142 20638 28194 20690
rect 1710 20526 1762 20578
rect 10782 20526 10834 20578
rect 13582 20526 13634 20578
rect 17278 20526 17330 20578
rect 19630 20526 19682 20578
rect 20750 20526 20802 20578
rect 26686 20526 26738 20578
rect 38222 20526 38274 20578
rect 10538 20358 10590 20410
rect 10642 20358 10694 20410
rect 10746 20358 10798 20410
rect 19862 20358 19914 20410
rect 19966 20358 20018 20410
rect 20070 20358 20122 20410
rect 29186 20358 29238 20410
rect 29290 20358 29342 20410
rect 29394 20358 29446 20410
rect 38510 20358 38562 20410
rect 38614 20358 38666 20410
rect 38718 20358 38770 20410
rect 11566 20190 11618 20242
rect 16158 20190 16210 20242
rect 17950 20190 18002 20242
rect 18510 20190 18562 20242
rect 20526 20190 20578 20242
rect 22206 20190 22258 20242
rect 23662 20190 23714 20242
rect 24334 20190 24386 20242
rect 25790 20190 25842 20242
rect 1710 20078 1762 20130
rect 10782 20078 10834 20130
rect 14142 20078 14194 20130
rect 14254 20078 14306 20130
rect 14702 20078 14754 20130
rect 15262 20078 15314 20130
rect 15374 20078 15426 20130
rect 19182 20078 19234 20130
rect 19966 20078 20018 20130
rect 21534 20078 21586 20130
rect 21646 20078 21698 20130
rect 21758 20078 21810 20130
rect 23998 20078 24050 20130
rect 26350 20078 26402 20130
rect 26686 20078 26738 20130
rect 27022 20078 27074 20130
rect 28254 20078 28306 20130
rect 28926 20078 28978 20130
rect 30382 20078 30434 20130
rect 37886 20078 37938 20130
rect 38222 20078 38274 20130
rect 2046 19966 2098 20018
rect 12126 19966 12178 20018
rect 14030 19966 14082 20018
rect 15038 19966 15090 20018
rect 16494 19966 16546 20018
rect 18958 19966 19010 20018
rect 19630 19966 19682 20018
rect 22654 19966 22706 20018
rect 23438 19966 23490 20018
rect 26014 19966 26066 20018
rect 27918 19966 27970 20018
rect 28590 19966 28642 20018
rect 30046 19966 30098 20018
rect 11230 19854 11282 19906
rect 13022 19854 13074 19906
rect 13582 19854 13634 19906
rect 17390 19854 17442 19906
rect 18398 19854 18450 19906
rect 30942 19854 30994 19906
rect 11902 19742 11954 19794
rect 12462 19742 12514 19794
rect 12798 19742 12850 19794
rect 15822 19742 15874 19794
rect 17614 19742 17666 19794
rect 5876 19574 5928 19626
rect 5980 19574 6032 19626
rect 6084 19574 6136 19626
rect 15200 19574 15252 19626
rect 15304 19574 15356 19626
rect 15408 19574 15460 19626
rect 24524 19574 24576 19626
rect 24628 19574 24680 19626
rect 24732 19574 24784 19626
rect 33848 19574 33900 19626
rect 33952 19574 34004 19626
rect 34056 19574 34108 19626
rect 27918 19406 27970 19458
rect 30046 19406 30098 19458
rect 11566 19294 11618 19346
rect 13582 19294 13634 19346
rect 18958 19294 19010 19346
rect 22542 19294 22594 19346
rect 2046 19182 2098 19234
rect 12238 19182 12290 19234
rect 12798 19182 12850 19234
rect 15262 19182 15314 19234
rect 17166 19182 17218 19234
rect 18510 19182 18562 19234
rect 20638 19182 20690 19234
rect 22878 19182 22930 19234
rect 26014 19182 26066 19234
rect 27470 19182 27522 19234
rect 29374 19182 29426 19234
rect 30382 19182 30434 19234
rect 37886 19182 37938 19234
rect 11902 19070 11954 19122
rect 14926 19070 14978 19122
rect 15934 19070 15986 19122
rect 18174 19070 18226 19122
rect 18846 19070 18898 19122
rect 19742 19070 19794 19122
rect 21534 19070 21586 19122
rect 21870 19070 21922 19122
rect 23102 19070 23154 19122
rect 23214 19070 23266 19122
rect 23998 19070 24050 19122
rect 24334 19070 24386 19122
rect 24670 19070 24722 19122
rect 25342 19070 25394 19122
rect 27246 19070 27298 19122
rect 27358 19070 27410 19122
rect 29486 19070 29538 19122
rect 29598 19070 29650 19122
rect 30606 19070 30658 19122
rect 30718 19070 30770 19122
rect 31166 19070 31218 19122
rect 31502 19070 31554 19122
rect 1710 18958 1762 19010
rect 12574 18958 12626 19010
rect 15598 18958 15650 19010
rect 16942 18958 16994 19010
rect 17726 18958 17778 19010
rect 19070 18958 19122 19010
rect 20078 18958 20130 19010
rect 20414 18958 20466 19010
rect 23662 18958 23714 19010
rect 25006 18958 25058 19010
rect 25678 18958 25730 19010
rect 26350 18958 26402 19010
rect 28366 18958 28418 19010
rect 31838 18958 31890 19010
rect 32398 18958 32450 19010
rect 38222 18958 38274 19010
rect 10538 18790 10590 18842
rect 10642 18790 10694 18842
rect 10746 18790 10798 18842
rect 19862 18790 19914 18842
rect 19966 18790 20018 18842
rect 20070 18790 20122 18842
rect 29186 18790 29238 18842
rect 29290 18790 29342 18842
rect 29394 18790 29446 18842
rect 38510 18790 38562 18842
rect 38614 18790 38666 18842
rect 38718 18790 38770 18842
rect 12462 18622 12514 18674
rect 13470 18622 13522 18674
rect 16830 18622 16882 18674
rect 19182 18622 19234 18674
rect 21534 18622 21586 18674
rect 23438 18622 23490 18674
rect 1710 18510 1762 18562
rect 10894 18510 10946 18562
rect 13918 18510 13970 18562
rect 15374 18510 15426 18562
rect 18174 18510 18226 18562
rect 19854 18510 19906 18562
rect 20974 18510 21026 18562
rect 24446 18510 24498 18562
rect 26574 18510 26626 18562
rect 27470 18510 27522 18562
rect 28926 18510 28978 18562
rect 29038 18510 29090 18562
rect 30046 18510 30098 18562
rect 30158 18510 30210 18562
rect 31278 18510 31330 18562
rect 38222 18510 38274 18562
rect 2046 18398 2098 18450
rect 10558 18398 10610 18450
rect 11230 18398 11282 18450
rect 11566 18398 11618 18450
rect 12126 18398 12178 18450
rect 13022 18398 13074 18450
rect 14030 18398 14082 18450
rect 14142 18398 14194 18450
rect 14590 18398 14642 18450
rect 15710 18398 15762 18450
rect 16046 18398 16098 18450
rect 16270 18398 16322 18450
rect 16382 18398 16434 18450
rect 17838 18398 17890 18450
rect 18510 18398 18562 18450
rect 18846 18398 18898 18450
rect 19518 18398 19570 18450
rect 20862 18398 20914 18450
rect 21086 18398 21138 18450
rect 23102 18398 23154 18450
rect 24110 18398 24162 18450
rect 26462 18398 26514 18450
rect 26798 18398 26850 18450
rect 27134 18398 27186 18450
rect 27358 18398 27410 18450
rect 27918 18398 27970 18450
rect 28814 18398 28866 18450
rect 29934 18398 29986 18450
rect 30606 18398 30658 18450
rect 30942 18398 30994 18450
rect 37886 18398 37938 18450
rect 15038 18286 15090 18338
rect 17726 18286 17778 18338
rect 21982 18286 22034 18338
rect 22766 18286 22818 18338
rect 28366 18286 28418 18338
rect 31726 18286 31778 18338
rect 11902 18174 11954 18226
rect 12798 18174 12850 18226
rect 26014 18174 26066 18226
rect 29486 18174 29538 18226
rect 5876 18006 5928 18058
rect 5980 18006 6032 18058
rect 6084 18006 6136 18058
rect 15200 18006 15252 18058
rect 15304 18006 15356 18058
rect 15408 18006 15460 18058
rect 24524 18006 24576 18058
rect 24628 18006 24680 18058
rect 24732 18006 24784 18058
rect 33848 18006 33900 18058
rect 33952 18006 34004 18058
rect 34056 18006 34108 18058
rect 11902 17838 11954 17890
rect 16830 17838 16882 17890
rect 23774 17838 23826 17890
rect 21310 17726 21362 17778
rect 30606 17726 30658 17778
rect 2718 17614 2770 17666
rect 11678 17614 11730 17666
rect 13806 17614 13858 17666
rect 14030 17614 14082 17666
rect 14142 17614 14194 17666
rect 14590 17614 14642 17666
rect 15150 17614 15202 17666
rect 16606 17614 16658 17666
rect 17166 17614 17218 17666
rect 17726 17614 17778 17666
rect 19966 17614 20018 17666
rect 20526 17614 20578 17666
rect 21758 17614 21810 17666
rect 22094 17614 22146 17666
rect 23214 17614 23266 17666
rect 23326 17614 23378 17666
rect 26462 17614 26514 17666
rect 27358 17614 27410 17666
rect 27470 17614 27522 17666
rect 29598 17614 29650 17666
rect 37886 17614 37938 17666
rect 1710 17502 1762 17554
rect 3166 17502 3218 17554
rect 12910 17502 12962 17554
rect 14926 17502 14978 17554
rect 15598 17502 15650 17554
rect 15934 17502 15986 17554
rect 21870 17502 21922 17554
rect 22654 17502 22706 17554
rect 23102 17502 23154 17554
rect 24334 17502 24386 17554
rect 24670 17502 24722 17554
rect 27246 17502 27298 17554
rect 27918 17502 27970 17554
rect 28254 17502 28306 17554
rect 37214 17502 37266 17554
rect 38222 17502 38274 17554
rect 2046 17390 2098 17442
rect 2382 17390 2434 17442
rect 11342 17390 11394 17442
rect 12238 17390 12290 17442
rect 12574 17390 12626 17442
rect 17502 17390 17554 17442
rect 18286 17390 18338 17442
rect 18958 17390 19010 17442
rect 19406 17390 19458 17442
rect 19742 17390 19794 17442
rect 20750 17390 20802 17442
rect 25006 17390 25058 17442
rect 26798 17390 26850 17442
rect 28590 17390 28642 17442
rect 29262 17390 29314 17442
rect 29934 17390 29986 17442
rect 37550 17390 37602 17442
rect 10538 17222 10590 17274
rect 10642 17222 10694 17274
rect 10746 17222 10798 17274
rect 19862 17222 19914 17274
rect 19966 17222 20018 17274
rect 20070 17222 20122 17274
rect 29186 17222 29238 17274
rect 29290 17222 29342 17274
rect 29394 17222 29446 17274
rect 38510 17222 38562 17274
rect 38614 17222 38666 17274
rect 38718 17222 38770 17274
rect 13470 17054 13522 17106
rect 13694 17054 13746 17106
rect 16494 17054 16546 17106
rect 17950 17054 18002 17106
rect 19630 17054 19682 17106
rect 23998 17054 24050 17106
rect 24670 17054 24722 17106
rect 26910 17054 26962 17106
rect 1710 16942 1762 16994
rect 12126 16942 12178 16994
rect 12910 16942 12962 16994
rect 14142 16942 14194 16994
rect 14366 16942 14418 16994
rect 18286 16942 18338 16994
rect 18622 16942 18674 16994
rect 18958 16942 19010 16994
rect 20078 16942 20130 16994
rect 21086 16942 21138 16994
rect 21198 16942 21250 16994
rect 22318 16942 22370 16994
rect 23438 16942 23490 16994
rect 23550 16942 23602 16994
rect 25566 16942 25618 16994
rect 28478 16942 28530 16994
rect 28814 16942 28866 16994
rect 29150 16942 29202 16994
rect 31950 16942 32002 16994
rect 37886 16942 37938 16994
rect 38222 16942 38274 16994
rect 2046 16830 2098 16882
rect 12350 16830 12402 16882
rect 14254 16830 14306 16882
rect 15934 16830 15986 16882
rect 16718 16830 16770 16882
rect 17614 16830 17666 16882
rect 19182 16830 19234 16882
rect 20190 16830 20242 16882
rect 20414 16830 20466 16882
rect 20974 16830 21026 16882
rect 21646 16830 21698 16882
rect 21982 16830 22034 16882
rect 22878 16830 22930 16882
rect 23326 16830 23378 16882
rect 24334 16830 24386 16882
rect 25342 16830 25394 16882
rect 26462 16830 26514 16882
rect 27806 16830 27858 16882
rect 28142 16830 28194 16882
rect 29822 16830 29874 16882
rect 30718 16830 30770 16882
rect 31278 16830 31330 16882
rect 31614 16830 31666 16882
rect 32398 16830 32450 16882
rect 15374 16718 15426 16770
rect 26238 16718 26290 16770
rect 27246 16718 27298 16770
rect 27470 16718 27522 16770
rect 15598 16606 15650 16658
rect 25902 16606 25954 16658
rect 30046 16606 30098 16658
rect 30382 16606 30434 16658
rect 30942 16606 30994 16658
rect 5876 16438 5928 16490
rect 5980 16438 6032 16490
rect 6084 16438 6136 16490
rect 15200 16438 15252 16490
rect 15304 16438 15356 16490
rect 15408 16438 15460 16490
rect 24524 16438 24576 16490
rect 24628 16438 24680 16490
rect 24732 16438 24784 16490
rect 33848 16438 33900 16490
rect 33952 16438 34004 16490
rect 34056 16438 34108 16490
rect 19182 16270 19234 16322
rect 19518 16270 19570 16322
rect 21534 16270 21586 16322
rect 23886 16270 23938 16322
rect 28254 16270 28306 16322
rect 28478 16270 28530 16322
rect 21310 16158 21362 16210
rect 24222 16158 24274 16210
rect 25902 16158 25954 16210
rect 1934 16046 1986 16098
rect 18398 16046 18450 16098
rect 19742 16046 19794 16098
rect 22430 16046 22482 16098
rect 23102 16046 23154 16098
rect 23326 16046 23378 16098
rect 23438 16046 23490 16098
rect 24446 16046 24498 16098
rect 26238 16046 26290 16098
rect 30494 16046 30546 16098
rect 37886 16046 37938 16098
rect 16718 15934 16770 15986
rect 22766 15934 22818 15986
rect 24782 15934 24834 15986
rect 25118 15934 25170 15986
rect 26574 15934 26626 15986
rect 27694 15934 27746 15986
rect 1710 15822 1762 15874
rect 20078 15822 20130 15874
rect 20414 15822 20466 15874
rect 21870 15822 21922 15874
rect 25454 15822 25506 15874
rect 28030 15822 28082 15874
rect 28478 15822 28530 15874
rect 30830 15822 30882 15874
rect 38222 15822 38274 15874
rect 10538 15654 10590 15706
rect 10642 15654 10694 15706
rect 10746 15654 10798 15706
rect 19862 15654 19914 15706
rect 19966 15654 20018 15706
rect 20070 15654 20122 15706
rect 29186 15654 29238 15706
rect 29290 15654 29342 15706
rect 29394 15654 29446 15706
rect 38510 15654 38562 15706
rect 38614 15654 38666 15706
rect 38718 15654 38770 15706
rect 27694 15486 27746 15538
rect 1710 15374 1762 15426
rect 20190 15374 20242 15426
rect 24110 15374 24162 15426
rect 25566 15374 25618 15426
rect 31054 15374 31106 15426
rect 38222 15374 38274 15426
rect 2046 15262 2098 15314
rect 14030 15262 14082 15314
rect 17390 15262 17442 15314
rect 23214 15262 23266 15314
rect 23774 15262 23826 15314
rect 24334 15262 24386 15314
rect 25230 15262 25282 15314
rect 27134 15262 27186 15314
rect 28030 15262 28082 15314
rect 28254 15262 28306 15314
rect 29150 15262 29202 15314
rect 29822 15262 29874 15314
rect 30046 15262 30098 15314
rect 30382 15262 30434 15314
rect 30718 15262 30770 15314
rect 31502 15262 31554 15314
rect 37886 15262 37938 15314
rect 14702 15150 14754 15202
rect 16830 15150 16882 15202
rect 23438 15150 23490 15202
rect 27358 15150 27410 15202
rect 28926 15150 28978 15202
rect 26798 15038 26850 15090
rect 29486 15038 29538 15090
rect 5876 14870 5928 14922
rect 5980 14870 6032 14922
rect 6084 14870 6136 14922
rect 15200 14870 15252 14922
rect 15304 14870 15356 14922
rect 15408 14870 15460 14922
rect 24524 14870 24576 14922
rect 24628 14870 24680 14922
rect 24732 14870 24784 14922
rect 33848 14870 33900 14922
rect 33952 14870 34004 14922
rect 34056 14870 34108 14922
rect 18286 14702 18338 14754
rect 18510 14702 18562 14754
rect 18958 14702 19010 14754
rect 20414 14702 20466 14754
rect 17054 14590 17106 14642
rect 28478 14590 28530 14642
rect 14254 14478 14306 14530
rect 18062 14478 18114 14530
rect 19406 14478 19458 14530
rect 19742 14478 19794 14530
rect 20190 14478 20242 14530
rect 21870 14478 21922 14530
rect 27134 14478 27186 14530
rect 29486 14478 29538 14530
rect 1710 14366 1762 14418
rect 14926 14366 14978 14418
rect 17614 14366 17666 14418
rect 19182 14366 19234 14418
rect 23550 14366 23602 14418
rect 27470 14366 27522 14418
rect 37886 14366 37938 14418
rect 2046 14254 2098 14306
rect 2494 14254 2546 14306
rect 17726 14254 17778 14306
rect 19070 14254 19122 14306
rect 20750 14254 20802 14306
rect 29822 14254 29874 14306
rect 38222 14254 38274 14306
rect 10538 14086 10590 14138
rect 10642 14086 10694 14138
rect 10746 14086 10798 14138
rect 19862 14086 19914 14138
rect 19966 14086 20018 14138
rect 20070 14086 20122 14138
rect 29186 14086 29238 14138
rect 29290 14086 29342 14138
rect 29394 14086 29446 14138
rect 38510 14086 38562 14138
rect 38614 14086 38666 14138
rect 38718 14086 38770 14138
rect 2046 13918 2098 13970
rect 15822 13918 15874 13970
rect 19854 13918 19906 13970
rect 15486 13806 15538 13858
rect 19518 13806 19570 13858
rect 19966 13806 20018 13858
rect 20974 13806 21026 13858
rect 25566 13806 25618 13858
rect 38222 13806 38274 13858
rect 1710 13694 1762 13746
rect 18062 13694 18114 13746
rect 18510 13694 18562 13746
rect 18958 13694 19010 13746
rect 19182 13694 19234 13746
rect 20750 13694 20802 13746
rect 21646 13694 21698 13746
rect 22990 13694 23042 13746
rect 23886 13694 23938 13746
rect 24222 13694 24274 13746
rect 25230 13694 25282 13746
rect 37886 13694 37938 13746
rect 2494 13582 2546 13634
rect 16830 13582 16882 13634
rect 17614 13582 17666 13634
rect 21310 13582 21362 13634
rect 21870 13582 21922 13634
rect 22318 13582 22370 13634
rect 22766 13582 22818 13634
rect 23662 13582 23714 13634
rect 24670 13582 24722 13634
rect 17726 13470 17778 13522
rect 18286 13470 18338 13522
rect 23326 13470 23378 13522
rect 5876 13302 5928 13354
rect 5980 13302 6032 13354
rect 6084 13302 6136 13354
rect 15200 13302 15252 13354
rect 15304 13302 15356 13354
rect 15408 13302 15460 13354
rect 24524 13302 24576 13354
rect 24628 13302 24680 13354
rect 24732 13302 24784 13354
rect 33848 13302 33900 13354
rect 33952 13302 34004 13354
rect 34056 13302 34108 13354
rect 17726 12910 17778 12962
rect 17950 12910 18002 12962
rect 21982 12910 22034 12962
rect 23326 12910 23378 12962
rect 37214 12910 37266 12962
rect 1710 12798 1762 12850
rect 2046 12798 2098 12850
rect 2494 12798 2546 12850
rect 37886 12798 37938 12850
rect 38222 12798 38274 12850
rect 17390 12686 17442 12738
rect 17502 12686 17554 12738
rect 21422 12686 21474 12738
rect 21758 12686 21810 12738
rect 23550 12686 23602 12738
rect 24446 12686 24498 12738
rect 37550 12686 37602 12738
rect 10538 12518 10590 12570
rect 10642 12518 10694 12570
rect 10746 12518 10798 12570
rect 19862 12518 19914 12570
rect 19966 12518 20018 12570
rect 20070 12518 20122 12570
rect 29186 12518 29238 12570
rect 29290 12518 29342 12570
rect 29394 12518 29446 12570
rect 38510 12518 38562 12570
rect 38614 12518 38666 12570
rect 38718 12518 38770 12570
rect 37886 12350 37938 12402
rect 37662 12126 37714 12178
rect 38222 12126 38274 12178
rect 5876 11734 5928 11786
rect 5980 11734 6032 11786
rect 6084 11734 6136 11786
rect 15200 11734 15252 11786
rect 15304 11734 15356 11786
rect 15408 11734 15460 11786
rect 24524 11734 24576 11786
rect 24628 11734 24680 11786
rect 24732 11734 24784 11786
rect 33848 11734 33900 11786
rect 33952 11734 34004 11786
rect 34056 11734 34108 11786
rect 37886 11230 37938 11282
rect 38222 11118 38274 11170
rect 10538 10950 10590 11002
rect 10642 10950 10694 11002
rect 10746 10950 10798 11002
rect 19862 10950 19914 11002
rect 19966 10950 20018 11002
rect 20070 10950 20122 11002
rect 29186 10950 29238 11002
rect 29290 10950 29342 11002
rect 29394 10950 29446 11002
rect 38510 10950 38562 11002
rect 38614 10950 38666 11002
rect 38718 10950 38770 11002
rect 38222 10670 38274 10722
rect 37886 10558 37938 10610
rect 5876 10166 5928 10218
rect 5980 10166 6032 10218
rect 6084 10166 6136 10218
rect 15200 10166 15252 10218
rect 15304 10166 15356 10218
rect 15408 10166 15460 10218
rect 24524 10166 24576 10218
rect 24628 10166 24680 10218
rect 24732 10166 24784 10218
rect 33848 10166 33900 10218
rect 33952 10166 34004 10218
rect 34056 10166 34108 10218
rect 37886 9662 37938 9714
rect 38222 9662 38274 9714
rect 37662 9550 37714 9602
rect 10538 9382 10590 9434
rect 10642 9382 10694 9434
rect 10746 9382 10798 9434
rect 19862 9382 19914 9434
rect 19966 9382 20018 9434
rect 20070 9382 20122 9434
rect 29186 9382 29238 9434
rect 29290 9382 29342 9434
rect 29394 9382 29446 9434
rect 38510 9382 38562 9434
rect 38614 9382 38666 9434
rect 38718 9382 38770 9434
rect 37886 9102 37938 9154
rect 38222 9102 38274 9154
rect 5876 8598 5928 8650
rect 5980 8598 6032 8650
rect 6084 8598 6136 8650
rect 15200 8598 15252 8650
rect 15304 8598 15356 8650
rect 15408 8598 15460 8650
rect 24524 8598 24576 8650
rect 24628 8598 24680 8650
rect 24732 8598 24784 8650
rect 33848 8598 33900 8650
rect 33952 8598 34004 8650
rect 34056 8598 34108 8650
rect 37214 8094 37266 8146
rect 37886 8094 37938 8146
rect 38222 8094 38274 8146
rect 36430 7982 36482 8034
rect 37550 7982 37602 8034
rect 10538 7814 10590 7866
rect 10642 7814 10694 7866
rect 10746 7814 10798 7866
rect 19862 7814 19914 7866
rect 19966 7814 20018 7866
rect 20070 7814 20122 7866
rect 29186 7814 29238 7866
rect 29290 7814 29342 7866
rect 29394 7814 29446 7866
rect 38510 7814 38562 7866
rect 38614 7814 38666 7866
rect 38718 7814 38770 7866
rect 37662 7646 37714 7698
rect 38222 7534 38274 7586
rect 37886 7422 37938 7474
rect 37214 7310 37266 7362
rect 5876 7030 5928 7082
rect 5980 7030 6032 7082
rect 6084 7030 6136 7082
rect 15200 7030 15252 7082
rect 15304 7030 15356 7082
rect 15408 7030 15460 7082
rect 24524 7030 24576 7082
rect 24628 7030 24680 7082
rect 24732 7030 24784 7082
rect 33848 7030 33900 7082
rect 33952 7030 34004 7082
rect 34056 7030 34108 7082
rect 37550 6526 37602 6578
rect 37886 6526 37938 6578
rect 38222 6414 38274 6466
rect 10538 6246 10590 6298
rect 10642 6246 10694 6298
rect 10746 6246 10798 6298
rect 19862 6246 19914 6298
rect 19966 6246 20018 6298
rect 20070 6246 20122 6298
rect 29186 6246 29238 6298
rect 29290 6246 29342 6298
rect 29394 6246 29446 6298
rect 38510 6246 38562 6298
rect 38614 6246 38666 6298
rect 38718 6246 38770 6298
rect 38222 5966 38274 6018
rect 37886 5854 37938 5906
rect 37662 5742 37714 5794
rect 5876 5462 5928 5514
rect 5980 5462 6032 5514
rect 6084 5462 6136 5514
rect 15200 5462 15252 5514
rect 15304 5462 15356 5514
rect 15408 5462 15460 5514
rect 24524 5462 24576 5514
rect 24628 5462 24680 5514
rect 24732 5462 24784 5514
rect 33848 5462 33900 5514
rect 33952 5462 34004 5514
rect 34056 5462 34108 5514
rect 37550 5070 37602 5122
rect 37998 5070 38050 5122
rect 38222 4846 38274 4898
rect 10538 4678 10590 4730
rect 10642 4678 10694 4730
rect 10746 4678 10798 4730
rect 19862 4678 19914 4730
rect 19966 4678 20018 4730
rect 20070 4678 20122 4730
rect 29186 4678 29238 4730
rect 29290 4678 29342 4730
rect 29394 4678 29446 4730
rect 38510 4678 38562 4730
rect 38614 4678 38666 4730
rect 38718 4678 38770 4730
rect 16382 4398 16434 4450
rect 38222 4398 38274 4450
rect 16606 4286 16658 4338
rect 37886 4286 37938 4338
rect 15934 4174 15986 4226
rect 25678 4174 25730 4226
rect 26350 4174 26402 4226
rect 37662 4174 37714 4226
rect 5876 3894 5928 3946
rect 5980 3894 6032 3946
rect 6084 3894 6136 3946
rect 15200 3894 15252 3946
rect 15304 3894 15356 3946
rect 15408 3894 15460 3946
rect 24524 3894 24576 3946
rect 24628 3894 24680 3946
rect 24732 3894 24784 3946
rect 33848 3894 33900 3946
rect 33952 3894 34004 3946
rect 34056 3894 34108 3946
rect 15486 3502 15538 3554
rect 16046 3502 16098 3554
rect 17278 3502 17330 3554
rect 17950 3502 18002 3554
rect 18622 3502 18674 3554
rect 19294 3502 19346 3554
rect 19854 3502 19906 3554
rect 21422 3502 21474 3554
rect 21982 3502 22034 3554
rect 22766 3502 22818 3554
rect 23326 3502 23378 3554
rect 24782 3502 24834 3554
rect 25566 3502 25618 3554
rect 26238 3502 26290 3554
rect 26798 3502 26850 3554
rect 27470 3502 27522 3554
rect 15710 3390 15762 3442
rect 16382 3390 16434 3442
rect 24110 3390 24162 3442
rect 24558 3390 24610 3442
rect 25230 3390 25282 3442
rect 25902 3390 25954 3442
rect 26574 3390 26626 3442
rect 27246 3390 27298 3442
rect 36430 3390 36482 3442
rect 36990 3390 37042 3442
rect 37214 3390 37266 3442
rect 37550 3390 37602 3442
rect 37886 3390 37938 3442
rect 38222 3390 38274 3442
rect 17502 3278 17554 3330
rect 18174 3278 18226 3330
rect 18846 3278 18898 3330
rect 19518 3278 19570 3330
rect 20190 3278 20242 3330
rect 21086 3278 21138 3330
rect 21758 3278 21810 3330
rect 22430 3278 22482 3330
rect 23102 3278 23154 3330
rect 10538 3110 10590 3162
rect 10642 3110 10694 3162
rect 10746 3110 10798 3162
rect 19862 3110 19914 3162
rect 19966 3110 20018 3162
rect 20070 3110 20122 3162
rect 29186 3110 29238 3162
rect 29290 3110 29342 3162
rect 29394 3110 29446 3162
rect 38510 3110 38562 3162
rect 38614 3110 38666 3162
rect 38718 3110 38770 3162
rect 25566 2494 25618 2546
rect 26350 2494 26402 2546
rect 26798 2494 26850 2546
<< metal2 >>
rect 14784 39200 14896 40000
rect 15456 39200 15568 40000
rect 16128 39200 16240 40000
rect 16800 39200 16912 40000
rect 17472 39200 17584 40000
rect 18144 39200 18256 40000
rect 18816 39200 18928 40000
rect 19488 39200 19600 40000
rect 20160 39200 20272 40000
rect 20832 39200 20944 40000
rect 21504 39200 21616 40000
rect 22176 39200 22288 40000
rect 22848 39200 22960 40000
rect 23520 39200 23632 40000
rect 24192 39200 24304 40000
rect 24864 39200 24976 40000
rect 5874 36876 6138 36886
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 5874 36810 6138 36820
rect 14812 36484 14868 39200
rect 15484 37044 15540 39200
rect 15484 36988 15652 37044
rect 15198 36876 15462 36886
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15198 36810 15462 36820
rect 14812 36482 15316 36484
rect 14812 36430 14814 36482
rect 14866 36430 15316 36482
rect 14812 36428 15316 36430
rect 14812 36418 14868 36428
rect 15036 36258 15092 36270
rect 15036 36206 15038 36258
rect 15090 36206 15092 36258
rect 10536 36092 10800 36102
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10536 36026 10800 36036
rect 5874 35308 6138 35318
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 5874 35242 6138 35252
rect 10536 34524 10800 34534
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10536 34458 10800 34468
rect 5874 33740 6138 33750
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 5874 33674 6138 33684
rect 10536 32956 10800 32966
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10536 32890 10800 32900
rect 5874 32172 6138 32182
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 5874 32106 6138 32116
rect 10536 31388 10800 31398
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10536 31322 10800 31332
rect 5874 30604 6138 30614
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 5874 30538 6138 30548
rect 10536 29820 10800 29830
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10536 29754 10800 29764
rect 5874 29036 6138 29046
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 5874 28970 6138 28980
rect 10536 28252 10800 28262
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10536 28186 10800 28196
rect 5874 27468 6138 27478
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 5874 27402 6138 27412
rect 1820 27074 1876 27086
rect 1820 27022 1822 27074
rect 1874 27022 1876 27074
rect 1820 26852 1876 27022
rect 2492 26962 2548 26974
rect 2492 26910 2494 26962
rect 2546 26910 2548 26962
rect 1708 26402 1764 26414
rect 1708 26350 1710 26402
rect 1762 26350 1764 26402
rect 1708 25620 1764 26350
rect 1820 26292 1876 26796
rect 2044 26852 2100 26862
rect 2492 26852 2548 26910
rect 2044 26850 2436 26852
rect 2044 26798 2046 26850
rect 2098 26798 2436 26850
rect 2044 26796 2436 26798
rect 2044 26786 2100 26796
rect 1820 26226 1876 26236
rect 2044 26290 2100 26302
rect 2044 26238 2046 26290
rect 2098 26238 2100 26290
rect 2044 26068 2100 26238
rect 2268 26068 2324 26078
rect 2044 26066 2324 26068
rect 2044 26014 2270 26066
rect 2322 26014 2324 26066
rect 2044 26012 2324 26014
rect 2268 26002 2324 26012
rect 1708 25554 1764 25564
rect 1820 25506 1876 25518
rect 1820 25454 1822 25506
rect 1874 25454 1876 25506
rect 1820 24948 1876 25454
rect 2380 25508 2436 26796
rect 2492 26786 2548 26796
rect 10536 26684 10800 26694
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10536 26618 10800 26628
rect 2492 26180 2548 26190
rect 2492 26178 2884 26180
rect 2492 26126 2494 26178
rect 2546 26126 2884 26178
rect 2492 26124 2884 26126
rect 2492 26066 2548 26124
rect 2492 26014 2494 26066
rect 2546 26014 2548 26066
rect 2492 26002 2548 26014
rect 2380 25452 2660 25508
rect 2044 25284 2100 25294
rect 1820 24882 1876 24892
rect 1932 25282 2100 25284
rect 1932 25230 2046 25282
rect 2098 25230 2100 25282
rect 1932 25228 2100 25230
rect 1708 24834 1764 24846
rect 1708 24782 1710 24834
rect 1762 24782 1764 24834
rect 1708 24276 1764 24782
rect 1708 24210 1764 24220
rect 1708 23716 1764 23726
rect 1708 23622 1764 23660
rect 1708 23266 1764 23278
rect 1708 23214 1710 23266
rect 1762 23214 1764 23266
rect 1708 22932 1764 23214
rect 1708 22866 1764 22876
rect 1708 22260 1764 22270
rect 1708 22166 1764 22204
rect 1708 21698 1764 21710
rect 1708 21646 1710 21698
rect 1762 21646 1764 21698
rect 1708 20916 1764 21646
rect 1932 21364 1988 25228
rect 2044 25218 2100 25228
rect 2492 25282 2548 25294
rect 2492 25230 2494 25282
rect 2546 25230 2548 25282
rect 2492 24948 2548 25230
rect 2492 24882 2548 24892
rect 2044 24722 2100 24734
rect 2044 24670 2046 24722
rect 2098 24670 2100 24722
rect 2044 24612 2100 24670
rect 2492 24612 2548 24622
rect 2044 24610 2548 24612
rect 2044 24558 2494 24610
rect 2546 24558 2548 24610
rect 2044 24556 2548 24558
rect 2044 23828 2100 23838
rect 2044 23826 2212 23828
rect 2044 23774 2046 23826
rect 2098 23774 2212 23826
rect 2044 23772 2212 23774
rect 2044 23762 2100 23772
rect 2044 23156 2100 23166
rect 2044 23062 2100 23100
rect 2044 22260 2100 22270
rect 2044 22166 2100 22204
rect 2044 21588 2100 21598
rect 2044 21494 2100 21532
rect 1932 21298 1988 21308
rect 1708 20850 1764 20860
rect 2044 20690 2100 20702
rect 2044 20638 2046 20690
rect 2098 20638 2100 20690
rect 1708 20580 1764 20590
rect 1708 20486 1764 20524
rect 2044 20244 2100 20638
rect 2156 20692 2212 23772
rect 2380 22146 2436 22158
rect 2380 22094 2382 22146
rect 2434 22094 2436 22146
rect 2380 21812 2436 22094
rect 2380 21746 2436 21756
rect 2492 20916 2548 24556
rect 2492 20850 2548 20860
rect 2156 20626 2212 20636
rect 2044 20178 2100 20188
rect 1708 20130 1764 20142
rect 1708 20078 1710 20130
rect 1762 20078 1764 20130
rect 1708 19572 1764 20078
rect 2604 20132 2660 25452
rect 2716 22258 2772 22270
rect 2716 22206 2718 22258
rect 2770 22206 2772 22258
rect 2716 21028 2772 22206
rect 2716 20962 2772 20972
rect 2604 20066 2660 20076
rect 2044 20020 2100 20030
rect 2044 19926 2100 19964
rect 1708 19506 1764 19516
rect 2044 19460 2100 19470
rect 2044 19234 2100 19404
rect 2044 19182 2046 19234
rect 2098 19182 2100 19234
rect 2044 19170 2100 19182
rect 2828 19236 2884 26124
rect 5874 25900 6138 25910
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 5874 25834 6138 25844
rect 10536 25116 10800 25126
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10536 25050 10800 25060
rect 5874 24332 6138 24342
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 5874 24266 6138 24276
rect 15036 24052 15092 36206
rect 15260 35922 15316 36428
rect 15372 36372 15428 36382
rect 15596 36372 15652 36988
rect 15372 36370 15652 36372
rect 15372 36318 15374 36370
rect 15426 36318 15652 36370
rect 15372 36316 15652 36318
rect 15708 36370 15764 36382
rect 15708 36318 15710 36370
rect 15762 36318 15764 36370
rect 15372 36306 15428 36316
rect 15260 35870 15262 35922
rect 15314 35870 15316 35922
rect 15260 35858 15316 35870
rect 15198 35308 15462 35318
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15198 35242 15462 35252
rect 15198 33740 15462 33750
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15198 33674 15462 33684
rect 15198 32172 15462 32182
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15198 32106 15462 32116
rect 15198 30604 15462 30614
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15198 30538 15462 30548
rect 15198 29036 15462 29046
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15198 28970 15462 28980
rect 15708 28644 15764 36318
rect 16044 36370 16100 36382
rect 16044 36318 16046 36370
rect 16098 36318 16100 36370
rect 16044 35364 16100 36318
rect 16156 35924 16212 39200
rect 16828 36932 16884 39200
rect 16380 36876 16884 36932
rect 16380 36370 16436 36876
rect 17276 36484 17332 36494
rect 17276 36482 17444 36484
rect 17276 36430 17278 36482
rect 17330 36430 17444 36482
rect 17276 36428 17444 36430
rect 17276 36418 17332 36428
rect 16380 36318 16382 36370
rect 16434 36318 16436 36370
rect 16380 36306 16436 36318
rect 16380 35924 16436 35934
rect 16156 35922 16436 35924
rect 16156 35870 16158 35922
rect 16210 35870 16382 35922
rect 16434 35870 16436 35922
rect 16156 35868 16436 35870
rect 16156 35858 16212 35868
rect 16380 35858 16436 35868
rect 16044 35298 16100 35308
rect 16716 35810 16772 35822
rect 16716 35758 16718 35810
rect 16770 35758 16772 35810
rect 15708 28578 15764 28588
rect 15198 27468 15462 27478
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15198 27402 15462 27412
rect 15198 25900 15462 25910
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15198 25834 15462 25844
rect 15198 24332 15462 24342
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15198 24266 15462 24276
rect 15036 23986 15092 23996
rect 16604 24052 16660 24062
rect 16604 23958 16660 23996
rect 16716 24052 16772 35758
rect 17276 35364 17332 35374
rect 17276 31948 17332 35308
rect 17388 34132 17444 36428
rect 17500 36370 17556 39200
rect 17500 36318 17502 36370
rect 17554 36318 17556 36370
rect 17500 36306 17556 36318
rect 17836 36370 17892 36382
rect 17836 36318 17838 36370
rect 17890 36318 17892 36370
rect 17388 34076 17780 34132
rect 17276 31892 17556 31948
rect 17500 24724 17556 31892
rect 17612 28644 17668 28654
rect 17612 24948 17668 28588
rect 17724 25394 17780 34076
rect 17724 25342 17726 25394
rect 17778 25342 17780 25394
rect 17724 25330 17780 25342
rect 17724 24948 17780 24958
rect 17612 24946 17780 24948
rect 17612 24894 17726 24946
rect 17778 24894 17780 24946
rect 17612 24892 17780 24894
rect 17724 24882 17780 24892
rect 17500 24668 17780 24724
rect 17612 24500 17668 24510
rect 17612 24162 17668 24444
rect 17612 24110 17614 24162
rect 17666 24110 17668 24162
rect 17612 24098 17668 24110
rect 17052 24052 17108 24062
rect 17388 24052 17444 24062
rect 16716 24050 17108 24052
rect 16716 23998 17054 24050
rect 17106 23998 17108 24050
rect 16716 23996 17108 23998
rect 10536 23548 10800 23558
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10536 23482 10800 23492
rect 15596 23156 15652 23166
rect 5874 22764 6138 22774
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 5874 22698 6138 22708
rect 15198 22764 15462 22774
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15198 22698 15462 22708
rect 14700 22260 14756 22270
rect 10536 21980 10800 21990
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10536 21914 10800 21924
rect 14700 21810 14756 22204
rect 14700 21758 14702 21810
rect 14754 21758 14756 21810
rect 14700 21746 14756 21758
rect 15372 21812 15428 21822
rect 15596 21812 15652 23100
rect 16716 22596 16772 23996
rect 17052 23940 17108 23996
rect 17052 23874 17108 23884
rect 17164 23996 17388 24052
rect 16716 22482 16772 22540
rect 16716 22430 16718 22482
rect 16770 22430 16772 22482
rect 16716 22418 16772 22430
rect 17052 22484 17108 22494
rect 17164 22484 17220 23996
rect 17388 23958 17444 23996
rect 17724 23378 17780 24668
rect 17724 23326 17726 23378
rect 17778 23326 17780 23378
rect 17724 23314 17780 23326
rect 17052 22482 17164 22484
rect 17052 22430 17054 22482
rect 17106 22430 17164 22482
rect 17052 22428 17164 22430
rect 17052 22418 17108 22428
rect 17164 22390 17220 22428
rect 17388 22596 17444 22606
rect 17388 22482 17444 22540
rect 17388 22430 17390 22482
rect 17442 22430 17444 22482
rect 17388 22418 17444 22430
rect 17612 22372 17668 22382
rect 17612 22278 17668 22316
rect 15372 21810 15652 21812
rect 15372 21758 15374 21810
rect 15426 21758 15652 21810
rect 15372 21756 15652 21758
rect 17724 21812 17780 21822
rect 17836 21812 17892 36318
rect 18172 36370 18228 39200
rect 18172 36318 18174 36370
rect 18226 36318 18228 36370
rect 18172 36306 18228 36318
rect 18508 36370 18564 36382
rect 18508 36318 18510 36370
rect 18562 36318 18564 36370
rect 18508 34020 18564 36318
rect 18844 36370 18900 39200
rect 18844 36318 18846 36370
rect 18898 36318 18900 36370
rect 18844 36306 18900 36318
rect 19180 36370 19236 36382
rect 19180 36318 19182 36370
rect 19234 36318 19236 36370
rect 18508 33954 18564 33964
rect 19068 32004 19124 32014
rect 19068 30100 19124 31948
rect 19068 30034 19124 30044
rect 19180 26908 19236 36318
rect 19516 36370 19572 39200
rect 19852 36372 19908 36382
rect 19516 36318 19518 36370
rect 19570 36318 19572 36370
rect 19516 36306 19572 36318
rect 19740 36370 19908 36372
rect 19740 36318 19854 36370
rect 19906 36318 19908 36370
rect 19740 36316 19908 36318
rect 19292 34020 19348 34030
rect 19348 33964 19684 34020
rect 19292 33954 19348 33964
rect 19180 26852 19572 26908
rect 19292 25508 19348 25518
rect 18956 25452 19292 25508
rect 18060 25396 18116 25406
rect 18060 25394 18340 25396
rect 18060 25342 18062 25394
rect 18114 25342 18340 25394
rect 18060 25340 18340 25342
rect 18060 25330 18116 25340
rect 17948 24722 18004 24734
rect 17948 24670 17950 24722
rect 18002 24670 18004 24722
rect 17948 24162 18004 24670
rect 17948 24110 17950 24162
rect 18002 24110 18004 24162
rect 17948 24098 18004 24110
rect 18284 24162 18340 25340
rect 18956 24946 19012 25452
rect 19292 25442 19348 25452
rect 19180 25284 19236 25294
rect 19404 25284 19460 25294
rect 19180 25190 19236 25228
rect 19292 25228 19404 25284
rect 18956 24894 18958 24946
rect 19010 24894 19012 24946
rect 18956 24882 19012 24894
rect 18396 24836 18452 24846
rect 18396 24722 18452 24780
rect 18396 24670 18398 24722
rect 18450 24670 18452 24722
rect 18396 24658 18452 24670
rect 19292 24722 19348 25228
rect 19404 25218 19460 25228
rect 19516 25172 19572 26852
rect 19628 25394 19684 33964
rect 19740 32004 19796 36316
rect 19852 36306 19908 36316
rect 20188 36370 20244 39200
rect 20188 36318 20190 36370
rect 20242 36318 20244 36370
rect 20188 36306 20244 36318
rect 20860 36372 20916 39200
rect 21308 36484 21364 36494
rect 21196 36482 21364 36484
rect 21196 36430 21310 36482
rect 21362 36430 21364 36482
rect 21196 36428 21364 36430
rect 21084 36372 21140 36382
rect 20860 36370 21140 36372
rect 20860 36318 21086 36370
rect 21138 36318 21140 36370
rect 20860 36316 21140 36318
rect 21084 36306 21140 36316
rect 19860 36092 20124 36102
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 19860 36026 20124 36036
rect 19860 34524 20124 34534
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 19860 34458 20124 34468
rect 19860 32956 20124 32966
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 19860 32890 20124 32900
rect 21196 31948 21252 36428
rect 21308 36418 21364 36428
rect 21532 36484 21588 39200
rect 21756 36484 21812 36494
rect 21532 36482 21812 36484
rect 21532 36430 21758 36482
rect 21810 36430 21812 36482
rect 21532 36428 21812 36430
rect 21532 35922 21588 36428
rect 21756 36418 21812 36428
rect 22204 36372 22260 39200
rect 22428 36372 22484 36382
rect 22204 36370 22484 36372
rect 22204 36318 22430 36370
rect 22482 36318 22484 36370
rect 22204 36316 22484 36318
rect 22428 36306 22484 36316
rect 22764 36370 22820 36382
rect 22764 36318 22766 36370
rect 22818 36318 22820 36370
rect 21532 35870 21534 35922
rect 21586 35870 21588 35922
rect 21532 35858 21588 35870
rect 22092 36258 22148 36270
rect 22092 36206 22094 36258
rect 22146 36206 22148 36258
rect 19740 31938 19796 31948
rect 20860 31892 21252 31948
rect 22092 31948 22148 36206
rect 22092 31892 22260 31948
rect 19860 31388 20124 31398
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 19860 31322 20124 31332
rect 20188 30100 20244 30110
rect 19860 29820 20124 29830
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 19860 29754 20124 29764
rect 19860 28252 20124 28262
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 19860 28186 20124 28196
rect 19860 26684 20124 26694
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 19860 26618 20124 26628
rect 19852 25508 19908 25518
rect 19852 25414 19908 25452
rect 19628 25342 19630 25394
rect 19682 25342 19684 25394
rect 19628 25330 19684 25342
rect 19740 25284 19796 25294
rect 19516 25116 19684 25172
rect 19292 24670 19294 24722
rect 19346 24670 19348 24722
rect 19292 24658 19348 24670
rect 18284 24110 18286 24162
rect 18338 24110 18340 24162
rect 18284 24098 18340 24110
rect 18620 24500 18676 24510
rect 19516 24500 19572 24510
rect 18620 24162 18676 24444
rect 18620 24110 18622 24162
rect 18674 24110 18676 24162
rect 18620 24098 18676 24110
rect 19404 24444 19516 24500
rect 18844 23940 18900 23950
rect 18844 23846 18900 23884
rect 19292 23828 19348 23838
rect 19404 23828 19460 24444
rect 19516 24406 19572 24444
rect 19292 23826 19460 23828
rect 19292 23774 19294 23826
rect 19346 23774 19460 23826
rect 19292 23772 19460 23774
rect 19516 23938 19572 23950
rect 19516 23886 19518 23938
rect 19570 23886 19572 23938
rect 19292 23762 19348 23772
rect 18060 23156 18116 23166
rect 19404 23156 19460 23166
rect 18060 23154 18340 23156
rect 18060 23102 18062 23154
rect 18114 23102 18340 23154
rect 18060 23100 18340 23102
rect 18060 23090 18116 23100
rect 18284 22594 18340 23100
rect 18284 22542 18286 22594
rect 18338 22542 18340 22594
rect 18284 22530 18340 22542
rect 19292 23154 19460 23156
rect 19292 23102 19406 23154
rect 19458 23102 19460 23154
rect 19292 23100 19460 23102
rect 19292 22594 19348 23100
rect 19404 23090 19460 23100
rect 19292 22542 19294 22594
rect 19346 22542 19348 22594
rect 19292 22530 19348 22542
rect 18844 22484 18900 22494
rect 18844 22390 18900 22428
rect 18620 22372 18676 22382
rect 18676 22316 18788 22372
rect 18620 22278 18676 22316
rect 17724 21810 17892 21812
rect 17724 21758 17726 21810
rect 17778 21758 17892 21810
rect 17724 21756 17892 21758
rect 17948 22146 18004 22158
rect 17948 22094 17950 22146
rect 18002 22094 18004 22146
rect 15372 21746 15428 21756
rect 17724 21746 17780 21756
rect 12348 21700 12404 21710
rect 12348 21606 12404 21644
rect 12572 21588 12628 21598
rect 14924 21588 14980 21598
rect 12460 21586 12628 21588
rect 12460 21534 12574 21586
rect 12626 21534 12628 21586
rect 12460 21532 12628 21534
rect 10332 21364 10388 21374
rect 5874 21196 6138 21206
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 5874 21130 6138 21140
rect 10332 20580 10388 21308
rect 12348 21028 12404 21038
rect 12460 21028 12516 21532
rect 12572 21522 12628 21532
rect 14812 21586 14980 21588
rect 14812 21534 14926 21586
rect 14978 21534 14980 21586
rect 14812 21532 14980 21534
rect 12348 21026 12516 21028
rect 12348 20974 12350 21026
rect 12402 20974 12516 21026
rect 12348 20972 12516 20974
rect 14700 21028 14756 21038
rect 14812 21028 14868 21532
rect 14924 21522 14980 21532
rect 15596 21586 15652 21598
rect 15596 21534 15598 21586
rect 15650 21534 15652 21586
rect 15198 21196 15462 21206
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15198 21130 15462 21140
rect 14700 21026 14868 21028
rect 14700 20974 14702 21026
rect 14754 20974 14868 21026
rect 14700 20972 14868 20974
rect 12348 20962 12404 20972
rect 14700 20962 14756 20972
rect 11788 20802 11844 20814
rect 12012 20804 12068 20814
rect 11788 20750 11790 20802
rect 11842 20750 11844 20802
rect 11116 20692 11172 20702
rect 10780 20580 10836 20618
rect 11116 20598 11172 20636
rect 11452 20690 11508 20702
rect 11452 20638 11454 20690
rect 11506 20638 11508 20690
rect 10332 20524 10780 20580
rect 5874 19628 6138 19638
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 5874 19562 6138 19572
rect 2828 19170 2884 19180
rect 1708 19012 1764 19022
rect 1708 18918 1764 18956
rect 1708 18562 1764 18574
rect 1708 18510 1710 18562
rect 1762 18510 1764 18562
rect 1708 18228 1764 18510
rect 2044 18452 2100 18462
rect 10332 18452 10388 20524
rect 10780 20514 10836 20524
rect 10536 20412 10800 20422
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10536 20346 10800 20356
rect 11452 20244 11508 20638
rect 11788 20580 11844 20750
rect 11788 20514 11844 20524
rect 11900 20802 12068 20804
rect 11900 20750 12014 20802
rect 12066 20750 12068 20802
rect 11900 20748 12068 20750
rect 11564 20244 11620 20254
rect 11452 20242 11620 20244
rect 11452 20190 11566 20242
rect 11618 20190 11620 20242
rect 11452 20188 11620 20190
rect 11564 20178 11620 20188
rect 11788 20244 11844 20254
rect 10780 20132 10836 20142
rect 10780 20038 10836 20076
rect 11676 20132 11732 20142
rect 11228 19908 11284 19918
rect 11116 19906 11284 19908
rect 11116 19854 11230 19906
rect 11282 19854 11284 19906
rect 11116 19852 11284 19854
rect 10536 18844 10800 18854
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10536 18778 10800 18788
rect 10892 18562 10948 18574
rect 10892 18510 10894 18562
rect 10946 18510 10948 18562
rect 10556 18452 10612 18462
rect 10332 18450 10612 18452
rect 10332 18398 10558 18450
rect 10610 18398 10612 18450
rect 10332 18396 10612 18398
rect 2044 18358 2100 18396
rect 10556 18386 10612 18396
rect 1708 18162 1764 18172
rect 5874 18060 6138 18070
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 5874 17994 6138 18004
rect 2044 17892 2100 17902
rect 1932 17836 2044 17892
rect 1708 17556 1764 17566
rect 1708 17462 1764 17500
rect 1708 16994 1764 17006
rect 1708 16942 1710 16994
rect 1762 16942 1764 16994
rect 1708 16212 1764 16942
rect 1708 16146 1764 16156
rect 1932 16098 1988 17836
rect 2044 17826 2100 17836
rect 2716 17668 2772 17678
rect 2716 17574 2772 17612
rect 10892 17668 10948 18510
rect 10892 17602 10948 17612
rect 3164 17556 3220 17566
rect 3164 17462 3220 17500
rect 2044 17444 2100 17454
rect 2044 17350 2100 17388
rect 2380 17442 2436 17454
rect 2380 17390 2382 17442
rect 2434 17390 2436 17442
rect 2380 17108 2436 17390
rect 11116 17444 11172 19852
rect 11228 19842 11284 19852
rect 11564 19348 11620 19358
rect 11676 19348 11732 20076
rect 11564 19346 11676 19348
rect 11564 19294 11566 19346
rect 11618 19294 11676 19346
rect 11564 19292 11676 19294
rect 11564 19282 11620 19292
rect 11676 19254 11732 19292
rect 11788 19124 11844 20188
rect 11900 19796 11956 20748
rect 12012 20738 12068 20748
rect 13916 20802 13972 20814
rect 13916 20750 13918 20802
rect 13970 20750 13972 20802
rect 11900 19702 11956 19740
rect 12012 20580 12068 20590
rect 11900 19124 11956 19134
rect 11788 19122 11956 19124
rect 11788 19070 11902 19122
rect 11954 19070 11956 19122
rect 11788 19068 11956 19070
rect 11900 19058 11956 19068
rect 11228 18452 11284 18462
rect 11564 18452 11620 18462
rect 11228 18450 11620 18452
rect 11228 18398 11230 18450
rect 11282 18398 11566 18450
rect 11618 18398 11620 18450
rect 11228 18396 11620 18398
rect 12012 18452 12068 20524
rect 13580 20580 13636 20590
rect 13916 20580 13972 20750
rect 14700 20804 14756 20814
rect 13636 20524 13972 20580
rect 14140 20692 14196 20702
rect 13580 20486 13636 20524
rect 12124 20132 12180 20142
rect 12124 20018 12180 20076
rect 14140 20130 14196 20636
rect 14140 20078 14142 20130
rect 14194 20078 14196 20130
rect 14140 20066 14196 20078
rect 14252 20690 14308 20702
rect 14252 20638 14254 20690
rect 14306 20638 14308 20690
rect 14252 20132 14308 20638
rect 14252 20038 14308 20076
rect 14700 20130 14756 20748
rect 15596 20804 15652 21534
rect 17948 21586 18004 22094
rect 18732 21812 18788 22316
rect 18844 21812 18900 21822
rect 18732 21810 19460 21812
rect 18732 21758 18846 21810
rect 18898 21758 19460 21810
rect 18732 21756 19460 21758
rect 18844 21746 18900 21756
rect 17948 21534 17950 21586
rect 18002 21534 18004 21586
rect 17948 21522 18004 21534
rect 18508 21586 18564 21598
rect 18508 21534 18510 21586
rect 18562 21534 18564 21586
rect 16828 21028 16884 21038
rect 15820 20916 15876 20926
rect 15820 20914 16548 20916
rect 15820 20862 15822 20914
rect 15874 20862 16548 20914
rect 15820 20860 16548 20862
rect 15820 20850 15876 20860
rect 15596 20738 15652 20748
rect 14700 20078 14702 20130
rect 14754 20078 14756 20130
rect 14700 20066 14756 20078
rect 15260 20692 15316 20702
rect 15260 20130 15316 20636
rect 16268 20692 16324 20702
rect 16268 20598 16324 20636
rect 16380 20690 16436 20702
rect 16380 20638 16382 20690
rect 16434 20638 16436 20690
rect 16380 20356 16436 20638
rect 16156 20300 16436 20356
rect 16492 20690 16548 20860
rect 16492 20638 16494 20690
rect 16546 20638 16548 20690
rect 15260 20078 15262 20130
rect 15314 20078 15316 20130
rect 15260 20066 15316 20078
rect 15372 20244 15428 20254
rect 15372 20130 15428 20188
rect 16156 20244 16212 20300
rect 16492 20244 16548 20638
rect 16828 20580 16884 20972
rect 17948 20916 18004 20926
rect 16940 20804 16996 20814
rect 17500 20804 17556 20814
rect 16940 20802 17556 20804
rect 16940 20750 16942 20802
rect 16994 20750 17502 20802
rect 17554 20750 17556 20802
rect 16940 20748 17556 20750
rect 16940 20738 16996 20748
rect 17500 20738 17556 20748
rect 17948 20690 18004 20860
rect 18172 20804 18228 20814
rect 17948 20638 17950 20690
rect 18002 20638 18004 20690
rect 17948 20626 18004 20638
rect 18060 20802 18228 20804
rect 18060 20750 18174 20802
rect 18226 20750 18228 20802
rect 18060 20748 18228 20750
rect 17276 20580 17332 20590
rect 16828 20578 17332 20580
rect 16828 20526 17278 20578
rect 17330 20526 17332 20578
rect 16828 20524 17332 20526
rect 17276 20514 17332 20524
rect 16156 20150 16212 20188
rect 16380 20188 16548 20244
rect 17948 20244 18004 20254
rect 18060 20244 18116 20748
rect 18172 20738 18228 20748
rect 18508 20468 18564 21534
rect 19180 21588 19236 21598
rect 19180 21494 19236 21532
rect 19404 21586 19460 21756
rect 19404 21534 19406 21586
rect 19458 21534 19460 21586
rect 19404 21522 19460 21534
rect 19068 20802 19124 20814
rect 19068 20750 19070 20802
rect 19122 20750 19124 20802
rect 18844 20692 18900 20702
rect 18844 20598 18900 20636
rect 18396 20412 18564 20468
rect 19068 20580 19124 20750
rect 18396 20244 18452 20412
rect 17948 20242 18116 20244
rect 17948 20190 17950 20242
rect 18002 20190 18116 20242
rect 17948 20188 18116 20190
rect 18284 20188 18452 20244
rect 18508 20244 18564 20254
rect 19068 20244 19124 20524
rect 19516 20356 19572 23886
rect 19628 22596 19684 25116
rect 19740 24948 19796 25228
rect 19860 25116 20124 25126
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 19860 25050 20124 25060
rect 19740 24892 20132 24948
rect 19852 24724 19908 24734
rect 19852 24630 19908 24668
rect 20076 24050 20132 24892
rect 20188 24946 20244 30044
rect 20188 24894 20190 24946
rect 20242 24894 20244 24946
rect 20188 24882 20244 24894
rect 20076 23998 20078 24050
rect 20130 23998 20132 24050
rect 20076 23716 20132 23998
rect 20300 24836 20356 24846
rect 20076 23660 20244 23716
rect 19860 23548 20124 23558
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 19860 23482 20124 23492
rect 20188 23380 20244 23660
rect 19964 23324 20244 23380
rect 19740 23268 19796 23278
rect 19740 23174 19796 23212
rect 19964 22596 20020 23324
rect 19628 22540 19796 22596
rect 19628 22372 19684 22382
rect 19628 22278 19684 22316
rect 19740 21812 19796 22540
rect 19852 22484 19908 22494
rect 19964 22484 20020 22540
rect 19852 22482 20020 22484
rect 19852 22430 19854 22482
rect 19906 22430 20020 22482
rect 19852 22428 20020 22430
rect 20188 23154 20244 23166
rect 20188 23102 20190 23154
rect 20242 23102 20244 23154
rect 19852 22418 19908 22428
rect 19860 21980 20124 21990
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 19860 21914 20124 21924
rect 20076 21812 20132 21822
rect 19740 21810 20132 21812
rect 19740 21758 20078 21810
rect 20130 21758 20132 21810
rect 19740 21756 20132 21758
rect 20076 21746 20132 21756
rect 19740 21476 19796 21486
rect 19740 21382 19796 21420
rect 20188 20804 20244 23102
rect 20300 22820 20356 24780
rect 20524 24724 20580 24734
rect 20524 24630 20580 24668
rect 20636 23940 20692 23950
rect 20636 23604 20692 23884
rect 20412 23266 20468 23278
rect 20412 23214 20414 23266
rect 20466 23214 20468 23266
rect 20412 23156 20468 23214
rect 20412 23090 20468 23100
rect 20300 22764 20468 22820
rect 20300 22596 20356 22606
rect 20300 22482 20356 22540
rect 20300 22430 20302 22482
rect 20354 22430 20356 22482
rect 20300 22260 20356 22430
rect 20300 22194 20356 22204
rect 20300 21586 20356 21598
rect 20300 21534 20302 21586
rect 20354 21534 20356 21586
rect 20300 21476 20356 21534
rect 20412 21588 20468 22764
rect 20636 22484 20692 23548
rect 20860 23380 20916 31892
rect 21420 26516 21476 26526
rect 21420 25506 21476 26460
rect 21420 25454 21422 25506
rect 21474 25454 21476 25506
rect 21420 25284 21476 25454
rect 22092 25508 22148 25518
rect 22092 25414 22148 25452
rect 21420 25218 21476 25228
rect 21532 25394 21588 25406
rect 21532 25342 21534 25394
rect 21586 25342 21588 25394
rect 21532 25060 21588 25342
rect 21196 25004 21588 25060
rect 21644 25394 21700 25406
rect 21644 25342 21646 25394
rect 21698 25342 21700 25394
rect 21084 24836 21140 24846
rect 21084 24742 21140 24780
rect 20860 23314 20916 23324
rect 21196 24722 21252 25004
rect 21644 24948 21700 25342
rect 21308 24892 21700 24948
rect 21308 24834 21364 24892
rect 21308 24782 21310 24834
rect 21362 24782 21364 24834
rect 21308 24770 21364 24782
rect 21196 24670 21198 24722
rect 21250 24670 21252 24722
rect 21084 23268 21140 23278
rect 21084 23174 21140 23212
rect 20860 23154 20916 23166
rect 20860 23102 20862 23154
rect 20914 23102 20916 23154
rect 20860 22596 20916 23102
rect 21196 23156 21252 24670
rect 21644 24052 21700 24892
rect 21756 25396 21812 25406
rect 21756 24946 21812 25340
rect 21756 24894 21758 24946
rect 21810 24894 21812 24946
rect 21756 24882 21812 24894
rect 22204 24946 22260 31892
rect 22316 26516 22372 26526
rect 22316 26422 22372 26460
rect 22428 25396 22484 25406
rect 22428 25302 22484 25340
rect 22764 25394 22820 36318
rect 22876 36372 22932 39200
rect 23548 37828 23604 39200
rect 23548 37772 24164 37828
rect 24108 36484 24164 37772
rect 24220 36708 24276 39200
rect 24522 36876 24786 36886
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24522 36810 24786 36820
rect 24220 36642 24276 36652
rect 24780 36484 24836 36494
rect 24108 36428 24612 36484
rect 23100 36372 23156 36382
rect 22876 36370 23156 36372
rect 22876 36318 23102 36370
rect 23154 36318 23156 36370
rect 22876 36316 23156 36318
rect 23100 36306 23156 36316
rect 23324 36372 23380 36382
rect 23100 25508 23156 25518
rect 23100 25414 23156 25452
rect 22764 25342 22766 25394
rect 22818 25342 22820 25394
rect 22764 25330 22820 25342
rect 22204 24894 22206 24946
rect 22258 24894 22260 24946
rect 22204 24836 22260 24894
rect 23324 24948 23380 36316
rect 23436 36370 23492 36382
rect 23436 36318 23438 36370
rect 23490 36318 23492 36370
rect 23436 25394 23492 36318
rect 24556 36370 24612 36428
rect 24556 36318 24558 36370
rect 24610 36318 24612 36370
rect 24556 36306 24612 36318
rect 24668 36482 24836 36484
rect 24668 36430 24782 36482
rect 24834 36430 24836 36482
rect 24668 36428 24836 36430
rect 24668 35476 24724 36428
rect 24780 36418 24836 36428
rect 24892 36484 24948 39200
rect 37548 36932 37604 36942
rect 33846 36876 34110 36886
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 33846 36810 34110 36820
rect 24892 36418 24948 36428
rect 25228 36708 25284 36718
rect 25228 36370 25284 36652
rect 25676 36484 25732 36494
rect 25228 36318 25230 36370
rect 25282 36318 25284 36370
rect 25228 36306 25284 36318
rect 25564 36372 25620 36382
rect 25564 36278 25620 36316
rect 25676 35922 25732 36428
rect 26124 36484 26180 36494
rect 26124 36390 26180 36428
rect 35532 36484 35588 36494
rect 37548 36484 37604 36876
rect 35532 36482 36484 36484
rect 35532 36430 35534 36482
rect 35586 36430 36484 36482
rect 35532 36428 36484 36430
rect 35532 36418 35588 36428
rect 36428 36372 36484 36428
rect 37548 36482 37716 36484
rect 37548 36430 37550 36482
rect 37602 36430 37716 36482
rect 37548 36428 37716 36430
rect 37548 36418 37604 36428
rect 36540 36372 36596 36382
rect 36428 36370 36596 36372
rect 36428 36318 36542 36370
rect 36594 36318 36596 36370
rect 36428 36316 36596 36318
rect 25676 35870 25678 35922
rect 25730 35870 25732 35922
rect 25676 35858 25732 35870
rect 25900 36258 25956 36270
rect 25900 36206 25902 36258
rect 25954 36206 25956 36258
rect 24108 35420 24724 35476
rect 23436 25342 23438 25394
rect 23490 25342 23492 25394
rect 23436 25330 23492 25342
rect 23996 31556 24052 31566
rect 23436 24948 23492 24958
rect 23324 24946 23492 24948
rect 23324 24894 23438 24946
rect 23490 24894 23492 24946
rect 23324 24892 23492 24894
rect 23436 24882 23492 24892
rect 22204 24770 22260 24780
rect 23100 24724 23156 24734
rect 22540 24722 23156 24724
rect 22540 24670 23102 24722
rect 23154 24670 23156 24722
rect 22540 24668 23156 24670
rect 22540 24162 22596 24668
rect 23100 24658 23156 24668
rect 23772 24722 23828 24734
rect 23772 24670 23774 24722
rect 23826 24670 23828 24722
rect 22764 24164 22820 24174
rect 22540 24110 22542 24162
rect 22594 24110 22596 24162
rect 22540 24098 22596 24110
rect 22652 24108 22764 24164
rect 21644 23996 22148 24052
rect 22092 23938 22148 23996
rect 22092 23886 22094 23938
rect 22146 23886 22148 23938
rect 21868 23828 21924 23838
rect 21756 23826 21924 23828
rect 21756 23774 21870 23826
rect 21922 23774 21924 23826
rect 21756 23772 21924 23774
rect 21196 23090 21252 23100
rect 21420 23716 21476 23726
rect 21756 23716 21812 23772
rect 21868 23762 21924 23772
rect 21980 23826 22036 23838
rect 21980 23774 21982 23826
rect 22034 23774 22036 23826
rect 21420 23714 21812 23716
rect 21420 23662 21422 23714
rect 21474 23662 21812 23714
rect 21420 23660 21812 23662
rect 20860 22540 21140 22596
rect 20748 22484 20804 22494
rect 20636 22482 21028 22484
rect 20636 22430 20750 22482
rect 20802 22430 21028 22482
rect 20636 22428 21028 22430
rect 20748 22418 20804 22428
rect 20972 21810 21028 22428
rect 20972 21758 20974 21810
rect 21026 21758 21028 21810
rect 20972 21746 21028 21758
rect 20468 21532 20580 21588
rect 20412 21522 20468 21532
rect 20300 21410 20356 21420
rect 19964 20748 20188 20804
rect 19964 20690 20020 20748
rect 20188 20710 20244 20748
rect 20412 20692 20468 20702
rect 19964 20638 19966 20690
rect 20018 20638 20020 20690
rect 19964 20626 20020 20638
rect 20300 20690 20468 20692
rect 20300 20638 20414 20690
rect 20466 20638 20468 20690
rect 20300 20636 20468 20638
rect 19628 20580 19684 20590
rect 19628 20486 19684 20524
rect 18508 20242 19124 20244
rect 18508 20190 18510 20242
rect 18562 20190 19124 20242
rect 18508 20188 19124 20190
rect 19180 20300 19572 20356
rect 19860 20412 20124 20422
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 19860 20346 20124 20356
rect 15372 20078 15374 20130
rect 15426 20078 15428 20130
rect 15372 20066 15428 20078
rect 12124 19966 12126 20018
rect 12178 19966 12180 20018
rect 12124 19954 12180 19966
rect 14028 20018 14084 20030
rect 14028 19966 14030 20018
rect 14082 19966 14084 20018
rect 13020 19908 13076 19918
rect 13580 19908 13636 19918
rect 12908 19906 13580 19908
rect 12908 19854 13022 19906
rect 13074 19854 13580 19906
rect 12908 19852 13580 19854
rect 12460 19796 12516 19806
rect 12236 19794 12516 19796
rect 12236 19742 12462 19794
rect 12514 19742 12516 19794
rect 12236 19740 12516 19742
rect 12236 19234 12292 19740
rect 12460 19730 12516 19740
rect 12796 19796 12852 19806
rect 12796 19702 12852 19740
rect 12796 19236 12852 19246
rect 12236 19182 12238 19234
rect 12290 19182 12292 19234
rect 12236 19170 12292 19182
rect 12460 19234 12852 19236
rect 12460 19182 12798 19234
rect 12850 19182 12852 19234
rect 12460 19180 12852 19182
rect 12460 18674 12516 19180
rect 12796 19170 12852 19180
rect 12460 18622 12462 18674
rect 12514 18622 12516 18674
rect 12460 18610 12516 18622
rect 12572 19010 12628 19022
rect 12572 18958 12574 19010
rect 12626 18958 12628 19010
rect 12124 18452 12180 18462
rect 12012 18396 12124 18452
rect 11228 18386 11284 18396
rect 11564 18386 11620 18396
rect 12124 18358 12180 18396
rect 11900 18228 11956 18238
rect 11900 17890 11956 18172
rect 11900 17838 11902 17890
rect 11954 17838 11956 17890
rect 11900 17826 11956 17838
rect 12572 17892 12628 18958
rect 12796 18228 12852 18238
rect 12908 18228 12964 19852
rect 13020 19842 13076 19852
rect 13580 19814 13636 19852
rect 13580 19348 13636 19358
rect 14028 19348 14084 19966
rect 15036 20018 15092 20030
rect 15036 19966 15038 20018
rect 15090 19966 15092 20018
rect 14924 19908 14980 19918
rect 15036 19908 15092 19966
rect 15820 20020 15876 20030
rect 15876 19964 15988 20020
rect 15820 19954 15876 19964
rect 14980 19852 15092 19908
rect 14924 19842 14980 19852
rect 15820 19796 15876 19806
rect 15596 19794 15876 19796
rect 15596 19742 15822 19794
rect 15874 19742 15876 19794
rect 15596 19740 15876 19742
rect 15198 19628 15462 19638
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15198 19562 15462 19572
rect 13468 19292 13580 19348
rect 13468 18676 13524 19292
rect 13580 19254 13636 19292
rect 13916 19292 14028 19348
rect 13020 18674 13524 18676
rect 13020 18622 13470 18674
rect 13522 18622 13524 18674
rect 13020 18620 13524 18622
rect 13020 18450 13076 18620
rect 13468 18610 13524 18620
rect 13916 18562 13972 19292
rect 14028 19282 14084 19292
rect 14924 19236 14980 19246
rect 13916 18510 13918 18562
rect 13970 18510 13972 18562
rect 13916 18498 13972 18510
rect 14588 19124 14644 19134
rect 13020 18398 13022 18450
rect 13074 18398 13076 18450
rect 13020 18386 13076 18398
rect 13804 18452 13860 18462
rect 12908 18172 13076 18228
rect 12796 18134 12852 18172
rect 12572 17826 12628 17836
rect 11676 17666 11732 17678
rect 11676 17614 11678 17666
rect 11730 17614 11732 17666
rect 11340 17444 11396 17454
rect 11676 17444 11732 17614
rect 12908 17556 12964 17566
rect 12908 17462 12964 17500
rect 11116 17442 11732 17444
rect 11116 17390 11342 17442
rect 11394 17390 11732 17442
rect 11116 17388 11732 17390
rect 12236 17442 12292 17454
rect 12236 17390 12238 17442
rect 12290 17390 12292 17442
rect 10536 17276 10800 17286
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10536 17210 10800 17220
rect 2380 17042 2436 17052
rect 2268 16996 2324 17006
rect 2044 16884 2100 16894
rect 2044 16790 2100 16828
rect 1932 16046 1934 16098
rect 1986 16046 1988 16098
rect 1932 16034 1988 16046
rect 1708 15876 1764 15886
rect 1708 15782 1764 15820
rect 1708 15426 1764 15438
rect 1708 15374 1710 15426
rect 1762 15374 1764 15426
rect 1708 14868 1764 15374
rect 2044 15316 2100 15326
rect 2044 15222 2100 15260
rect 1708 14802 1764 14812
rect 2156 15204 2212 15214
rect 1708 14418 1764 14430
rect 1708 14366 1710 14418
rect 1762 14366 1764 14418
rect 1708 14196 1764 14366
rect 2044 14308 2100 14318
rect 2044 14214 2100 14252
rect 1708 14130 1764 14140
rect 2044 13972 2100 13982
rect 2156 13972 2212 15148
rect 2044 13970 2212 13972
rect 2044 13918 2046 13970
rect 2098 13918 2212 13970
rect 2044 13916 2212 13918
rect 2044 13906 2100 13916
rect 1708 13746 1764 13758
rect 1708 13694 1710 13746
rect 1762 13694 1764 13746
rect 1708 13524 1764 13694
rect 1708 13458 1764 13468
rect 1708 12852 1764 12862
rect 1708 12758 1764 12796
rect 2044 12852 2100 12862
rect 2268 12852 2324 16940
rect 11340 16996 11396 17388
rect 11340 16930 11396 16940
rect 12124 16994 12180 17006
rect 12124 16942 12126 16994
rect 12178 16942 12180 16994
rect 5874 16492 6138 16502
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 5874 16426 6138 16436
rect 10536 15708 10800 15718
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10536 15642 10800 15652
rect 12124 15316 12180 16942
rect 12236 16884 12292 17390
rect 12572 17442 12628 17454
rect 12572 17390 12574 17442
rect 12626 17390 12628 17442
rect 12348 16884 12404 16894
rect 12236 16882 12404 16884
rect 12236 16830 12350 16882
rect 12402 16830 12404 16882
rect 12236 16828 12404 16830
rect 12348 16818 12404 16828
rect 12572 16884 12628 17390
rect 12908 16996 12964 17006
rect 13020 16996 13076 18172
rect 13804 17780 13860 18396
rect 13468 17724 13860 17780
rect 13468 17106 13524 17724
rect 13804 17666 13860 17724
rect 13804 17614 13806 17666
rect 13858 17614 13860 17666
rect 13804 17602 13860 17614
rect 14028 18452 14084 18462
rect 14028 17666 14084 18396
rect 14028 17614 14030 17666
rect 14082 17614 14084 17666
rect 13468 17054 13470 17106
rect 13522 17054 13524 17106
rect 13468 17042 13524 17054
rect 13692 17556 13748 17566
rect 13692 17106 13748 17500
rect 13692 17054 13694 17106
rect 13746 17054 13748 17106
rect 13692 17042 13748 17054
rect 12964 16940 13076 16996
rect 12908 16902 12964 16940
rect 12572 16818 12628 16828
rect 14028 16772 14084 17614
rect 14140 18450 14196 18462
rect 14140 18398 14142 18450
rect 14194 18398 14196 18450
rect 14140 17892 14196 18398
rect 14588 18450 14644 19068
rect 14924 19122 14980 19180
rect 15260 19236 15316 19246
rect 15596 19236 15652 19740
rect 15820 19730 15876 19740
rect 15932 19348 15988 19964
rect 15260 19234 15652 19236
rect 15260 19182 15262 19234
rect 15314 19182 15652 19234
rect 15260 19180 15652 19182
rect 15708 19292 15988 19348
rect 15260 19170 15316 19180
rect 14924 19070 14926 19122
rect 14978 19070 14980 19122
rect 14924 19058 14980 19070
rect 15596 19012 15652 19022
rect 15708 19012 15764 19292
rect 15932 19124 15988 19134
rect 15932 19030 15988 19068
rect 15596 19010 15764 19012
rect 15596 18958 15598 19010
rect 15650 18958 15764 19010
rect 15596 18956 15764 18958
rect 15596 18946 15652 18956
rect 14588 18398 14590 18450
rect 14642 18398 14644 18450
rect 14588 18386 14644 18398
rect 15372 18562 15428 18574
rect 15372 18510 15374 18562
rect 15426 18510 15428 18562
rect 15372 18452 15428 18510
rect 15820 18564 15876 18574
rect 15372 18386 15428 18396
rect 15708 18452 15764 18462
rect 15820 18452 15876 18508
rect 15708 18450 15876 18452
rect 15708 18398 15710 18450
rect 15762 18398 15876 18450
rect 15708 18396 15876 18398
rect 15708 18386 15764 18396
rect 14140 17666 14196 17836
rect 14924 18340 14980 18350
rect 14140 17614 14142 17666
rect 14194 17614 14196 17666
rect 14140 16994 14196 17614
rect 14588 17668 14644 17678
rect 14588 17574 14644 17612
rect 14924 17554 14980 18284
rect 14924 17502 14926 17554
rect 14978 17502 14980 17554
rect 14924 17490 14980 17502
rect 15036 18338 15092 18350
rect 15036 18286 15038 18338
rect 15090 18286 15092 18338
rect 15036 17444 15092 18286
rect 15198 18060 15462 18070
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15198 17994 15462 18004
rect 15148 17668 15204 17678
rect 15148 17574 15204 17612
rect 15036 17378 15092 17388
rect 15596 17554 15652 17566
rect 15596 17502 15598 17554
rect 15650 17502 15652 17554
rect 14140 16942 14142 16994
rect 14194 16942 14196 16994
rect 14140 16930 14196 16942
rect 14364 16996 14420 17006
rect 14364 16902 14420 16940
rect 14252 16882 14308 16894
rect 14252 16830 14254 16882
rect 14306 16830 14308 16882
rect 14252 16772 14308 16830
rect 14028 16716 14308 16772
rect 15372 16770 15428 16782
rect 15372 16718 15374 16770
rect 15426 16718 15428 16770
rect 15372 16660 15428 16718
rect 15036 16604 15428 16660
rect 15596 16658 15652 17502
rect 15596 16606 15598 16658
rect 15650 16606 15652 16658
rect 15036 16324 15092 16604
rect 15198 16492 15462 16502
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15198 16426 15462 16436
rect 15036 16268 15204 16324
rect 14252 15988 14308 15998
rect 12124 15250 12180 15260
rect 14028 15316 14084 15326
rect 14252 15316 14308 15932
rect 14028 15314 14308 15316
rect 14028 15262 14030 15314
rect 14082 15262 14308 15314
rect 14028 15260 14308 15262
rect 14028 15250 14084 15260
rect 5874 14924 6138 14934
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 5874 14858 6138 14868
rect 14252 14530 14308 15260
rect 14700 15204 14756 15214
rect 14700 15110 14756 15148
rect 15148 15092 15204 16268
rect 15596 15204 15652 16606
rect 15596 15138 15652 15148
rect 14252 14478 14254 14530
rect 14306 14478 14308 14530
rect 14252 14466 14308 14478
rect 15036 15036 15204 15092
rect 14924 14420 14980 14430
rect 15036 14420 15092 15036
rect 15198 14924 15462 14934
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15198 14858 15462 14868
rect 14924 14418 15092 14420
rect 14924 14366 14926 14418
rect 14978 14366 15092 14418
rect 14924 14364 15092 14366
rect 15708 14532 15764 14542
rect 2492 14306 2548 14318
rect 2492 14254 2494 14306
rect 2546 14254 2548 14306
rect 2492 14196 2548 14254
rect 14924 14308 14980 14364
rect 14924 14242 14980 14252
rect 15484 14308 15540 14318
rect 2492 14130 2548 14140
rect 10536 14140 10800 14150
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10536 14074 10800 14084
rect 15484 13858 15540 14252
rect 15484 13806 15486 13858
rect 15538 13806 15540 13858
rect 15484 13794 15540 13806
rect 2492 13634 2548 13646
rect 2492 13582 2494 13634
rect 2546 13582 2548 13634
rect 2492 13524 2548 13582
rect 2492 13458 2548 13468
rect 14812 13636 14868 13646
rect 5874 13356 6138 13366
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 5874 13290 6138 13300
rect 2044 12850 2324 12852
rect 2044 12798 2046 12850
rect 2098 12798 2324 12850
rect 2044 12796 2324 12798
rect 2492 12852 2548 12862
rect 2044 12786 2100 12796
rect 2492 12758 2548 12796
rect 10536 12572 10800 12582
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10536 12506 10800 12516
rect 5874 11788 6138 11798
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 5874 11722 6138 11732
rect 10536 11004 10800 11014
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10536 10938 10800 10948
rect 5874 10220 6138 10230
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 5874 10154 6138 10164
rect 10536 9436 10800 9446
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10536 9370 10800 9380
rect 5874 8652 6138 8662
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 5874 8586 6138 8596
rect 10536 7868 10800 7878
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10536 7802 10800 7812
rect 5874 7084 6138 7094
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 5874 7018 6138 7028
rect 10536 6300 10800 6310
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10536 6234 10800 6244
rect 5874 5516 6138 5526
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 5874 5450 6138 5460
rect 10536 4732 10800 4742
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10536 4666 10800 4676
rect 5874 3948 6138 3958
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 5874 3882 6138 3892
rect 10536 3164 10800 3174
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10536 3098 10800 3108
rect 14812 800 14868 13580
rect 15198 13356 15462 13366
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15198 13290 15462 13300
rect 15198 11788 15462 11798
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15198 11722 15462 11732
rect 15198 10220 15462 10230
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15198 10154 15462 10164
rect 15198 8652 15462 8662
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15198 8586 15462 8596
rect 15198 7084 15462 7094
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15198 7018 15462 7028
rect 15198 5516 15462 5526
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15198 5450 15462 5460
rect 15198 3948 15462 3958
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15198 3882 15462 3892
rect 15484 3554 15540 3566
rect 15484 3502 15486 3554
rect 15538 3502 15540 3554
rect 15484 3220 15540 3502
rect 15708 3442 15764 14476
rect 15820 13970 15876 18396
rect 16044 18452 16100 18462
rect 16044 18358 16100 18396
rect 16268 18450 16324 18462
rect 16268 18398 16270 18450
rect 16322 18398 16324 18450
rect 15932 18340 15988 18350
rect 15932 17554 15988 18284
rect 16268 17892 16324 18398
rect 16268 17826 16324 17836
rect 16380 18452 16436 20188
rect 17948 20178 18004 20188
rect 15932 17502 15934 17554
rect 15986 17502 15988 17554
rect 15932 17490 15988 17502
rect 16380 17444 16436 18396
rect 16492 20018 16548 20030
rect 16492 19966 16494 20018
rect 16546 19966 16548 20018
rect 16492 18340 16548 19966
rect 17388 19906 17444 19918
rect 17388 19854 17390 19906
rect 17442 19854 17444 19906
rect 17164 19236 17220 19246
rect 16828 19234 17220 19236
rect 16828 19182 17166 19234
rect 17218 19182 17220 19234
rect 16828 19180 17220 19182
rect 16828 18674 16884 19180
rect 17164 19170 17220 19180
rect 16940 19012 16996 19022
rect 17388 19012 17444 19854
rect 17612 19796 17668 19806
rect 17612 19702 17668 19740
rect 18172 19796 18228 19806
rect 18172 19122 18228 19740
rect 18172 19070 18174 19122
rect 18226 19070 18228 19122
rect 18172 19058 18228 19070
rect 17724 19012 17780 19022
rect 17388 19010 17780 19012
rect 17388 18958 17726 19010
rect 17778 18958 17780 19010
rect 17388 18956 17780 18958
rect 16940 18918 16996 18956
rect 16828 18622 16830 18674
rect 16882 18622 16884 18674
rect 16828 18610 16884 18622
rect 17500 18452 17556 18462
rect 17612 18452 17668 18956
rect 17724 18946 17780 18956
rect 18172 18562 18228 18574
rect 18172 18510 18174 18562
rect 18226 18510 18228 18562
rect 17556 18396 17668 18452
rect 17836 18452 17892 18462
rect 17500 18386 17556 18396
rect 17836 18358 17892 18396
rect 16492 18274 16548 18284
rect 17724 18340 17780 18350
rect 17724 18246 17780 18284
rect 16828 18228 16884 18238
rect 16828 17892 16884 18172
rect 16380 17378 16436 17388
rect 16492 17890 16884 17892
rect 16492 17838 16830 17890
rect 16882 17838 16884 17890
rect 16492 17836 16884 17838
rect 16492 17106 16548 17836
rect 16828 17826 16884 17836
rect 18172 17892 18228 18510
rect 18172 17826 18228 17836
rect 16604 17666 16660 17678
rect 16604 17614 16606 17666
rect 16658 17614 16660 17666
rect 16604 17444 16660 17614
rect 17164 17668 17220 17678
rect 17724 17668 17780 17678
rect 18284 17668 18340 20188
rect 18508 20178 18564 20188
rect 19180 20130 19236 20300
rect 19180 20078 19182 20130
rect 19234 20078 19236 20130
rect 19180 20066 19236 20078
rect 18396 20020 18452 20030
rect 18396 19906 18452 19964
rect 18396 19854 18398 19906
rect 18450 19854 18452 19906
rect 18396 18564 18452 19854
rect 18956 20018 19012 20030
rect 18956 19966 18958 20018
rect 19010 19966 19012 20018
rect 18956 19348 19012 19966
rect 19516 19684 19572 20300
rect 19964 20132 20020 20142
rect 19964 20038 20020 20076
rect 19628 20020 19684 20030
rect 19628 19926 19684 19964
rect 19516 19618 19572 19628
rect 18508 19346 19012 19348
rect 18508 19294 18958 19346
rect 19010 19294 19012 19346
rect 18508 19292 19012 19294
rect 18508 19234 18564 19292
rect 18956 19282 19012 19292
rect 18508 19182 18510 19234
rect 18562 19182 18564 19234
rect 18508 19170 18564 19182
rect 18396 18498 18452 18508
rect 18844 19122 18900 19134
rect 18844 19070 18846 19122
rect 18898 19070 18900 19122
rect 18508 18452 18564 18462
rect 18508 18358 18564 18396
rect 18844 18450 18900 19070
rect 19740 19124 19796 19134
rect 19068 19010 19124 19022
rect 19068 18958 19070 19010
rect 19122 18958 19124 19010
rect 19068 18564 19124 18958
rect 19180 18676 19236 18686
rect 19740 18676 19796 19068
rect 20076 19012 20132 19022
rect 20076 19010 20244 19012
rect 20076 18958 20078 19010
rect 20130 18958 20244 19010
rect 20076 18956 20244 18958
rect 20076 18946 20132 18956
rect 19860 18844 20124 18854
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 19860 18778 20124 18788
rect 19180 18674 19796 18676
rect 19180 18622 19182 18674
rect 19234 18622 19796 18674
rect 19180 18620 19796 18622
rect 19180 18610 19236 18620
rect 19068 18498 19124 18508
rect 19852 18562 19908 18574
rect 19852 18510 19854 18562
rect 19906 18510 19908 18562
rect 18844 18398 18846 18450
rect 18898 18398 18900 18450
rect 18844 18340 18900 18398
rect 19516 18452 19572 18462
rect 19516 18358 19572 18396
rect 18844 18274 18900 18284
rect 19852 18228 19908 18510
rect 19852 18162 19908 18172
rect 20188 18452 20244 18956
rect 19964 17668 20020 17678
rect 17164 17666 17780 17668
rect 17164 17614 17166 17666
rect 17218 17614 17726 17666
rect 17778 17614 17780 17666
rect 17164 17612 17780 17614
rect 17164 17602 17220 17612
rect 17724 17602 17780 17612
rect 18172 17612 18340 17668
rect 19628 17666 20020 17668
rect 19628 17614 19966 17666
rect 20018 17614 20020 17666
rect 19628 17612 20020 17614
rect 16604 17378 16660 17388
rect 17500 17442 17556 17454
rect 17500 17390 17502 17442
rect 17554 17390 17556 17442
rect 16492 17054 16494 17106
rect 16546 17054 16548 17106
rect 16492 17042 16548 17054
rect 15932 16884 15988 16894
rect 15932 16790 15988 16828
rect 16716 16884 16772 16894
rect 16716 16790 16772 16828
rect 16716 15988 16772 15998
rect 16716 15894 16772 15932
rect 17388 15314 17444 15326
rect 17388 15262 17390 15314
rect 17442 15262 17444 15314
rect 16828 15202 16884 15214
rect 16828 15150 16830 15202
rect 16882 15150 16884 15202
rect 16828 14756 16884 15150
rect 16828 14690 16884 14700
rect 17052 14642 17108 14654
rect 17052 14590 17054 14642
rect 17106 14590 17108 14642
rect 17052 14420 17108 14590
rect 17052 14354 17108 14364
rect 16156 14308 16212 14318
rect 15820 13918 15822 13970
rect 15874 13918 15876 13970
rect 15820 13906 15876 13918
rect 16044 14252 16156 14308
rect 15708 3390 15710 3442
rect 15762 3390 15764 3442
rect 15708 3378 15764 3390
rect 15932 4226 15988 4238
rect 15932 4174 15934 4226
rect 15986 4174 15988 4226
rect 15932 3220 15988 4174
rect 16044 3554 16100 14252
rect 16156 14242 16212 14252
rect 16828 13636 16884 13646
rect 16828 13542 16884 13580
rect 17388 13636 17444 15262
rect 17388 13570 17444 13580
rect 17500 12964 17556 17390
rect 17948 17108 18004 17118
rect 18172 17108 18228 17612
rect 18284 17444 18340 17454
rect 18284 17350 18340 17388
rect 18956 17444 19012 17454
rect 19404 17444 19460 17454
rect 18956 17442 19460 17444
rect 18956 17390 18958 17442
rect 19010 17390 19406 17442
rect 19458 17390 19460 17442
rect 18956 17388 19460 17390
rect 18956 17378 19012 17388
rect 18284 17108 18340 17118
rect 17948 17106 18284 17108
rect 17948 17054 17950 17106
rect 18002 17054 18284 17106
rect 17948 17052 18284 17054
rect 17948 17042 18004 17052
rect 18284 16994 18340 17052
rect 18284 16942 18286 16994
rect 18338 16942 18340 16994
rect 18284 16930 18340 16942
rect 18620 16994 18676 17006
rect 18620 16942 18622 16994
rect 18674 16942 18676 16994
rect 17612 16884 17668 16894
rect 17612 16790 17668 16828
rect 18620 16324 18676 16942
rect 18620 16258 18676 16268
rect 18956 16994 19012 17006
rect 18956 16942 18958 16994
rect 19010 16942 19012 16994
rect 18956 16212 19012 16942
rect 18844 16156 19012 16212
rect 18396 16100 18452 16110
rect 18396 16006 18452 16044
rect 18508 15988 18564 15998
rect 18284 14756 18340 14766
rect 18060 14530 18116 14542
rect 18060 14478 18062 14530
rect 18114 14478 18116 14530
rect 17612 14418 17668 14430
rect 17612 14366 17614 14418
rect 17666 14366 17668 14418
rect 17612 13860 17668 14366
rect 18060 14420 18116 14478
rect 17724 14308 17780 14318
rect 17724 14306 17892 14308
rect 17724 14254 17726 14306
rect 17778 14254 17892 14306
rect 17724 14252 17892 14254
rect 17724 14242 17780 14252
rect 17612 13794 17668 13804
rect 17612 13636 17668 13674
rect 17612 13570 17668 13580
rect 17724 13522 17780 13534
rect 17724 13470 17726 13522
rect 17778 13470 17780 13522
rect 17276 12908 17556 12964
rect 17612 13412 17668 13422
rect 16604 12740 16660 12750
rect 16380 4452 16436 4462
rect 16044 3502 16046 3554
rect 16098 3502 16100 3554
rect 16044 3490 16100 3502
rect 16156 4450 16436 4452
rect 16156 4398 16382 4450
rect 16434 4398 16436 4450
rect 16156 4396 16436 4398
rect 15484 3164 15988 3220
rect 15484 800 15540 3164
rect 16156 800 16212 4396
rect 16380 4386 16436 4396
rect 16604 4338 16660 12684
rect 16604 4286 16606 4338
rect 16658 4286 16660 4338
rect 16604 4274 16660 4286
rect 17276 3554 17332 12908
rect 17388 12740 17444 12750
rect 17388 12646 17444 12684
rect 17500 12740 17556 12750
rect 17612 12740 17668 13356
rect 17724 12964 17780 13470
rect 17836 13300 17892 14252
rect 18060 13746 18116 14364
rect 18060 13694 18062 13746
rect 18114 13694 18116 13746
rect 18060 13636 18116 13694
rect 18284 13748 18340 14700
rect 18508 14754 18564 15932
rect 18732 15988 18788 15998
rect 18732 15148 18788 15932
rect 18508 14702 18510 14754
rect 18562 14702 18564 14754
rect 18508 14690 18564 14702
rect 18620 15092 18788 15148
rect 18284 13682 18340 13692
rect 18508 13860 18564 13870
rect 18508 13746 18564 13804
rect 18508 13694 18510 13746
rect 18562 13694 18564 13746
rect 18508 13682 18564 13694
rect 18060 13570 18116 13580
rect 18284 13522 18340 13534
rect 18284 13470 18286 13522
rect 18338 13470 18340 13522
rect 17836 13244 18004 13300
rect 17724 12962 17892 12964
rect 17724 12910 17726 12962
rect 17778 12910 17892 12962
rect 17724 12908 17892 12910
rect 17724 12898 17780 12908
rect 17500 12738 17668 12740
rect 17500 12686 17502 12738
rect 17554 12686 17668 12738
rect 17500 12684 17668 12686
rect 17836 12740 17892 12908
rect 17948 12962 18004 13244
rect 17948 12910 17950 12962
rect 18002 12910 18004 12962
rect 17948 12898 18004 12910
rect 18284 12740 18340 13470
rect 17836 12684 18340 12740
rect 17500 12674 17556 12684
rect 17276 3502 17278 3554
rect 17330 3502 17332 3554
rect 17276 3490 17332 3502
rect 17948 11844 18004 11854
rect 17948 3554 18004 11788
rect 17948 3502 17950 3554
rect 18002 3502 18004 3554
rect 17948 3490 18004 3502
rect 18620 3554 18676 15092
rect 18844 11844 18900 16156
rect 18956 15876 19012 15886
rect 18956 14754 19012 15820
rect 18956 14702 18958 14754
rect 19010 14702 19012 14754
rect 18956 14690 19012 14702
rect 19068 15092 19124 17388
rect 19180 16882 19236 16894
rect 19180 16830 19182 16882
rect 19234 16830 19236 16882
rect 19180 16322 19236 16830
rect 19404 16884 19460 17388
rect 19628 17106 19684 17612
rect 19964 17602 20020 17612
rect 19628 17054 19630 17106
rect 19682 17054 19684 17106
rect 19628 17042 19684 17054
rect 19740 17442 19796 17454
rect 19740 17390 19742 17442
rect 19794 17390 19796 17442
rect 19404 16818 19460 16828
rect 19180 16270 19182 16322
rect 19234 16270 19236 16322
rect 19180 16258 19236 16270
rect 19516 16324 19572 16334
rect 19740 16324 19796 17390
rect 19860 17276 20124 17286
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 19860 17210 20124 17220
rect 20188 17108 20244 18396
rect 20300 18228 20356 20636
rect 20412 20626 20468 20636
rect 20524 20242 20580 21532
rect 20524 20190 20526 20242
rect 20578 20190 20580 20242
rect 20524 20178 20580 20190
rect 20636 20804 20692 20814
rect 20636 19908 20692 20748
rect 20748 20580 20804 20590
rect 20748 20486 20804 20524
rect 20636 19234 20692 19852
rect 20636 19182 20638 19234
rect 20690 19182 20692 19234
rect 20636 19170 20692 19182
rect 21084 19796 21140 22540
rect 21420 22484 21476 23660
rect 21756 23492 21812 23502
rect 21756 23154 21812 23436
rect 21756 23102 21758 23154
rect 21810 23102 21812 23154
rect 21476 22428 21700 22484
rect 21420 21810 21476 22428
rect 21644 22370 21700 22428
rect 21644 22318 21646 22370
rect 21698 22318 21700 22370
rect 21644 22306 21700 22318
rect 21420 21758 21422 21810
rect 21474 21758 21476 21810
rect 21420 21746 21476 21758
rect 21532 22260 21588 22270
rect 21420 21588 21476 21598
rect 21420 20802 21476 21532
rect 21420 20750 21422 20802
rect 21474 20750 21476 20802
rect 21420 20020 21476 20750
rect 21420 19954 21476 19964
rect 21532 20130 21588 22204
rect 21756 21698 21812 23102
rect 21980 23156 22036 23774
rect 22092 23268 22148 23886
rect 22540 23380 22596 23390
rect 22652 23380 22708 24108
rect 22764 24098 22820 24108
rect 23772 24164 23828 24670
rect 23772 24098 23828 24108
rect 23772 23938 23828 23950
rect 23772 23886 23774 23938
rect 23826 23886 23828 23938
rect 23772 23604 23828 23886
rect 23996 23826 24052 31500
rect 24108 24946 24164 35420
rect 24522 35308 24786 35318
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24522 35242 24786 35252
rect 24522 33740 24786 33750
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24522 33674 24786 33684
rect 24522 32172 24786 32182
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24522 32106 24786 32116
rect 24522 30604 24786 30614
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24522 30538 24786 30548
rect 24522 29036 24786 29046
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24522 28970 24786 28980
rect 24522 27468 24786 27478
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24522 27402 24786 27412
rect 25900 26516 25956 36206
rect 36316 36260 36372 36270
rect 36316 36166 36372 36204
rect 29184 36092 29448 36102
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29184 36026 29448 36036
rect 33846 35308 34110 35318
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 33846 35242 34110 35252
rect 29184 34524 29448 34534
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29184 34458 29448 34468
rect 33846 33740 34110 33750
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 33846 33674 34110 33684
rect 28588 33236 28644 33246
rect 25900 26450 25956 26460
rect 27020 30884 27076 30894
rect 24522 25900 24786 25910
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24522 25834 24786 25844
rect 24108 24894 24110 24946
rect 24162 24894 24164 24946
rect 24108 24882 24164 24894
rect 25788 25506 25844 25518
rect 25788 25454 25790 25506
rect 25842 25454 25844 25506
rect 25788 24946 25844 25454
rect 26012 25508 26068 25518
rect 26012 25394 26068 25452
rect 26460 25508 26516 25518
rect 26460 25506 26628 25508
rect 26460 25454 26462 25506
rect 26514 25454 26628 25506
rect 26460 25452 26628 25454
rect 26460 25442 26516 25452
rect 26012 25342 26014 25394
rect 26066 25342 26068 25394
rect 26012 25330 26068 25342
rect 25788 24894 25790 24946
rect 25842 24894 25844 24946
rect 25788 24882 25844 24894
rect 26572 24948 26628 25452
rect 26684 25396 26740 25406
rect 26684 25302 26740 25340
rect 26684 24948 26740 24958
rect 26572 24946 26740 24948
rect 26572 24894 26686 24946
rect 26738 24894 26740 24946
rect 26572 24892 26740 24894
rect 26684 24882 26740 24892
rect 26124 24724 26180 24734
rect 26124 24630 26180 24668
rect 25228 24610 25284 24622
rect 25228 24558 25230 24610
rect 25282 24558 25284 24610
rect 24522 24332 24786 24342
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24522 24266 24786 24276
rect 24668 24164 24724 24174
rect 24668 24070 24724 24108
rect 23996 23774 23998 23826
rect 24050 23774 24052 23826
rect 23996 23762 24052 23774
rect 24892 23938 24948 23950
rect 24892 23886 24894 23938
rect 24946 23886 24948 23938
rect 24892 23828 24948 23886
rect 24892 23762 24948 23772
rect 24332 23714 24388 23726
rect 24332 23662 24334 23714
rect 24386 23662 24388 23714
rect 24332 23604 24388 23662
rect 23772 23548 24388 23604
rect 25228 23492 25284 24558
rect 25452 24500 25508 24510
rect 26348 24500 26404 24510
rect 25452 24498 26404 24500
rect 25452 24446 25454 24498
rect 25506 24446 26350 24498
rect 26402 24446 26404 24498
rect 25452 24444 26404 24446
rect 25452 24164 25508 24444
rect 25452 24098 25508 24108
rect 25340 23828 25396 23838
rect 25340 23734 25396 23772
rect 25116 23436 25228 23492
rect 22540 23378 22708 23380
rect 22540 23326 22542 23378
rect 22594 23326 22708 23378
rect 22540 23324 22708 23326
rect 23884 23380 23940 23390
rect 22540 23314 22596 23324
rect 23884 23286 23940 23324
rect 22092 23174 22148 23212
rect 23212 23266 23268 23278
rect 23212 23214 23214 23266
rect 23266 23214 23268 23266
rect 22876 23156 22932 23166
rect 21980 23062 22036 23100
rect 22428 23154 22932 23156
rect 22428 23102 22878 23154
rect 22930 23102 22932 23154
rect 22428 23100 22932 23102
rect 22428 22594 22484 23100
rect 22876 23090 22932 23100
rect 22428 22542 22430 22594
rect 22482 22542 22484 22594
rect 22428 22530 22484 22542
rect 23212 22596 23268 23214
rect 23212 22530 23268 22540
rect 23548 23154 23604 23166
rect 23548 23102 23550 23154
rect 23602 23102 23604 23154
rect 21756 21646 21758 21698
rect 21810 21646 21812 21698
rect 21756 21634 21812 21646
rect 21868 22258 21924 22270
rect 21868 22206 21870 22258
rect 21922 22206 21924 22258
rect 21868 21698 21924 22206
rect 21868 21646 21870 21698
rect 21922 21646 21924 21698
rect 21868 21028 21924 21646
rect 21532 20078 21534 20130
rect 21586 20078 21588 20130
rect 21084 19124 21140 19740
rect 21532 19348 21588 20078
rect 21644 20972 21924 21028
rect 21980 22258 22036 22270
rect 21980 22206 21982 22258
rect 22034 22206 22036 22258
rect 21980 21698 22036 22206
rect 22428 22260 22484 22270
rect 22428 21810 22484 22204
rect 23548 22260 23604 23102
rect 24522 22764 24786 22774
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24522 22698 24786 22708
rect 25116 22370 25172 23436
rect 25228 23426 25284 23436
rect 25564 23378 25620 24444
rect 26012 24162 26068 24444
rect 26348 24434 26404 24444
rect 26012 24110 26014 24162
rect 26066 24110 26068 24162
rect 26012 24098 26068 24110
rect 25788 23940 25844 23950
rect 25788 23846 25844 23884
rect 26236 23940 26292 23950
rect 25564 23326 25566 23378
rect 25618 23326 25620 23378
rect 25564 23314 25620 23326
rect 26012 23492 26068 23502
rect 26012 23378 26068 23436
rect 26012 23326 26014 23378
rect 26066 23326 26068 23378
rect 26012 23314 26068 23326
rect 25340 23156 25396 23166
rect 26124 23156 26180 23166
rect 25340 23154 25732 23156
rect 25340 23102 25342 23154
rect 25394 23102 25732 23154
rect 25340 23100 25732 23102
rect 25340 23090 25396 23100
rect 25116 22318 25118 22370
rect 25170 22318 25172 22370
rect 25116 22306 25172 22318
rect 23548 22194 23604 22204
rect 25228 22258 25284 22270
rect 25228 22206 25230 22258
rect 25282 22206 25284 22258
rect 22428 21758 22430 21810
rect 22482 21758 22484 21810
rect 22428 21746 22484 21758
rect 23100 21812 23156 21822
rect 23100 21718 23156 21756
rect 21980 21646 21982 21698
rect 22034 21646 22036 21698
rect 21644 20802 21700 20972
rect 21644 20750 21646 20802
rect 21698 20750 21700 20802
rect 21644 20692 21700 20750
rect 21644 20130 21700 20636
rect 21644 20078 21646 20130
rect 21698 20078 21700 20130
rect 21644 20066 21700 20078
rect 21756 20804 21812 20814
rect 21980 20804 22036 21646
rect 24444 21700 24500 21710
rect 22764 21588 22820 21598
rect 22204 21586 22820 21588
rect 22204 21534 22766 21586
rect 22818 21534 22820 21586
rect 22204 21532 22820 21534
rect 22204 21026 22260 21532
rect 22764 21522 22820 21532
rect 23660 21588 23716 21598
rect 22204 20974 22206 21026
rect 22258 20974 22260 21026
rect 22204 20962 22260 20974
rect 23548 20916 23604 20926
rect 21756 20802 22036 20804
rect 21756 20750 21758 20802
rect 21810 20750 22036 20802
rect 21756 20748 22036 20750
rect 22764 20802 22820 20814
rect 22764 20750 22766 20802
rect 22818 20750 22820 20802
rect 21756 20580 21812 20748
rect 22540 20692 22596 20702
rect 22540 20598 22596 20636
rect 21756 20130 21812 20524
rect 22764 20468 22820 20750
rect 23212 20692 23268 20702
rect 21756 20078 21758 20130
rect 21810 20078 21812 20130
rect 21756 20066 21812 20078
rect 22092 20412 22820 20468
rect 22988 20690 23268 20692
rect 22988 20638 23214 20690
rect 23266 20638 23268 20690
rect 22988 20636 23268 20638
rect 22092 20132 22148 20412
rect 22988 20356 23044 20636
rect 23212 20626 23268 20636
rect 23548 20690 23604 20860
rect 23548 20638 23550 20690
rect 23602 20638 23604 20690
rect 23548 20626 23604 20638
rect 22204 20300 23044 20356
rect 22204 20242 22260 20300
rect 22204 20190 22206 20242
rect 22258 20190 22260 20242
rect 22204 20178 22260 20190
rect 23660 20242 23716 21532
rect 24332 21588 24388 21598
rect 24332 21494 24388 21532
rect 23884 21364 23940 21374
rect 24444 21364 24500 21644
rect 25228 21700 25284 22206
rect 25340 22258 25396 22270
rect 25340 22206 25342 22258
rect 25394 22206 25396 22258
rect 25340 22148 25396 22206
rect 25340 22092 25620 22148
rect 25284 21644 25396 21700
rect 25228 21634 25284 21644
rect 23884 21362 24164 21364
rect 23884 21310 23886 21362
rect 23938 21310 24164 21362
rect 23884 21308 24164 21310
rect 23884 21298 23940 21308
rect 24108 20802 24164 21308
rect 24108 20750 24110 20802
rect 24162 20750 24164 20802
rect 24108 20738 24164 20750
rect 24332 21308 24500 21364
rect 24668 21586 24724 21598
rect 24668 21534 24670 21586
rect 24722 21534 24724 21586
rect 24668 21364 24724 21534
rect 23660 20190 23662 20242
rect 23714 20190 23716 20242
rect 23660 20178 23716 20190
rect 24332 20242 24388 21308
rect 24668 21298 24724 21308
rect 24522 21196 24786 21206
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24522 21130 24786 21140
rect 25340 21140 25396 21644
rect 25564 21588 25620 22092
rect 25452 21474 25508 21486
rect 25452 21422 25454 21474
rect 25506 21422 25508 21474
rect 25452 21364 25508 21422
rect 25452 21298 25508 21308
rect 25340 21084 25508 21140
rect 24444 21028 24500 21038
rect 24444 20690 24500 20972
rect 25452 20802 25508 21084
rect 25452 20750 25454 20802
rect 25506 20750 25508 20802
rect 25452 20738 25508 20750
rect 25564 20802 25620 21532
rect 25564 20750 25566 20802
rect 25618 20750 25620 20802
rect 25564 20738 25620 20750
rect 24444 20638 24446 20690
rect 24498 20638 24500 20690
rect 24444 20626 24500 20638
rect 25340 20692 25396 20702
rect 25340 20598 25396 20636
rect 24332 20190 24334 20242
rect 24386 20190 24388 20242
rect 24332 20178 24388 20190
rect 22092 20066 22148 20076
rect 23996 20132 24052 20142
rect 22652 20020 22708 20030
rect 22652 19926 22708 19964
rect 23436 20018 23492 20030
rect 23436 19966 23438 20018
rect 23490 19966 23492 20018
rect 21532 19282 21588 19292
rect 22428 19684 22484 19694
rect 21868 19236 21924 19246
rect 21084 19058 21140 19068
rect 21532 19122 21588 19134
rect 21532 19070 21534 19122
rect 21586 19070 21588 19122
rect 20300 18162 20356 18172
rect 20412 19012 20468 19022
rect 20412 19010 21028 19012
rect 20412 18958 20414 19010
rect 20466 18958 21028 19010
rect 20412 18956 21028 18958
rect 20412 17108 20468 18956
rect 20972 18562 21028 18956
rect 21532 18674 21588 19070
rect 21868 19122 21924 19180
rect 21868 19070 21870 19122
rect 21922 19070 21924 19122
rect 21868 19058 21924 19070
rect 21532 18622 21534 18674
rect 21586 18622 21588 18674
rect 21532 18610 21588 18622
rect 20972 18510 20974 18562
rect 21026 18510 21028 18562
rect 20972 18498 21028 18510
rect 20860 18450 20916 18462
rect 20860 18398 20862 18450
rect 20914 18398 20916 18450
rect 20860 18340 20916 18398
rect 21084 18452 21140 18462
rect 21084 18358 21140 18396
rect 21756 18452 21812 18462
rect 20860 18274 20916 18284
rect 21308 17780 21364 17790
rect 20524 17778 21364 17780
rect 20524 17726 21310 17778
rect 21362 17726 21364 17778
rect 20524 17724 21364 17726
rect 20524 17666 20580 17724
rect 21308 17714 21364 17724
rect 21756 17668 21812 18396
rect 20524 17614 20526 17666
rect 20578 17614 20580 17666
rect 20524 17602 20580 17614
rect 21420 17666 21812 17668
rect 21420 17614 21758 17666
rect 21810 17614 21812 17666
rect 21420 17612 21812 17614
rect 21420 17556 21476 17612
rect 21756 17602 21812 17612
rect 21980 18340 22036 18350
rect 21196 17500 21476 17556
rect 21868 17554 21924 17566
rect 21868 17502 21870 17554
rect 21922 17502 21924 17554
rect 20748 17444 20804 17454
rect 20748 17350 20804 17388
rect 20076 17052 20244 17108
rect 20300 17052 20468 17108
rect 20076 16994 20132 17052
rect 20076 16942 20078 16994
rect 20130 16942 20132 16994
rect 20076 16930 20132 16942
rect 20300 16996 20356 17052
rect 20188 16884 20244 16894
rect 20300 16884 20356 16940
rect 21084 16996 21140 17006
rect 21084 16902 21140 16940
rect 21196 16994 21252 17500
rect 21868 17444 21924 17502
rect 21196 16942 21198 16994
rect 21250 16942 21252 16994
rect 21196 16930 21252 16942
rect 21532 17388 21924 17444
rect 21532 16996 21588 17388
rect 21980 17332 22036 18284
rect 22092 17666 22148 17678
rect 22092 17614 22094 17666
rect 22146 17614 22148 17666
rect 22092 17556 22148 17614
rect 22092 17490 22148 17500
rect 21980 17276 22148 17332
rect 21532 16930 21588 16940
rect 20188 16882 20356 16884
rect 20188 16830 20190 16882
rect 20242 16830 20356 16882
rect 20188 16828 20356 16830
rect 20412 16884 20468 16894
rect 20188 16818 20244 16828
rect 20412 16790 20468 16828
rect 20972 16882 21028 16894
rect 20972 16830 20974 16882
rect 21026 16830 21028 16882
rect 19516 16230 19572 16268
rect 19628 16268 19796 16324
rect 20524 16324 20580 16334
rect 20972 16324 21028 16830
rect 21644 16884 21700 16894
rect 21980 16884 22036 16894
rect 21644 16882 22036 16884
rect 21644 16830 21646 16882
rect 21698 16830 21982 16882
rect 22034 16830 22036 16882
rect 21644 16828 22036 16830
rect 21644 16818 21700 16828
rect 21980 16818 22036 16828
rect 21532 16324 21588 16334
rect 20972 16268 21364 16324
rect 19068 14532 19124 15036
rect 19068 14466 19124 14476
rect 19404 14756 19460 14766
rect 19404 14530 19460 14700
rect 19404 14478 19406 14530
rect 19458 14478 19460 14530
rect 19404 14466 19460 14478
rect 19180 14420 19236 14430
rect 19180 14326 19236 14364
rect 19068 14308 19124 14318
rect 19068 14214 19124 14252
rect 19516 13860 19572 13870
rect 19292 13858 19572 13860
rect 19292 13806 19518 13858
rect 19570 13806 19572 13858
rect 19292 13804 19572 13806
rect 18956 13748 19012 13758
rect 19180 13748 19236 13758
rect 18956 13746 19236 13748
rect 18956 13694 18958 13746
rect 19010 13694 19182 13746
rect 19234 13694 19236 13746
rect 18956 13692 19236 13694
rect 18956 13682 19012 13692
rect 19180 13682 19236 13692
rect 18844 11778 18900 11788
rect 18620 3502 18622 3554
rect 18674 3502 18676 3554
rect 18620 3490 18676 3502
rect 19292 3554 19348 13804
rect 19516 13794 19572 13804
rect 19628 4564 19684 16268
rect 19740 16098 19796 16110
rect 19740 16046 19742 16098
rect 19794 16046 19796 16098
rect 19740 15092 19796 16046
rect 20188 16100 20244 16110
rect 20076 15988 20132 15998
rect 20076 15874 20132 15932
rect 20076 15822 20078 15874
rect 20130 15822 20132 15874
rect 20076 15810 20132 15822
rect 19860 15708 20124 15718
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 19860 15642 20124 15652
rect 20188 15428 20244 16044
rect 20412 15876 20468 15886
rect 20412 15782 20468 15820
rect 20188 15334 20244 15372
rect 19740 15026 19796 15036
rect 20412 14756 20468 14766
rect 20524 14756 20580 16268
rect 21308 16212 21364 16268
rect 21308 16118 21364 16156
rect 21532 15148 21588 16268
rect 21868 15876 21924 15886
rect 21868 15782 21924 15820
rect 21868 15428 21924 15438
rect 21532 15092 21700 15148
rect 20412 14754 20580 14756
rect 20412 14702 20414 14754
rect 20466 14702 20580 14754
rect 20412 14700 20580 14702
rect 20412 14690 20468 14700
rect 19740 14530 19796 14542
rect 19740 14478 19742 14530
rect 19794 14478 19796 14530
rect 19740 13972 19796 14478
rect 20188 14530 20244 14542
rect 20188 14478 20190 14530
rect 20242 14478 20244 14530
rect 19860 14140 20124 14150
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 19860 14074 20124 14084
rect 19852 13972 19908 13982
rect 19740 13970 19908 13972
rect 19740 13918 19854 13970
rect 19906 13918 19908 13970
rect 19740 13916 19908 13918
rect 19852 13906 19908 13916
rect 19964 13860 20020 13870
rect 19964 13766 20020 13804
rect 20188 12740 20244 14478
rect 20748 14308 20804 14318
rect 20636 14306 20804 14308
rect 20636 14254 20750 14306
rect 20802 14254 20804 14306
rect 20636 14252 20804 14254
rect 20636 12964 20692 14252
rect 20748 14242 20804 14252
rect 20972 13860 21028 13870
rect 20972 13858 21588 13860
rect 20972 13806 20974 13858
rect 21026 13806 21588 13858
rect 20972 13804 21588 13806
rect 20972 13794 21028 13804
rect 20748 13746 20804 13758
rect 20748 13694 20750 13746
rect 20802 13694 20804 13746
rect 20748 13636 20804 13694
rect 21308 13636 21364 13646
rect 20748 13634 21364 13636
rect 20748 13582 21310 13634
rect 21362 13582 21364 13634
rect 20748 13580 21364 13582
rect 21308 13570 21364 13580
rect 21532 12964 21588 13804
rect 21644 13746 21700 15092
rect 21868 14530 21924 15372
rect 21868 14478 21870 14530
rect 21922 14478 21924 14530
rect 21868 14466 21924 14478
rect 21644 13694 21646 13746
rect 21698 13694 21700 13746
rect 21644 13682 21700 13694
rect 21868 13636 21924 13646
rect 22092 13636 22148 17276
rect 22316 16994 22372 17006
rect 22316 16942 22318 16994
rect 22370 16942 22372 16994
rect 22316 15148 22372 16942
rect 22428 16098 22484 19628
rect 22540 19348 22596 19358
rect 22540 19254 22596 19292
rect 22988 19348 23044 19358
rect 22876 19236 22932 19246
rect 22764 19234 22932 19236
rect 22764 19182 22878 19234
rect 22930 19182 22932 19234
rect 22764 19180 22932 19182
rect 22764 18340 22820 19180
rect 22876 19170 22932 19180
rect 22764 18246 22820 18284
rect 22988 18452 23044 19292
rect 23436 19348 23492 19966
rect 23996 19460 24052 20076
rect 24522 19628 24786 19638
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24522 19562 24786 19572
rect 23996 19404 24388 19460
rect 23436 19282 23492 19292
rect 23100 19124 23156 19134
rect 23100 18676 23156 19068
rect 23212 19124 23268 19134
rect 23996 19124 24052 19134
rect 23212 19122 23492 19124
rect 23212 19070 23214 19122
rect 23266 19070 23492 19122
rect 23212 19068 23492 19070
rect 23212 19058 23268 19068
rect 23436 18676 23492 19068
rect 23996 19030 24052 19068
rect 24332 19124 24388 19404
rect 25676 19236 25732 23100
rect 25788 22146 25844 22158
rect 25788 22094 25790 22146
rect 25842 22094 25844 22146
rect 25788 21698 25844 22094
rect 26124 21810 26180 23100
rect 26236 22370 26292 23884
rect 26348 23828 26404 23838
rect 26684 23828 26740 23838
rect 26348 23826 26740 23828
rect 26348 23774 26350 23826
rect 26402 23774 26686 23826
rect 26738 23774 26740 23826
rect 26348 23772 26740 23774
rect 26348 23762 26404 23772
rect 26684 23762 26740 23772
rect 27020 23826 27076 30828
rect 27804 27188 27860 27198
rect 27692 27132 27804 27188
rect 27132 25284 27188 25294
rect 27132 25282 27300 25284
rect 27132 25230 27134 25282
rect 27186 25230 27300 25282
rect 27132 25228 27300 25230
rect 27132 25218 27188 25228
rect 27020 23774 27022 23826
rect 27074 23774 27076 23826
rect 27020 23762 27076 23774
rect 27132 24948 27188 24958
rect 27132 23716 27188 24892
rect 27244 24724 27300 25228
rect 27244 24658 27300 24668
rect 27580 24500 27636 24510
rect 27580 24162 27636 24444
rect 27580 24110 27582 24162
rect 27634 24110 27636 24162
rect 27580 24098 27636 24110
rect 27132 23650 27188 23660
rect 27356 23938 27412 23950
rect 27356 23886 27358 23938
rect 27410 23886 27412 23938
rect 27356 23828 27412 23886
rect 26236 22318 26238 22370
rect 26290 22318 26292 22370
rect 26236 22306 26292 22318
rect 27356 23268 27412 23772
rect 26124 21758 26126 21810
rect 26178 21758 26180 21810
rect 26124 21746 26180 21758
rect 26348 22258 26404 22270
rect 26348 22206 26350 22258
rect 26402 22206 26404 22258
rect 25788 21646 25790 21698
rect 25842 21646 25844 21698
rect 25788 21634 25844 21646
rect 26348 21700 26404 22206
rect 26460 22260 26516 22270
rect 26908 22260 26964 22270
rect 27244 22260 27300 22270
rect 26460 22258 26628 22260
rect 26460 22206 26462 22258
rect 26514 22206 26628 22258
rect 26460 22204 26628 22206
rect 26460 22194 26516 22204
rect 26348 21634 26404 21644
rect 26460 21586 26516 21598
rect 26460 21534 26462 21586
rect 26514 21534 26516 21586
rect 25788 20692 25844 20702
rect 25788 20242 25844 20636
rect 26012 20692 26068 20702
rect 26348 20692 26404 20702
rect 26012 20690 26404 20692
rect 26012 20638 26014 20690
rect 26066 20638 26350 20690
rect 26402 20638 26404 20690
rect 26012 20636 26404 20638
rect 26012 20626 26068 20636
rect 26348 20626 26404 20636
rect 26460 20356 26516 21534
rect 26572 21588 26628 22204
rect 26908 22258 27300 22260
rect 26908 22206 26910 22258
rect 26962 22206 27246 22258
rect 27298 22206 27300 22258
rect 26908 22204 27300 22206
rect 26908 22194 26964 22204
rect 27244 22194 27300 22204
rect 27356 22036 27412 23212
rect 27580 22260 27636 22270
rect 27692 22260 27748 27132
rect 27804 27122 27860 27132
rect 28364 25506 28420 25518
rect 28364 25454 28366 25506
rect 28418 25454 28420 25506
rect 28364 24946 28420 25454
rect 28588 25394 28644 33180
rect 29184 32956 29448 32966
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29184 32890 29448 32900
rect 33846 32172 34110 32182
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 33846 32106 34110 32116
rect 36540 31948 36596 36316
rect 36876 36372 36932 36382
rect 36876 36278 36932 36316
rect 37212 36258 37268 36270
rect 37212 36206 37214 36258
rect 37266 36206 37268 36258
rect 37100 35700 37156 35710
rect 37100 35606 37156 35644
rect 37212 35252 37268 36206
rect 37660 35922 37716 36428
rect 37884 36260 37940 36270
rect 37660 35870 37662 35922
rect 37714 35870 37716 35922
rect 37660 35858 37716 35870
rect 37772 36258 37940 36260
rect 37772 36206 37886 36258
rect 37938 36206 37940 36258
rect 37772 36204 37940 36206
rect 37212 35186 37268 35196
rect 37772 34916 37828 36204
rect 37884 36194 37940 36204
rect 38220 36260 38276 36270
rect 38276 36204 38388 36260
rect 38220 36166 38276 36204
rect 38220 35810 38276 35822
rect 38220 35758 38222 35810
rect 38274 35758 38276 35810
rect 37996 35700 38052 35710
rect 38052 35644 38164 35700
rect 37996 35606 38052 35644
rect 36428 31892 36596 31948
rect 36988 34860 37828 34916
rect 29184 31388 29448 31398
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29184 31322 29448 31332
rect 33846 30604 34110 30614
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 33846 30538 34110 30548
rect 29184 29820 29448 29830
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29184 29754 29448 29764
rect 33846 29036 34110 29046
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 33846 28970 34110 28980
rect 29184 28252 29448 28262
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29184 28186 29448 28196
rect 30380 27860 30436 27870
rect 29184 26684 29448 26694
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29184 26618 29448 26628
rect 29148 25396 29204 25406
rect 28588 25342 28590 25394
rect 28642 25342 28644 25394
rect 28588 25330 28644 25342
rect 29036 25394 29204 25396
rect 29036 25342 29150 25394
rect 29202 25342 29204 25394
rect 29036 25340 29204 25342
rect 28364 24894 28366 24946
rect 28418 24894 28420 24946
rect 28364 24882 28420 24894
rect 28700 24948 28756 24958
rect 29036 24948 29092 25340
rect 29148 25330 29204 25340
rect 29484 25396 29540 25406
rect 29484 25302 29540 25340
rect 29184 25116 29448 25126
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29184 25050 29448 25060
rect 29260 24948 29316 24958
rect 29036 24946 29316 24948
rect 29036 24894 29262 24946
rect 29314 24894 29316 24946
rect 29036 24892 29316 24894
rect 27804 24724 27860 24734
rect 27804 24630 27860 24668
rect 28588 24724 28644 24734
rect 28028 24500 28084 24510
rect 28028 24406 28084 24444
rect 28364 24500 28420 24510
rect 27916 23828 27972 23838
rect 28252 23828 28308 23838
rect 27916 23826 28308 23828
rect 27916 23774 27918 23826
rect 27970 23774 28254 23826
rect 28306 23774 28308 23826
rect 27916 23772 28308 23774
rect 27916 23762 27972 23772
rect 28252 23762 28308 23772
rect 28140 23380 28196 23390
rect 28364 23380 28420 24444
rect 28588 24052 28644 24668
rect 28700 24722 28756 24892
rect 29260 24882 29316 24892
rect 30156 24948 30212 24958
rect 28700 24670 28702 24722
rect 28754 24670 28756 24722
rect 28700 24658 28756 24670
rect 29708 24724 29764 24734
rect 29708 24630 29764 24668
rect 28924 24500 28980 24510
rect 28980 24444 29428 24500
rect 28924 24406 28980 24444
rect 28812 24164 28868 24174
rect 28588 23996 28756 24052
rect 28588 23828 28644 23838
rect 28588 23734 28644 23772
rect 28140 23378 28420 23380
rect 28140 23326 28142 23378
rect 28194 23326 28420 23378
rect 28140 23324 28420 23326
rect 28140 23314 28196 23324
rect 28476 23268 28532 23278
rect 27580 22258 27748 22260
rect 27580 22206 27582 22258
rect 27634 22206 27748 22258
rect 27580 22204 27748 22206
rect 28364 23154 28420 23166
rect 28364 23102 28366 23154
rect 28418 23102 28420 23154
rect 27580 22194 27636 22204
rect 27244 21980 27412 22036
rect 26796 21700 26852 21710
rect 26796 21606 26852 21644
rect 27244 21698 27300 21980
rect 27244 21646 27246 21698
rect 27298 21646 27300 21698
rect 26572 21522 26628 21532
rect 27244 21364 27300 21646
rect 27468 21700 27524 21710
rect 27468 21606 27524 21644
rect 27244 21298 27300 21308
rect 27356 21588 27412 21598
rect 27020 20692 27076 20702
rect 26908 20690 27076 20692
rect 26908 20638 27022 20690
rect 27074 20638 27076 20690
rect 26908 20636 27076 20638
rect 26684 20580 26740 20590
rect 26684 20486 26740 20524
rect 26460 20300 26740 20356
rect 25788 20190 25790 20242
rect 25842 20190 25844 20242
rect 25788 20178 25844 20190
rect 26348 20132 26404 20142
rect 26348 20130 26628 20132
rect 26348 20078 26350 20130
rect 26402 20078 26628 20130
rect 26348 20076 26628 20078
rect 26348 20066 26404 20076
rect 26012 20018 26068 20030
rect 26012 19966 26014 20018
rect 26066 19966 26068 20018
rect 26012 19908 26068 19966
rect 26012 19842 26068 19852
rect 25452 19180 25732 19236
rect 26012 19348 26068 19358
rect 26012 19234 26068 19292
rect 26012 19182 26014 19234
rect 26066 19182 26068 19234
rect 24332 19030 24388 19068
rect 24668 19122 24724 19134
rect 24668 19070 24670 19122
rect 24722 19070 24724 19122
rect 23660 19012 23716 19022
rect 23660 19010 23940 19012
rect 23660 18958 23662 19010
rect 23714 18958 23940 19010
rect 23660 18956 23940 18958
rect 23660 18946 23716 18956
rect 23884 18900 23940 18956
rect 24668 18900 24724 19070
rect 25340 19124 25396 19134
rect 25340 19030 25396 19068
rect 25004 19012 25060 19022
rect 25004 19010 25172 19012
rect 25004 18958 25006 19010
rect 25058 18958 25172 19010
rect 25004 18956 25172 18958
rect 25004 18946 25060 18956
rect 23884 18844 24724 18900
rect 23100 18620 23268 18676
rect 23100 18452 23156 18462
rect 22988 18450 23156 18452
rect 22988 18398 23102 18450
rect 23154 18398 23156 18450
rect 22988 18396 23156 18398
rect 22988 18228 23044 18396
rect 23100 18386 23156 18396
rect 22988 18162 23044 18172
rect 23212 17666 23268 18620
rect 23212 17614 23214 17666
rect 23266 17614 23268 17666
rect 22652 17556 22708 17566
rect 22652 17462 22708 17500
rect 23100 17556 23156 17566
rect 23100 17462 23156 17500
rect 23212 17444 23268 17614
rect 23324 18674 23492 18676
rect 23324 18622 23438 18674
rect 23490 18622 23492 18674
rect 23324 18620 23492 18622
rect 23324 17668 23380 18620
rect 23436 18610 23492 18620
rect 24444 18562 24500 18574
rect 24444 18510 24446 18562
rect 24498 18510 24500 18562
rect 24108 18452 24164 18462
rect 23772 18450 24164 18452
rect 23772 18398 24110 18450
rect 24162 18398 24164 18450
rect 23772 18396 24164 18398
rect 23772 17890 23828 18396
rect 24108 18386 24164 18396
rect 24444 18228 24500 18510
rect 24444 18162 24500 18172
rect 24522 18060 24786 18070
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24522 17994 24786 18004
rect 23772 17838 23774 17890
rect 23826 17838 23828 17890
rect 23772 17826 23828 17838
rect 23324 17666 23604 17668
rect 23324 17614 23326 17666
rect 23378 17614 23604 17666
rect 23324 17612 23604 17614
rect 23324 17602 23380 17612
rect 23212 17388 23492 17444
rect 22876 16884 22932 16894
rect 22876 16790 22932 16828
rect 23212 16660 23268 17388
rect 23436 16994 23492 17388
rect 23436 16942 23438 16994
rect 23490 16942 23492 16994
rect 23436 16930 23492 16942
rect 23548 16994 23604 17612
rect 23548 16942 23550 16994
rect 23602 16942 23604 16994
rect 23324 16884 23380 16894
rect 23324 16790 23380 16828
rect 23548 16660 23604 16942
rect 23212 16604 23380 16660
rect 23100 16212 23156 16222
rect 22428 16046 22430 16098
rect 22482 16046 22484 16098
rect 22428 16034 22484 16046
rect 22764 16100 22820 16110
rect 22764 15986 22820 16044
rect 23100 16100 23156 16156
rect 23100 16098 23268 16100
rect 23100 16046 23102 16098
rect 23154 16046 23268 16098
rect 23100 16044 23268 16046
rect 23100 16034 23156 16044
rect 22764 15934 22766 15986
rect 22818 15934 22820 15986
rect 22764 15922 22820 15934
rect 23212 15314 23268 16044
rect 23324 16098 23380 16604
rect 23324 16046 23326 16098
rect 23378 16046 23380 16098
rect 23324 16034 23380 16046
rect 23436 16604 23604 16660
rect 23660 17556 23716 17566
rect 23436 16098 23492 16604
rect 23436 16046 23438 16098
rect 23490 16046 23492 16098
rect 23436 16034 23492 16046
rect 23548 16100 23604 16110
rect 23212 15262 23214 15314
rect 23266 15262 23268 15314
rect 23212 15204 23268 15262
rect 23436 15204 23492 15242
rect 23548 15204 23604 16044
rect 23436 15202 23604 15204
rect 23436 15150 23438 15202
rect 23490 15150 23604 15202
rect 23436 15148 23604 15150
rect 22316 15092 22932 15148
rect 23212 15138 23268 15148
rect 21924 13580 22148 13636
rect 22316 13636 22372 13646
rect 21868 13542 21924 13580
rect 22316 13542 22372 13580
rect 22764 13636 22820 13646
rect 22764 13542 22820 13580
rect 21980 12964 22036 12974
rect 21532 12908 21924 12964
rect 20636 12898 20692 12908
rect 20188 12674 20244 12684
rect 21420 12740 21476 12750
rect 21756 12740 21812 12750
rect 21420 12646 21476 12684
rect 21532 12738 21812 12740
rect 21532 12686 21758 12738
rect 21810 12686 21812 12738
rect 21532 12684 21812 12686
rect 19860 12572 20124 12582
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 19860 12506 20124 12516
rect 19860 11004 20124 11014
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 19860 10938 20124 10948
rect 19860 9436 20124 9446
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 19860 9370 20124 9380
rect 19860 7868 20124 7878
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 19860 7802 20124 7812
rect 19860 6300 20124 6310
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 19860 6234 20124 6244
rect 19860 4732 20124 4742
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 19860 4666 20124 4676
rect 19628 4508 19908 4564
rect 19292 3502 19294 3554
rect 19346 3502 19348 3554
rect 19292 3490 19348 3502
rect 19852 3554 19908 4508
rect 19852 3502 19854 3554
rect 19906 3502 19908 3554
rect 19852 3490 19908 3502
rect 21420 3556 21476 3566
rect 21532 3556 21588 12684
rect 21756 12674 21812 12684
rect 21420 3554 21588 3556
rect 21420 3502 21422 3554
rect 21474 3502 21588 3554
rect 21420 3500 21588 3502
rect 21868 3556 21924 12908
rect 21980 12870 22036 12908
rect 22764 11844 22820 11854
rect 21980 3556 22036 3566
rect 21868 3554 22036 3556
rect 21868 3502 21982 3554
rect 22034 3502 22036 3554
rect 21868 3500 22036 3502
rect 21420 3490 21476 3500
rect 21980 3490 22036 3500
rect 22764 3554 22820 11788
rect 22876 9380 22932 15092
rect 23324 15092 23492 15148
rect 23324 13860 23380 15092
rect 22988 13804 23380 13860
rect 22988 13746 23044 13804
rect 22988 13694 22990 13746
rect 23042 13694 23044 13746
rect 22988 13682 23044 13694
rect 23324 13748 23380 13804
rect 23548 14418 23604 14430
rect 23548 14366 23550 14418
rect 23602 14366 23604 14418
rect 23548 13860 23604 14366
rect 23548 13794 23604 13804
rect 23324 13682 23380 13692
rect 23660 13634 23716 17500
rect 24332 17556 24388 17566
rect 24668 17556 24724 17566
rect 24332 17462 24388 17500
rect 24444 17554 24724 17556
rect 24444 17502 24670 17554
rect 24722 17502 24724 17554
rect 24444 17500 24724 17502
rect 24444 17220 24500 17500
rect 24668 17490 24724 17500
rect 24780 17556 24836 17566
rect 23996 17164 24500 17220
rect 23996 17106 24052 17164
rect 23996 17054 23998 17106
rect 24050 17054 24052 17106
rect 23996 17042 24052 17054
rect 24668 17108 24724 17118
rect 24780 17108 24836 17500
rect 25004 17444 25060 17454
rect 24668 17106 24836 17108
rect 24668 17054 24670 17106
rect 24722 17054 24836 17106
rect 24668 17052 24836 17054
rect 24892 17442 25060 17444
rect 24892 17390 25006 17442
rect 25058 17390 25060 17442
rect 24892 17388 25060 17390
rect 24668 17042 24724 17052
rect 24332 16884 24388 16894
rect 23884 16882 24388 16884
rect 23884 16830 24334 16882
rect 24386 16830 24388 16882
rect 23884 16828 24388 16830
rect 23884 16322 23940 16828
rect 24332 16818 24388 16828
rect 23884 16270 23886 16322
rect 23938 16270 23940 16322
rect 23884 16258 23940 16270
rect 24220 16660 24276 16670
rect 24220 16212 24276 16604
rect 24522 16492 24786 16502
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24522 16426 24786 16436
rect 24220 16118 24276 16156
rect 24444 16100 24500 16110
rect 24444 16006 24500 16044
rect 24780 15988 24836 15998
rect 24780 15894 24836 15932
rect 24332 15876 24388 15886
rect 24108 15426 24164 15438
rect 24108 15374 24110 15426
rect 24162 15374 24164 15426
rect 23772 15316 23828 15326
rect 23772 15222 23828 15260
rect 23884 13748 23940 13758
rect 23884 13654 23940 13692
rect 23660 13582 23662 13634
rect 23714 13582 23716 13634
rect 23324 13522 23380 13534
rect 23324 13470 23326 13522
rect 23378 13470 23380 13522
rect 23324 12962 23380 13470
rect 23324 12910 23326 12962
rect 23378 12910 23380 12962
rect 23324 12898 23380 12910
rect 23548 12738 23604 12750
rect 23548 12686 23550 12738
rect 23602 12686 23604 12738
rect 22876 9324 23380 9380
rect 22764 3502 22766 3554
rect 22818 3502 22820 3554
rect 22764 3490 22820 3502
rect 23324 3554 23380 9324
rect 23548 5012 23604 12686
rect 23660 12740 23716 13582
rect 23660 12674 23716 12684
rect 24108 11844 24164 15374
rect 24332 15314 24388 15820
rect 24332 15262 24334 15314
rect 24386 15262 24388 15314
rect 24332 15250 24388 15262
rect 24220 15204 24276 15214
rect 24220 15092 24388 15148
rect 24220 13748 24276 13758
rect 24220 13654 24276 13692
rect 24108 11778 24164 11788
rect 23548 4946 23604 4956
rect 23324 3502 23326 3554
rect 23378 3502 23380 3554
rect 23324 3490 23380 3502
rect 24108 3556 24164 3566
rect 16380 3442 16436 3454
rect 16380 3390 16382 3442
rect 16434 3390 16436 3442
rect 16380 3388 16436 3390
rect 24108 3442 24164 3500
rect 24108 3390 24110 3442
rect 24162 3390 24164 3442
rect 16380 3332 16884 3388
rect 16828 800 16884 3332
rect 17500 3330 17556 3342
rect 17500 3278 17502 3330
rect 17554 3278 17556 3330
rect 17500 800 17556 3278
rect 18172 3330 18228 3342
rect 18172 3278 18174 3330
rect 18226 3278 18228 3330
rect 18172 800 18228 3278
rect 18844 3330 18900 3342
rect 18844 3278 18846 3330
rect 18898 3278 18900 3330
rect 18844 800 18900 3278
rect 19516 3330 19572 3342
rect 19516 3278 19518 3330
rect 19570 3278 19572 3330
rect 19516 800 19572 3278
rect 20188 3330 20244 3342
rect 21084 3332 21140 3342
rect 21756 3332 21812 3342
rect 22428 3332 22484 3342
rect 23100 3332 23156 3342
rect 20188 3278 20190 3330
rect 20242 3278 20244 3330
rect 19860 3164 20124 3174
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 19860 3098 20124 3108
rect 20188 800 20244 3278
rect 20860 3330 21140 3332
rect 20860 3278 21086 3330
rect 21138 3278 21140 3330
rect 20860 3276 21140 3278
rect 20860 800 20916 3276
rect 21084 3266 21140 3276
rect 21532 3330 21812 3332
rect 21532 3278 21758 3330
rect 21810 3278 21812 3330
rect 21532 3276 21812 3278
rect 21532 800 21588 3276
rect 21756 3266 21812 3276
rect 22204 3330 22484 3332
rect 22204 3278 22430 3330
rect 22482 3278 22484 3330
rect 22204 3276 22484 3278
rect 22204 800 22260 3276
rect 22428 3266 22484 3276
rect 22876 3330 23156 3332
rect 22876 3278 23102 3330
rect 23154 3278 23156 3330
rect 22876 3276 23156 3278
rect 22876 800 22932 3276
rect 23100 3266 23156 3276
rect 24108 2212 24164 3390
rect 23548 2156 24164 2212
rect 24220 3444 24276 3454
rect 24332 3444 24388 15092
rect 24522 14924 24786 14934
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24522 14858 24786 14868
rect 24668 13636 24724 13646
rect 24668 13542 24724 13580
rect 24522 13356 24786 13366
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24522 13290 24786 13300
rect 24444 12740 24500 12750
rect 24444 12646 24500 12684
rect 24522 11788 24786 11798
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24522 11722 24786 11732
rect 24522 10220 24786 10230
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24522 10154 24786 10164
rect 24522 8652 24786 8662
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24522 8586 24786 8596
rect 24892 8036 24948 17388
rect 25004 17378 25060 17388
rect 25116 16212 25172 18956
rect 25452 17108 25508 19180
rect 26012 19170 26068 19182
rect 25676 19012 25732 19022
rect 25676 18918 25732 18956
rect 26348 19012 26404 19022
rect 26348 18918 26404 18956
rect 26572 18564 26628 20076
rect 26684 20130 26740 20300
rect 26684 20078 26686 20130
rect 26738 20078 26740 20130
rect 26684 19796 26740 20078
rect 26908 19908 26964 20636
rect 27020 20626 27076 20636
rect 27356 20690 27412 21532
rect 27916 21362 27972 21374
rect 27916 21310 27918 21362
rect 27970 21310 27972 21362
rect 27916 20802 27972 21310
rect 27916 20750 27918 20802
rect 27970 20750 27972 20802
rect 27916 20738 27972 20750
rect 27356 20638 27358 20690
rect 27410 20638 27412 20690
rect 27356 20626 27412 20638
rect 28140 20692 28196 20702
rect 28140 20598 28196 20636
rect 27020 20132 27076 20142
rect 27020 20130 27524 20132
rect 27020 20078 27022 20130
rect 27074 20078 27524 20130
rect 27020 20076 27524 20078
rect 27020 20066 27076 20076
rect 26908 19842 26964 19852
rect 26684 19730 26740 19740
rect 27468 19234 27524 20076
rect 28252 20130 28308 20142
rect 28252 20078 28254 20130
rect 28306 20078 28308 20130
rect 27916 20018 27972 20030
rect 27916 19966 27918 20018
rect 27970 19966 27972 20018
rect 27916 19458 27972 19966
rect 28252 20020 28308 20078
rect 28252 19954 28308 19964
rect 27916 19406 27918 19458
rect 27970 19406 27972 19458
rect 27916 19394 27972 19406
rect 28364 19460 28420 23102
rect 28476 21810 28532 23212
rect 28476 21758 28478 21810
rect 28530 21758 28532 21810
rect 28476 21746 28532 21758
rect 28700 21476 28756 23996
rect 28812 21586 28868 24108
rect 29148 24164 29204 24174
rect 29148 24050 29204 24108
rect 29372 24162 29428 24444
rect 29372 24110 29374 24162
rect 29426 24110 29428 24162
rect 29372 24098 29428 24110
rect 29148 23998 29150 24050
rect 29202 23998 29204 24050
rect 29148 23986 29204 23998
rect 29708 23828 29764 23838
rect 30044 23828 30100 23838
rect 29708 23826 30100 23828
rect 29708 23774 29710 23826
rect 29762 23774 30046 23826
rect 30098 23774 30100 23826
rect 29708 23772 30100 23774
rect 29708 23762 29764 23772
rect 30044 23762 30100 23772
rect 29184 23548 29448 23558
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29184 23482 29448 23492
rect 30156 23380 30212 24892
rect 30380 23826 30436 27804
rect 33846 27468 34110 27478
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 33846 27402 34110 27412
rect 33846 25900 34110 25910
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 33846 25834 34110 25844
rect 33846 24332 34110 24342
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 33846 24266 34110 24276
rect 30380 23774 30382 23826
rect 30434 23774 30436 23826
rect 30380 23762 30436 23774
rect 29820 23378 30212 23380
rect 29820 23326 30158 23378
rect 30210 23326 30212 23378
rect 29820 23324 30212 23326
rect 28924 23268 28980 23278
rect 28924 23174 28980 23212
rect 28812 21534 28814 21586
rect 28866 21534 28868 21586
rect 28812 21522 28868 21534
rect 29036 22428 29428 22484
rect 29036 21698 29092 22428
rect 29372 22370 29428 22428
rect 29372 22318 29374 22370
rect 29426 22318 29428 22370
rect 29372 22306 29428 22318
rect 29260 22260 29316 22270
rect 29260 22166 29316 22204
rect 29484 22260 29540 22270
rect 29820 22260 29876 23324
rect 30156 23314 30212 23324
rect 31276 23492 31332 23502
rect 30492 22372 30548 22382
rect 29484 22258 29764 22260
rect 29484 22206 29486 22258
rect 29538 22206 29764 22258
rect 29484 22204 29764 22206
rect 29484 22194 29540 22204
rect 29184 21980 29448 21990
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29184 21914 29448 21924
rect 29596 21924 29652 21934
rect 29596 21810 29652 21868
rect 29596 21758 29598 21810
rect 29650 21758 29652 21810
rect 29596 21746 29652 21758
rect 29036 21646 29038 21698
rect 29090 21646 29092 21698
rect 29036 21588 29092 21646
rect 29148 21700 29204 21710
rect 29148 21606 29204 21644
rect 29708 21700 29764 22204
rect 29820 22194 29876 22204
rect 29932 22260 29988 22270
rect 30268 22260 30324 22270
rect 29932 22258 30324 22260
rect 29932 22206 29934 22258
rect 29986 22206 30270 22258
rect 30322 22206 30324 22258
rect 29932 22204 30324 22206
rect 29932 22194 29988 22204
rect 30268 22194 30324 22204
rect 30268 22036 30324 22046
rect 30268 21810 30324 21980
rect 30268 21758 30270 21810
rect 30322 21758 30324 21810
rect 30268 21746 30324 21758
rect 28700 21410 28756 21420
rect 29036 21364 29092 21532
rect 29036 21308 29428 21364
rect 29260 21140 29316 21150
rect 29260 20804 29316 21084
rect 29260 20710 29316 20748
rect 29372 20802 29428 21308
rect 29372 20750 29374 20802
rect 29426 20750 29428 20802
rect 29372 20738 29428 20750
rect 29484 20804 29540 20814
rect 29708 20804 29764 21644
rect 29932 21586 29988 21598
rect 29932 21534 29934 21586
rect 29986 21534 29988 21586
rect 29932 21026 29988 21534
rect 29932 20974 29934 21026
rect 29986 20974 29988 21026
rect 29932 20962 29988 20974
rect 30380 21476 30436 21486
rect 30380 20914 30436 21420
rect 30380 20862 30382 20914
rect 30434 20862 30436 20914
rect 30380 20850 30436 20862
rect 29484 20802 29764 20804
rect 29484 20750 29486 20802
rect 29538 20750 29764 20802
rect 29484 20748 29764 20750
rect 29484 20738 29540 20748
rect 29184 20412 29448 20422
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29184 20346 29448 20356
rect 28924 20132 28980 20142
rect 28924 20038 28980 20076
rect 30380 20132 30436 20142
rect 30492 20132 30548 22316
rect 30604 22260 30660 22270
rect 30604 22166 30660 22204
rect 30940 22258 30996 22270
rect 30940 22206 30942 22258
rect 30994 22206 30996 22258
rect 30940 21924 30996 22206
rect 31276 22258 31332 23436
rect 33846 22764 34110 22774
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 33846 22698 34110 22708
rect 31276 22206 31278 22258
rect 31330 22206 31332 22258
rect 31276 22194 31332 22206
rect 36428 22260 36484 31892
rect 36540 31556 36596 31566
rect 36540 31462 36596 31500
rect 36988 24948 37044 34860
rect 37884 34804 37940 34814
rect 37100 34802 37940 34804
rect 37100 34750 37886 34802
rect 37938 34750 37940 34802
rect 37100 34748 37940 34750
rect 37100 25396 37156 34748
rect 37884 34738 37940 34748
rect 37996 34130 38052 34142
rect 37996 34078 37998 34130
rect 38050 34078 38052 34130
rect 37548 34020 37604 34030
rect 37996 34020 38052 34078
rect 37548 34018 38052 34020
rect 37548 33966 37550 34018
rect 37602 33966 38052 34018
rect 37548 33964 38052 33966
rect 37548 33954 37604 33964
rect 37996 33348 38052 33964
rect 38108 33460 38164 35644
rect 38220 35028 38276 35758
rect 38332 35700 38388 36204
rect 38508 36092 38772 36102
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38508 36026 38772 36036
rect 38332 35634 38388 35644
rect 39116 35252 39172 35262
rect 39172 35196 39284 35252
rect 39116 35186 39172 35196
rect 38220 34962 38276 34972
rect 38220 34692 38276 34702
rect 38220 34690 38388 34692
rect 38220 34638 38222 34690
rect 38274 34638 38388 34690
rect 38220 34636 38388 34638
rect 38220 34626 38276 34636
rect 38332 34356 38388 34636
rect 38508 34524 38772 34534
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38508 34458 38772 34468
rect 38444 34356 38500 34366
rect 38332 34300 38444 34356
rect 38444 34290 38500 34300
rect 38220 34242 38276 34254
rect 38220 34190 38222 34242
rect 38274 34190 38276 34242
rect 38220 33684 38276 34190
rect 38220 33618 38276 33628
rect 38108 33404 39172 33460
rect 37996 33292 39060 33348
rect 37884 33236 37940 33246
rect 37884 33142 37940 33180
rect 38220 33124 38276 33134
rect 38220 33030 38276 33068
rect 38508 32956 38772 32966
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38508 32890 38772 32900
rect 37884 32676 37940 32686
rect 37884 32674 38052 32676
rect 37884 32622 37886 32674
rect 37938 32622 38052 32674
rect 37884 32620 38052 32622
rect 37884 32610 37940 32620
rect 37212 32450 37268 32462
rect 37212 32398 37214 32450
rect 37266 32398 37268 32450
rect 37212 32340 37268 32398
rect 37212 32274 37268 32284
rect 37660 32450 37716 32462
rect 37660 32398 37662 32450
rect 37714 32398 37716 32450
rect 37660 31948 37716 32398
rect 37996 31948 38052 32620
rect 38220 32562 38276 32574
rect 38220 32510 38222 32562
rect 38274 32510 38276 32562
rect 38220 32340 38276 32510
rect 38220 32274 38276 32284
rect 37324 31892 37940 31948
rect 37996 31892 38948 31948
rect 37212 31666 37268 31678
rect 37212 31614 37214 31666
rect 37266 31614 37268 31666
rect 37212 31556 37268 31614
rect 37212 31490 37268 31500
rect 37212 27188 37268 27198
rect 37212 27074 37268 27132
rect 37212 27022 37214 27074
rect 37266 27022 37268 27074
rect 37212 27010 37268 27022
rect 37100 25330 37156 25340
rect 37212 26628 37268 26638
rect 36988 24882 37044 24892
rect 37212 22484 37268 26572
rect 37324 25508 37380 31892
rect 37884 31778 37940 31892
rect 37884 31726 37886 31778
rect 37938 31726 37940 31778
rect 37884 31714 37940 31726
rect 37548 31668 37604 31678
rect 37548 31574 37604 31612
rect 38220 31556 38276 31566
rect 38220 31554 38388 31556
rect 38220 31502 38222 31554
rect 38274 31502 38388 31554
rect 38220 31500 38388 31502
rect 38220 31490 38276 31500
rect 38220 31106 38276 31118
rect 38220 31054 38222 31106
rect 38274 31054 38276 31106
rect 37884 30994 37940 31006
rect 37884 30942 37886 30994
rect 37938 30942 37940 30994
rect 37548 30884 37604 30894
rect 37884 30884 37940 30942
rect 37604 30828 37940 30884
rect 37548 30790 37604 30828
rect 38220 30324 38276 31054
rect 38332 30996 38388 31500
rect 38508 31388 38772 31398
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38508 31322 38772 31332
rect 38444 30996 38500 31006
rect 38332 30940 38444 30996
rect 38444 30930 38500 30940
rect 38220 30258 38276 30268
rect 37884 30098 37940 30110
rect 37884 30046 37886 30098
rect 37938 30046 37940 30098
rect 37660 29988 37716 29998
rect 37884 29988 37940 30046
rect 37660 29986 37940 29988
rect 37660 29934 37662 29986
rect 37714 29934 37940 29986
rect 37660 29932 37940 29934
rect 38220 29986 38276 29998
rect 38220 29934 38222 29986
rect 38274 29934 38276 29986
rect 37660 28644 37716 29932
rect 38220 29764 38276 29934
rect 38508 29820 38772 29830
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38508 29754 38772 29764
rect 38220 29698 38276 29708
rect 38220 29538 38276 29550
rect 38220 29486 38222 29538
rect 38274 29486 38276 29538
rect 37884 29428 37940 29438
rect 37884 29426 38052 29428
rect 37884 29374 37886 29426
rect 37938 29374 38052 29426
rect 37884 29372 38052 29374
rect 37884 29362 37940 29372
rect 37324 25442 37380 25452
rect 37436 28588 37716 28644
rect 37884 28642 37940 28654
rect 37884 28590 37886 28642
rect 37938 28590 37940 28642
rect 37324 25282 37380 25294
rect 37324 25230 37326 25282
rect 37378 25230 37380 25282
rect 37324 24164 37380 25230
rect 37324 24098 37380 24108
rect 37436 23380 37492 28588
rect 37660 28420 37716 28430
rect 37884 28420 37940 28590
rect 37660 28418 37940 28420
rect 37660 28366 37662 28418
rect 37714 28366 37940 28418
rect 37660 28364 37940 28366
rect 37548 27076 37604 27086
rect 37548 26962 37604 27020
rect 37548 26910 37550 26962
rect 37602 26910 37604 26962
rect 37548 26898 37604 26910
rect 37660 26628 37716 28364
rect 37884 27860 37940 27870
rect 37884 27766 37940 27804
rect 37996 27300 38052 29372
rect 38220 28980 38276 29486
rect 38220 28914 38276 28924
rect 38220 28420 38276 28430
rect 38220 28326 38276 28364
rect 38508 28252 38772 28262
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38508 28186 38772 28196
rect 38220 27970 38276 27982
rect 38220 27918 38222 27970
rect 38274 27918 38276 27970
rect 38220 27636 38276 27918
rect 38220 27570 38276 27580
rect 37884 27244 38052 27300
rect 37884 26908 37940 27244
rect 37660 26562 37716 26572
rect 37772 26852 37940 26908
rect 37996 27074 38052 27086
rect 37996 27022 37998 27074
rect 38050 27022 38052 27074
rect 37772 26404 37828 26852
rect 37548 26348 37828 26404
rect 37884 26402 37940 26414
rect 37884 26350 37886 26402
rect 37938 26350 37940 26402
rect 37548 23492 37604 26348
rect 37660 26180 37716 26190
rect 37660 26086 37716 26124
rect 37660 25732 37716 25742
rect 37884 25732 37940 26350
rect 37660 25730 37940 25732
rect 37660 25678 37662 25730
rect 37714 25678 37940 25730
rect 37660 25676 37940 25678
rect 37660 25666 37716 25676
rect 37884 25394 37940 25406
rect 37884 25342 37886 25394
rect 37938 25342 37940 25394
rect 37548 23426 37604 23436
rect 37660 25284 37716 25294
rect 37884 25284 37940 25342
rect 37660 25282 37940 25284
rect 37660 25230 37662 25282
rect 37714 25230 37940 25282
rect 37660 25228 37940 25230
rect 37436 23314 37492 23324
rect 36428 22194 36484 22204
rect 37100 22428 37268 22484
rect 30940 21858 30996 21868
rect 37100 21812 37156 22428
rect 37100 21746 37156 21756
rect 37212 22258 37268 22270
rect 37212 22206 37214 22258
rect 37266 22206 37268 22258
rect 33846 21196 34110 21206
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 33846 21130 34110 21140
rect 37212 20916 37268 22206
rect 37548 22146 37604 22158
rect 37548 22094 37550 22146
rect 37602 22094 37604 22146
rect 37548 21588 37604 22094
rect 37548 21522 37604 21532
rect 37660 21028 37716 25228
rect 37996 24948 38052 27022
rect 38220 26964 38276 26974
rect 38108 26962 38276 26964
rect 38108 26910 38222 26962
rect 38274 26910 38276 26962
rect 38108 26908 38276 26910
rect 38108 26404 38164 26908
rect 38220 26898 38276 26908
rect 38508 26684 38772 26694
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38508 26618 38772 26628
rect 38108 26338 38164 26348
rect 38220 26290 38276 26302
rect 38220 26238 38222 26290
rect 38274 26238 38276 26290
rect 38220 26180 38276 26238
rect 38220 25620 38276 26124
rect 38220 25554 38276 25564
rect 38220 25282 38276 25294
rect 38220 25230 38222 25282
rect 38274 25230 38276 25282
rect 38220 25060 38276 25230
rect 38508 25116 38772 25126
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38508 25050 38772 25060
rect 38220 24994 38276 25004
rect 37996 24892 38164 24948
rect 37996 24722 38052 24734
rect 37996 24670 37998 24722
rect 38050 24670 38052 24722
rect 37884 23828 37940 23838
rect 37772 23826 37940 23828
rect 37772 23774 37886 23826
rect 37938 23774 37940 23826
rect 37772 23772 37940 23774
rect 37772 22596 37828 23772
rect 37884 23762 37940 23772
rect 37884 23156 37940 23166
rect 37884 23062 37940 23100
rect 37772 22530 37828 22540
rect 37996 22372 38052 24670
rect 37996 22306 38052 22316
rect 37884 22258 37940 22270
rect 37884 22206 37886 22258
rect 37938 22206 37940 22258
rect 37884 22036 37940 22206
rect 37884 21970 37940 21980
rect 37660 20962 37716 20972
rect 37884 21586 37940 21598
rect 37884 21534 37886 21586
rect 37938 21534 37940 21586
rect 37212 20850 37268 20860
rect 37884 20580 37940 21534
rect 37884 20514 37940 20524
rect 37996 20802 38052 20814
rect 37996 20750 37998 20802
rect 38050 20750 38052 20802
rect 30380 20130 30548 20132
rect 30380 20078 30382 20130
rect 30434 20078 30548 20130
rect 30380 20076 30548 20078
rect 37884 20132 37940 20142
rect 30380 20066 30436 20076
rect 37884 20038 37940 20076
rect 28588 20018 28644 20030
rect 28588 19966 28590 20018
rect 28642 19966 28644 20018
rect 28420 19404 28532 19460
rect 28364 19394 28420 19404
rect 27468 19182 27470 19234
rect 27522 19182 27524 19234
rect 27244 19124 27300 19134
rect 27244 19030 27300 19068
rect 27356 19122 27412 19134
rect 27356 19070 27358 19122
rect 27410 19070 27412 19122
rect 26572 18470 26628 18508
rect 27356 18564 27412 19070
rect 26460 18452 26516 18462
rect 26460 18358 26516 18396
rect 26796 18450 26852 18462
rect 26796 18398 26798 18450
rect 26850 18398 26852 18450
rect 26796 18340 26852 18398
rect 27132 18450 27188 18462
rect 27132 18398 27134 18450
rect 27186 18398 27188 18450
rect 26796 18284 26964 18340
rect 26012 18228 26068 18238
rect 26012 18226 26516 18228
rect 26012 18174 26014 18226
rect 26066 18174 26516 18226
rect 26012 18172 26516 18174
rect 26012 18162 26068 18172
rect 26460 17666 26516 18172
rect 26460 17614 26462 17666
rect 26514 17614 26516 17666
rect 26460 17602 26516 17614
rect 26796 17444 26852 17454
rect 26684 17442 26852 17444
rect 26684 17390 26798 17442
rect 26850 17390 26852 17442
rect 26684 17388 26852 17390
rect 25340 16884 25396 16894
rect 25452 16884 25508 17052
rect 26572 17108 26628 17118
rect 25340 16882 25508 16884
rect 25340 16830 25342 16882
rect 25394 16830 25508 16882
rect 25340 16828 25508 16830
rect 25564 16994 25620 17006
rect 25564 16942 25566 16994
rect 25618 16942 25620 16994
rect 25340 16818 25396 16828
rect 25564 16772 25620 16942
rect 26460 16884 26516 16894
rect 26460 16790 26516 16828
rect 25564 16706 25620 16716
rect 26236 16772 26292 16782
rect 26236 16678 26292 16716
rect 25900 16660 25956 16670
rect 25900 16658 26180 16660
rect 25900 16606 25902 16658
rect 25954 16606 26180 16658
rect 25900 16604 26180 16606
rect 25900 16594 25956 16604
rect 25900 16212 25956 16222
rect 25116 16156 25284 16212
rect 25116 15988 25172 15998
rect 25116 15894 25172 15932
rect 25228 15764 25284 16156
rect 25900 16118 25956 16156
rect 26124 16100 26180 16604
rect 26236 16100 26292 16110
rect 26124 16098 26292 16100
rect 26124 16046 26238 16098
rect 26290 16046 26292 16098
rect 26124 16044 26292 16046
rect 26236 16034 26292 16044
rect 26572 15986 26628 17052
rect 26572 15934 26574 15986
rect 26626 15934 26628 15986
rect 26572 15922 26628 15934
rect 24892 7970 24948 7980
rect 25004 15708 25284 15764
rect 25452 15874 25508 15886
rect 25452 15822 25454 15874
rect 25506 15822 25508 15874
rect 24522 7084 24786 7094
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24522 7018 24786 7028
rect 24522 5516 24786 5526
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24522 5450 24786 5460
rect 25004 4228 25060 15708
rect 25228 15316 25284 15326
rect 25228 15222 25284 15260
rect 25228 13748 25284 13758
rect 25228 13654 25284 13692
rect 25452 11284 25508 15822
rect 25564 15426 25620 15438
rect 25564 15374 25566 15426
rect 25618 15374 25620 15426
rect 25564 14532 25620 15374
rect 25564 14466 25620 14476
rect 25452 11218 25508 11228
rect 25564 13858 25620 13870
rect 25564 13806 25566 13858
rect 25618 13806 25620 13858
rect 25004 4162 25060 4172
rect 24522 3948 24786 3958
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24522 3882 24786 3892
rect 24892 3668 24948 3678
rect 24780 3556 24836 3566
rect 24780 3462 24836 3500
rect 24556 3444 24612 3454
rect 24332 3442 24612 3444
rect 24332 3390 24558 3442
rect 24610 3390 24612 3442
rect 24332 3388 24612 3390
rect 23548 800 23604 2156
rect 24220 800 24276 3388
rect 24556 3378 24612 3388
rect 24892 800 24948 3612
rect 25564 3554 25620 13806
rect 25900 13636 25956 13646
rect 25676 4226 25732 4238
rect 25676 4174 25678 4226
rect 25730 4174 25732 4226
rect 25676 3668 25732 4174
rect 25676 3602 25732 3612
rect 25564 3502 25566 3554
rect 25618 3502 25620 3554
rect 25564 3490 25620 3502
rect 25228 3444 25284 3482
rect 25228 3378 25284 3388
rect 25900 3442 25956 13580
rect 26572 12740 26628 12750
rect 26348 4226 26404 4238
rect 26348 4174 26350 4226
rect 26402 4174 26404 4226
rect 26124 3668 26180 3678
rect 26180 3612 26292 3668
rect 26124 3602 26180 3612
rect 26236 3554 26292 3612
rect 26236 3502 26238 3554
rect 26290 3502 26292 3554
rect 26236 3490 26292 3502
rect 25900 3390 25902 3442
rect 25954 3390 25956 3442
rect 25900 3378 25956 3390
rect 26124 3444 26180 3454
rect 26124 3332 26292 3388
rect 25564 2546 25620 2558
rect 25564 2494 25566 2546
rect 25618 2494 25620 2546
rect 25564 800 25620 2494
rect 26236 800 26292 3332
rect 26348 2546 26404 4174
rect 26572 3442 26628 12684
rect 26684 6580 26740 17388
rect 26796 17378 26852 17388
rect 26908 17106 26964 18284
rect 26908 17054 26910 17106
rect 26962 17054 26964 17106
rect 26908 16884 26964 17054
rect 27132 17444 27188 18398
rect 27356 18450 27412 18508
rect 27356 18398 27358 18450
rect 27410 18398 27412 18450
rect 27356 17666 27412 18398
rect 27356 17614 27358 17666
rect 27410 17614 27412 17666
rect 27356 17602 27412 17614
rect 27468 18562 27524 19182
rect 28364 19124 28420 19134
rect 28364 19010 28420 19068
rect 28364 18958 28366 19010
rect 28418 18958 28420 19010
rect 27468 18510 27470 18562
rect 27522 18510 27524 18562
rect 27468 18452 27524 18510
rect 27468 17666 27524 18396
rect 27916 18676 27972 18686
rect 27916 18450 27972 18620
rect 28364 18564 28420 18958
rect 28364 18498 28420 18508
rect 27916 18398 27918 18450
rect 27970 18398 27972 18450
rect 27916 18386 27972 18398
rect 28476 18452 28532 19404
rect 28588 18676 28644 19966
rect 30044 20018 30100 20030
rect 30044 19966 30046 20018
rect 30098 19966 30100 20018
rect 30044 19458 30100 19966
rect 37996 20020 38052 20750
rect 38108 20692 38164 24892
rect 38220 24834 38276 24846
rect 38220 24782 38222 24834
rect 38274 24782 38276 24834
rect 38220 24276 38276 24782
rect 38220 24210 38276 24220
rect 38220 23716 38276 23726
rect 38220 23622 38276 23660
rect 38508 23548 38772 23558
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38508 23482 38772 23492
rect 38220 23266 38276 23278
rect 38220 23214 38222 23266
rect 38274 23214 38276 23266
rect 38220 22932 38276 23214
rect 38892 23268 38948 31892
rect 39004 23828 39060 33292
rect 39116 25396 39172 33404
rect 39116 25330 39172 25340
rect 39228 24836 39284 35196
rect 39116 24780 39284 24836
rect 39116 24724 39172 24780
rect 39116 24658 39172 24668
rect 39004 23762 39060 23772
rect 38892 23202 38948 23212
rect 38220 22866 38276 22876
rect 38220 22260 38276 22270
rect 38220 22166 38276 22204
rect 38508 21980 38772 21990
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38508 21914 38772 21924
rect 38220 21698 38276 21710
rect 38220 21646 38222 21698
rect 38274 21646 38276 21698
rect 38220 20916 38276 21646
rect 38220 20850 38276 20860
rect 38108 20626 38164 20636
rect 38220 20580 38276 20590
rect 38220 20578 38388 20580
rect 38220 20526 38222 20578
rect 38274 20526 38388 20578
rect 38220 20524 38388 20526
rect 38220 20514 38276 20524
rect 38332 20244 38388 20524
rect 38508 20412 38772 20422
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38508 20346 38772 20356
rect 38444 20244 38500 20254
rect 38332 20188 38444 20244
rect 38444 20178 38500 20188
rect 37996 19954 38052 19964
rect 38220 20130 38276 20142
rect 38220 20078 38222 20130
rect 38274 20078 38276 20130
rect 30044 19406 30046 19458
rect 30098 19406 30100 19458
rect 30044 19394 30100 19406
rect 30940 19906 30996 19918
rect 30940 19854 30942 19906
rect 30994 19854 30996 19906
rect 29372 19292 29764 19348
rect 29372 19234 29428 19292
rect 29372 19182 29374 19234
rect 29426 19182 29428 19234
rect 29372 19170 29428 19182
rect 29036 19124 29092 19134
rect 28700 19012 28756 19022
rect 29036 19012 29092 19068
rect 28756 18956 29092 19012
rect 28700 18946 28756 18956
rect 28588 18610 28644 18620
rect 28924 18788 28980 18798
rect 28924 18562 28980 18732
rect 28924 18510 28926 18562
rect 28978 18510 28980 18562
rect 28924 18498 28980 18510
rect 29036 18562 29092 18956
rect 29484 19122 29540 19134
rect 29484 19070 29486 19122
rect 29538 19070 29540 19122
rect 29484 19012 29540 19070
rect 29596 19124 29652 19134
rect 29596 19030 29652 19068
rect 29484 18946 29540 18956
rect 29184 18844 29448 18854
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29184 18778 29448 18788
rect 29036 18510 29038 18562
rect 29090 18510 29092 18562
rect 29036 18498 29092 18510
rect 29596 18564 29652 18574
rect 29708 18564 29764 19292
rect 30380 19234 30436 19246
rect 30380 19182 30382 19234
rect 30434 19182 30436 19234
rect 30156 19124 30212 19134
rect 29652 18508 29764 18564
rect 30044 19012 30100 19022
rect 30044 18562 30100 18956
rect 30044 18510 30046 18562
rect 30098 18510 30100 18562
rect 29596 18498 29652 18508
rect 30044 18498 30100 18510
rect 30156 18562 30212 19068
rect 30156 18510 30158 18562
rect 30210 18510 30212 18562
rect 30156 18498 30212 18510
rect 30268 18564 30324 18574
rect 28476 18396 28756 18452
rect 28364 18340 28420 18350
rect 28364 18246 28420 18284
rect 27468 17614 27470 17666
rect 27522 17614 27524 17666
rect 27468 17602 27524 17614
rect 27132 16884 27188 17388
rect 27244 17554 27300 17566
rect 27244 17502 27246 17554
rect 27298 17502 27300 17554
rect 27244 16996 27300 17502
rect 27916 17556 27972 17566
rect 28252 17556 28308 17566
rect 27916 17554 28308 17556
rect 27916 17502 27918 17554
rect 27970 17502 28254 17554
rect 28306 17502 28308 17554
rect 27916 17500 28308 17502
rect 27916 17490 27972 17500
rect 28252 17490 28308 17500
rect 28476 17444 28532 17454
rect 28364 17388 28476 17444
rect 27244 16940 27412 16996
rect 27132 16828 27300 16884
rect 26908 16818 26964 16828
rect 27020 16772 27076 16782
rect 27076 16716 27188 16772
rect 27020 16706 27076 16716
rect 27132 15316 27188 16716
rect 27244 16770 27300 16828
rect 27244 16718 27246 16770
rect 27298 16718 27300 16770
rect 27244 16706 27300 16718
rect 27132 15222 27188 15260
rect 27356 15204 27412 16940
rect 27804 16884 27860 16894
rect 28140 16884 28196 16894
rect 27804 16882 28196 16884
rect 27804 16830 27806 16882
rect 27858 16830 28142 16882
rect 28194 16830 28196 16882
rect 27804 16828 28196 16830
rect 27804 16818 27860 16828
rect 28140 16818 28196 16828
rect 27468 16772 27524 16782
rect 27468 16678 27524 16716
rect 28252 16324 28308 16334
rect 27916 16322 28308 16324
rect 27916 16270 28254 16322
rect 28306 16270 28308 16322
rect 27916 16268 28308 16270
rect 27692 15986 27748 15998
rect 27692 15934 27694 15986
rect 27746 15934 27748 15986
rect 27692 15538 27748 15934
rect 27692 15486 27694 15538
rect 27746 15486 27748 15538
rect 27692 15474 27748 15486
rect 27356 15138 27412 15148
rect 26796 15092 26852 15102
rect 26796 15090 27076 15092
rect 26796 15038 26798 15090
rect 26850 15038 27076 15090
rect 26796 15036 27076 15038
rect 26796 15026 26852 15036
rect 27020 14532 27076 15036
rect 27132 14532 27188 14542
rect 27020 14530 27188 14532
rect 27020 14478 27134 14530
rect 27186 14478 27188 14530
rect 27020 14476 27188 14478
rect 27132 14466 27188 14476
rect 27468 14420 27524 14430
rect 27468 14326 27524 14364
rect 27916 10612 27972 16268
rect 28252 16258 28308 16268
rect 28028 15876 28084 15886
rect 28364 15876 28420 17388
rect 28476 17378 28532 17388
rect 28588 17442 28644 17454
rect 28588 17390 28590 17442
rect 28642 17390 28644 17442
rect 28476 16994 28532 17006
rect 28476 16942 28478 16994
rect 28530 16942 28532 16994
rect 28476 16322 28532 16942
rect 28476 16270 28478 16322
rect 28530 16270 28532 16322
rect 28476 16258 28532 16270
rect 28476 15876 28532 15886
rect 28028 15874 28196 15876
rect 28028 15822 28030 15874
rect 28082 15822 28196 15874
rect 28028 15820 28196 15822
rect 28364 15874 28532 15876
rect 28364 15822 28478 15874
rect 28530 15822 28532 15874
rect 28364 15820 28532 15822
rect 28028 15810 28084 15820
rect 28028 15316 28084 15326
rect 28028 15222 28084 15260
rect 28140 13748 28196 15820
rect 28476 15810 28532 15820
rect 28252 15316 28308 15326
rect 28476 15316 28532 15326
rect 28252 15314 28476 15316
rect 28252 15262 28254 15314
rect 28306 15262 28476 15314
rect 28252 15260 28476 15262
rect 28252 15250 28308 15260
rect 28476 14642 28532 15260
rect 28476 14590 28478 14642
rect 28530 14590 28532 14642
rect 28476 14578 28532 14590
rect 28140 13682 28196 13692
rect 27916 10546 27972 10556
rect 28588 7364 28644 17390
rect 28700 16996 28756 18396
rect 28812 18450 28868 18462
rect 28812 18398 28814 18450
rect 28866 18398 28868 18450
rect 28812 17220 28868 18398
rect 29932 18450 29988 18462
rect 29932 18398 29934 18450
rect 29986 18398 29988 18450
rect 29932 18340 29988 18398
rect 29932 18274 29988 18284
rect 29484 18226 29540 18238
rect 29484 18174 29486 18226
rect 29538 18174 29540 18226
rect 29484 17668 29540 18174
rect 29596 17668 29652 17678
rect 29484 17666 29652 17668
rect 29484 17614 29598 17666
rect 29650 17614 29652 17666
rect 29484 17612 29652 17614
rect 29596 17602 29652 17612
rect 29260 17444 29316 17482
rect 29260 17378 29316 17388
rect 29932 17442 29988 17454
rect 29932 17390 29934 17442
rect 29986 17390 29988 17442
rect 29184 17276 29448 17286
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 28812 17164 28980 17220
rect 29184 17210 29448 17220
rect 28812 16996 28868 17006
rect 28700 16994 28868 16996
rect 28700 16942 28814 16994
rect 28866 16942 28868 16994
rect 28700 16940 28868 16942
rect 28812 16930 28868 16940
rect 28924 15204 28980 17164
rect 29148 16994 29204 17006
rect 29148 16942 29150 16994
rect 29202 16942 29204 16994
rect 29148 16660 29204 16942
rect 29820 16884 29876 16894
rect 29820 16790 29876 16828
rect 29036 16604 29148 16660
rect 29036 15316 29092 16604
rect 29148 16594 29204 16604
rect 29184 15708 29448 15718
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29184 15642 29448 15652
rect 29148 15316 29204 15326
rect 29036 15314 29204 15316
rect 29036 15262 29150 15314
rect 29202 15262 29204 15314
rect 29036 15260 29204 15262
rect 29148 15250 29204 15260
rect 29820 15316 29876 15326
rect 29820 15222 29876 15260
rect 28924 15138 28980 15148
rect 29484 15090 29540 15102
rect 29484 15038 29486 15090
rect 29538 15038 29540 15090
rect 29484 14530 29540 15038
rect 29484 14478 29486 14530
rect 29538 14478 29540 14530
rect 29484 14466 29540 14478
rect 29820 14308 29876 14318
rect 29820 14214 29876 14252
rect 29184 14140 29448 14150
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29184 14074 29448 14084
rect 29184 12572 29448 12582
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29184 12506 29448 12516
rect 29184 11004 29448 11014
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29184 10938 29448 10948
rect 29184 9436 29448 9446
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29184 9370 29448 9380
rect 29184 7868 29448 7878
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29184 7802 29448 7812
rect 28588 7298 28644 7308
rect 26684 6514 26740 6524
rect 29184 6300 29448 6310
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29184 6234 29448 6244
rect 29932 5796 29988 17390
rect 30044 16660 30100 16670
rect 30044 15314 30100 16604
rect 30044 15262 30046 15314
rect 30098 15262 30100 15314
rect 30044 15250 30100 15262
rect 30156 15316 30212 15326
rect 30268 15316 30324 18508
rect 30380 17444 30436 19182
rect 30604 19122 30660 19134
rect 30604 19070 30606 19122
rect 30658 19070 30660 19122
rect 30604 19012 30660 19070
rect 30716 19124 30772 19134
rect 30716 19030 30772 19068
rect 30604 18946 30660 18956
rect 30940 18676 30996 19854
rect 33846 19628 34110 19638
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 33846 19562 34110 19572
rect 38220 19572 38276 20078
rect 38220 19506 38276 19516
rect 37884 19236 37940 19246
rect 37884 19142 37940 19180
rect 31164 19124 31220 19134
rect 31500 19124 31556 19134
rect 31164 19122 31556 19124
rect 31164 19070 31166 19122
rect 31218 19070 31502 19122
rect 31554 19070 31556 19122
rect 31164 19068 31556 19070
rect 31164 19058 31220 19068
rect 31500 19058 31556 19068
rect 30940 18610 30996 18620
rect 31836 19010 31892 19022
rect 31836 18958 31838 19010
rect 31890 18958 31892 19010
rect 31276 18562 31332 18574
rect 31276 18510 31278 18562
rect 31330 18510 31332 18562
rect 30604 18452 30660 18462
rect 30940 18452 30996 18462
rect 30604 18450 30996 18452
rect 30604 18398 30606 18450
rect 30658 18398 30942 18450
rect 30994 18398 30996 18450
rect 30604 18396 30996 18398
rect 30604 18386 30660 18396
rect 30940 18386 30996 18396
rect 30380 17378 30436 17388
rect 30492 18340 30548 18350
rect 30492 17780 30548 18284
rect 30604 17780 30660 17790
rect 30492 17778 30660 17780
rect 30492 17726 30606 17778
rect 30658 17726 30660 17778
rect 30492 17724 30660 17726
rect 30492 16884 30548 17724
rect 30604 17714 30660 17724
rect 30492 16818 30548 16828
rect 30716 17444 30772 17454
rect 30716 16884 30772 17388
rect 31276 17108 31332 18510
rect 31724 18340 31780 18350
rect 31724 18246 31780 18284
rect 30716 16790 30772 16828
rect 31164 17052 31332 17108
rect 30380 16660 30436 16670
rect 30940 16660 30996 16670
rect 30380 16658 30548 16660
rect 30380 16606 30382 16658
rect 30434 16606 30548 16658
rect 30380 16604 30548 16606
rect 30380 16594 30436 16604
rect 30492 16098 30548 16604
rect 30940 16566 30996 16604
rect 30492 16046 30494 16098
rect 30546 16046 30548 16098
rect 30492 16034 30548 16046
rect 30828 15874 30884 15886
rect 30828 15822 30830 15874
rect 30882 15822 30884 15874
rect 30212 15260 30324 15316
rect 30380 15316 30436 15326
rect 30716 15316 30772 15326
rect 30380 15314 30772 15316
rect 30380 15262 30382 15314
rect 30434 15262 30718 15314
rect 30770 15262 30772 15314
rect 30380 15260 30772 15262
rect 30156 15250 30212 15260
rect 30380 15250 30436 15260
rect 30716 15250 30772 15260
rect 30828 10948 30884 15822
rect 31052 15426 31108 15438
rect 31052 15374 31054 15426
rect 31106 15374 31108 15426
rect 31052 12852 31108 15374
rect 31052 12786 31108 12796
rect 30828 10882 30884 10892
rect 31164 8428 31220 17052
rect 31276 16884 31332 16894
rect 31612 16884 31668 16894
rect 31276 16882 31668 16884
rect 31276 16830 31278 16882
rect 31330 16830 31614 16882
rect 31666 16830 31668 16882
rect 31276 16828 31668 16830
rect 31276 16818 31332 16828
rect 31612 16818 31668 16828
rect 31500 15316 31556 15326
rect 31500 15222 31556 15260
rect 31164 8372 31332 8428
rect 29932 5730 29988 5740
rect 31276 5124 31332 8372
rect 31276 5058 31332 5068
rect 27468 5012 27524 5022
rect 26572 3390 26574 3442
rect 26626 3390 26628 3442
rect 26572 3378 26628 3390
rect 26796 3554 26852 3566
rect 26796 3502 26798 3554
rect 26850 3502 26852 3554
rect 26348 2494 26350 2546
rect 26402 2494 26404 2546
rect 26348 2482 26404 2494
rect 26796 2546 26852 3502
rect 27468 3554 27524 4956
rect 29184 4732 29448 4742
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29184 4666 29448 4676
rect 27468 3502 27470 3554
rect 27522 3502 27524 3554
rect 27468 3490 27524 3502
rect 27244 3444 27300 3454
rect 27244 3350 27300 3388
rect 31836 3444 31892 18958
rect 32396 19010 32452 19022
rect 32396 18958 32398 19010
rect 32450 18958 32452 19010
rect 31948 16994 32004 17006
rect 31948 16942 31950 16994
rect 32002 16942 32004 16994
rect 31948 16100 32004 16942
rect 32396 16884 32452 18958
rect 38220 19012 38276 19022
rect 38220 18918 38276 18956
rect 38508 18844 38772 18854
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38508 18778 38772 18788
rect 38220 18562 38276 18574
rect 38220 18510 38222 18562
rect 38274 18510 38276 18562
rect 37884 18452 37940 18462
rect 37884 18358 37940 18396
rect 37436 18340 37492 18350
rect 33846 18060 34110 18070
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 33846 17994 34110 18004
rect 37212 17556 37268 17566
rect 37212 17462 37268 17500
rect 32396 16790 32452 16828
rect 37100 16884 37156 16894
rect 33846 16492 34110 16502
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 33846 16426 34110 16436
rect 31948 16034 32004 16044
rect 33846 14924 34110 14934
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 33846 14858 34110 14868
rect 33846 13356 34110 13366
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 33846 13290 34110 13300
rect 33846 11788 34110 11798
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 33846 11722 34110 11732
rect 33846 10220 34110 10230
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 33846 10154 34110 10164
rect 33846 8652 34110 8662
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 33846 8586 34110 8596
rect 36428 8036 36484 8046
rect 36428 7942 36484 7980
rect 33846 7084 34110 7094
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 33846 7018 34110 7028
rect 33846 5516 34110 5526
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 33846 5450 34110 5460
rect 33846 3948 34110 3958
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 33846 3882 34110 3892
rect 31836 3378 31892 3388
rect 36428 3444 36484 3454
rect 36428 3350 36484 3388
rect 36988 3442 37044 3454
rect 36988 3390 36990 3442
rect 37042 3390 37044 3442
rect 36988 3220 37044 3390
rect 37100 3444 37156 16828
rect 37212 14532 37268 14542
rect 37212 12962 37268 14476
rect 37212 12910 37214 12962
rect 37266 12910 37268 12962
rect 37212 12898 37268 12910
rect 37324 10948 37380 10958
rect 37324 9156 37380 10892
rect 37436 10388 37492 18284
rect 38220 18228 38276 18510
rect 38220 18162 38276 18172
rect 37884 17668 37940 17678
rect 37884 17574 37940 17612
rect 38220 17556 38276 17566
rect 38220 17462 38276 17500
rect 37548 17442 37604 17454
rect 37548 17390 37550 17442
rect 37602 17390 37604 17442
rect 37548 16884 37604 17390
rect 38508 17276 38772 17286
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38508 17210 38772 17220
rect 37884 16996 37940 17006
rect 37884 16902 37940 16940
rect 38220 16994 38276 17006
rect 38220 16942 38222 16994
rect 38274 16942 38276 16994
rect 37548 16818 37604 16828
rect 38220 16212 38276 16942
rect 38220 16146 38276 16156
rect 37884 16100 37940 16110
rect 37884 16006 37940 16044
rect 38220 15876 38276 15886
rect 38220 15874 38388 15876
rect 38220 15822 38222 15874
rect 38274 15822 38388 15874
rect 38220 15820 38388 15822
rect 38220 15810 38276 15820
rect 38332 15540 38388 15820
rect 38508 15708 38772 15718
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38508 15642 38772 15652
rect 38444 15540 38500 15550
rect 38332 15484 38444 15540
rect 38444 15474 38500 15484
rect 38220 15426 38276 15438
rect 38220 15374 38222 15426
rect 38274 15374 38276 15426
rect 37884 15314 37940 15326
rect 37884 15262 37886 15314
rect 37938 15262 37940 15314
rect 37772 15204 37828 15214
rect 37548 12738 37604 12750
rect 37548 12686 37550 12738
rect 37602 12686 37604 12738
rect 37548 12292 37604 12686
rect 37772 12404 37828 15148
rect 37884 14644 37940 15262
rect 37884 14578 37940 14588
rect 37996 15316 38052 15326
rect 37884 14420 37940 14430
rect 37884 14326 37940 14364
rect 37884 13748 37940 13758
rect 37884 13654 37940 13692
rect 37884 12852 37940 12862
rect 37884 12758 37940 12796
rect 37884 12404 37940 12414
rect 37772 12402 37940 12404
rect 37772 12350 37886 12402
rect 37938 12350 37940 12402
rect 37772 12348 37940 12350
rect 37884 12338 37940 12348
rect 37548 12226 37604 12236
rect 37660 12180 37716 12190
rect 37660 12086 37716 12124
rect 37884 11284 37940 11294
rect 37884 11190 37940 11228
rect 37884 10612 37940 10622
rect 37884 10518 37940 10556
rect 37436 10332 37940 10388
rect 37884 9714 37940 10332
rect 37884 9662 37886 9714
rect 37938 9662 37940 9714
rect 37884 9650 37940 9662
rect 37660 9604 37716 9614
rect 37660 9510 37716 9548
rect 37884 9156 37940 9166
rect 37324 9154 37940 9156
rect 37324 9102 37886 9154
rect 37938 9102 37940 9154
rect 37324 9100 37940 9102
rect 37884 9090 37940 9100
rect 37996 8428 38052 15260
rect 38220 14868 38276 15374
rect 38220 14802 38276 14812
rect 38220 14308 38276 14318
rect 38220 14214 38276 14252
rect 38508 14140 38772 14150
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38508 14074 38772 14084
rect 38220 13858 38276 13870
rect 38220 13806 38222 13858
rect 38274 13806 38276 13858
rect 38220 13524 38276 13806
rect 38220 13458 38276 13468
rect 38220 12852 38276 12862
rect 38220 12758 38276 12796
rect 38508 12572 38772 12582
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38508 12506 38772 12516
rect 38220 12180 38276 12190
rect 38220 11508 38276 12124
rect 38220 11442 38276 11452
rect 38220 11172 38276 11182
rect 38220 11170 38388 11172
rect 38220 11118 38222 11170
rect 38274 11118 38388 11170
rect 38220 11116 38388 11118
rect 38220 11106 38276 11116
rect 38332 10836 38388 11116
rect 38508 11004 38772 11014
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38508 10938 38772 10948
rect 38444 10836 38500 10846
rect 38332 10780 38444 10836
rect 38444 10770 38500 10780
rect 38220 10722 38276 10734
rect 38220 10670 38222 10722
rect 38274 10670 38276 10722
rect 38220 10164 38276 10670
rect 38220 10098 38276 10108
rect 38220 9714 38276 9726
rect 38220 9662 38222 9714
rect 38274 9662 38276 9714
rect 38220 9604 38276 9662
rect 38220 9538 38276 9548
rect 38508 9436 38772 9446
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38508 9370 38772 9380
rect 38220 9154 38276 9166
rect 38220 9102 38222 9154
rect 38274 9102 38276 9154
rect 38220 8820 38276 9102
rect 38220 8754 38276 8764
rect 37884 8372 38052 8428
rect 37212 8146 37268 8158
rect 37212 8094 37214 8146
rect 37266 8094 37268 8146
rect 37212 8036 37268 8094
rect 37660 8148 37716 8158
rect 37212 7970 37268 7980
rect 37548 8034 37604 8046
rect 37548 7982 37550 8034
rect 37602 7982 37604 8034
rect 37548 7476 37604 7982
rect 37660 7698 37716 8092
rect 37884 8146 37940 8372
rect 37884 8094 37886 8146
rect 37938 8094 37940 8146
rect 37884 8082 37940 8094
rect 38220 8148 38276 8158
rect 38220 8054 38276 8092
rect 38508 7868 38772 7878
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38508 7802 38772 7812
rect 37660 7646 37662 7698
rect 37714 7646 37716 7698
rect 37660 7634 37716 7646
rect 38220 7586 38276 7598
rect 38220 7534 38222 7586
rect 38274 7534 38276 7586
rect 37548 7410 37604 7420
rect 37884 7474 37940 7486
rect 37884 7422 37886 7474
rect 37938 7422 37940 7474
rect 37212 7364 37268 7374
rect 37212 7270 37268 7308
rect 37884 7364 37940 7422
rect 37884 7298 37940 7308
rect 38220 6804 38276 7534
rect 38220 6738 38276 6748
rect 37548 6580 37604 6590
rect 37884 6580 37940 6590
rect 37604 6578 37940 6580
rect 37604 6526 37886 6578
rect 37938 6526 37940 6578
rect 37604 6524 37940 6526
rect 37548 6486 37604 6524
rect 37884 6514 37940 6524
rect 38220 6466 38276 6478
rect 38220 6414 38222 6466
rect 38274 6414 38276 6466
rect 38220 6244 38276 6414
rect 38508 6300 38772 6310
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38508 6234 38772 6244
rect 38220 6178 38276 6188
rect 38220 6018 38276 6030
rect 38220 5966 38222 6018
rect 38274 5966 38276 6018
rect 37884 5906 37940 5918
rect 37884 5854 37886 5906
rect 37938 5854 37940 5906
rect 37660 5796 37716 5806
rect 37884 5796 37940 5854
rect 37716 5740 37940 5796
rect 37660 5702 37716 5740
rect 38220 5460 38276 5966
rect 38220 5394 38276 5404
rect 37548 5124 37604 5134
rect 37548 5030 37604 5068
rect 37996 5124 38052 5134
rect 37996 5030 38052 5068
rect 38220 4900 38276 4910
rect 38220 4806 38276 4844
rect 38508 4732 38772 4742
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38508 4666 38772 4676
rect 38220 4450 38276 4462
rect 38220 4398 38222 4450
rect 38274 4398 38276 4450
rect 37884 4338 37940 4350
rect 37884 4286 37886 4338
rect 37938 4286 37940 4338
rect 37660 4228 37716 4238
rect 37884 4228 37940 4286
rect 37716 4172 37940 4228
rect 37660 4134 37716 4172
rect 38220 4116 38276 4398
rect 38220 4050 38276 4060
rect 37212 3444 37268 3454
rect 37100 3442 37268 3444
rect 37100 3390 37214 3442
rect 37266 3390 37268 3442
rect 37100 3388 37268 3390
rect 37212 3378 37268 3388
rect 37548 3442 37604 3454
rect 37548 3390 37550 3442
rect 37602 3390 37604 3442
rect 37548 3220 37604 3390
rect 37884 3444 37940 3454
rect 37884 3350 37940 3388
rect 38220 3444 38276 3454
rect 38220 3350 38276 3388
rect 29184 3164 29448 3174
rect 36988 3164 37604 3220
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29184 3098 29448 3108
rect 37548 2772 37604 3164
rect 38508 3164 38772 3174
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38508 3098 38772 3108
rect 37548 2706 37604 2716
rect 26796 2494 26798 2546
rect 26850 2494 26852 2546
rect 26796 2482 26852 2494
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 22176 0 22288 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
rect 25536 0 25648 800
rect 26208 0 26320 800
<< via2 >>
rect 5874 36874 5930 36876
rect 5874 36822 5876 36874
rect 5876 36822 5928 36874
rect 5928 36822 5930 36874
rect 5874 36820 5930 36822
rect 5978 36874 6034 36876
rect 5978 36822 5980 36874
rect 5980 36822 6032 36874
rect 6032 36822 6034 36874
rect 5978 36820 6034 36822
rect 6082 36874 6138 36876
rect 6082 36822 6084 36874
rect 6084 36822 6136 36874
rect 6136 36822 6138 36874
rect 6082 36820 6138 36822
rect 15198 36874 15254 36876
rect 15198 36822 15200 36874
rect 15200 36822 15252 36874
rect 15252 36822 15254 36874
rect 15198 36820 15254 36822
rect 15302 36874 15358 36876
rect 15302 36822 15304 36874
rect 15304 36822 15356 36874
rect 15356 36822 15358 36874
rect 15302 36820 15358 36822
rect 15406 36874 15462 36876
rect 15406 36822 15408 36874
rect 15408 36822 15460 36874
rect 15460 36822 15462 36874
rect 15406 36820 15462 36822
rect 10536 36090 10592 36092
rect 10536 36038 10538 36090
rect 10538 36038 10590 36090
rect 10590 36038 10592 36090
rect 10536 36036 10592 36038
rect 10640 36090 10696 36092
rect 10640 36038 10642 36090
rect 10642 36038 10694 36090
rect 10694 36038 10696 36090
rect 10640 36036 10696 36038
rect 10744 36090 10800 36092
rect 10744 36038 10746 36090
rect 10746 36038 10798 36090
rect 10798 36038 10800 36090
rect 10744 36036 10800 36038
rect 5874 35306 5930 35308
rect 5874 35254 5876 35306
rect 5876 35254 5928 35306
rect 5928 35254 5930 35306
rect 5874 35252 5930 35254
rect 5978 35306 6034 35308
rect 5978 35254 5980 35306
rect 5980 35254 6032 35306
rect 6032 35254 6034 35306
rect 5978 35252 6034 35254
rect 6082 35306 6138 35308
rect 6082 35254 6084 35306
rect 6084 35254 6136 35306
rect 6136 35254 6138 35306
rect 6082 35252 6138 35254
rect 10536 34522 10592 34524
rect 10536 34470 10538 34522
rect 10538 34470 10590 34522
rect 10590 34470 10592 34522
rect 10536 34468 10592 34470
rect 10640 34522 10696 34524
rect 10640 34470 10642 34522
rect 10642 34470 10694 34522
rect 10694 34470 10696 34522
rect 10640 34468 10696 34470
rect 10744 34522 10800 34524
rect 10744 34470 10746 34522
rect 10746 34470 10798 34522
rect 10798 34470 10800 34522
rect 10744 34468 10800 34470
rect 5874 33738 5930 33740
rect 5874 33686 5876 33738
rect 5876 33686 5928 33738
rect 5928 33686 5930 33738
rect 5874 33684 5930 33686
rect 5978 33738 6034 33740
rect 5978 33686 5980 33738
rect 5980 33686 6032 33738
rect 6032 33686 6034 33738
rect 5978 33684 6034 33686
rect 6082 33738 6138 33740
rect 6082 33686 6084 33738
rect 6084 33686 6136 33738
rect 6136 33686 6138 33738
rect 6082 33684 6138 33686
rect 10536 32954 10592 32956
rect 10536 32902 10538 32954
rect 10538 32902 10590 32954
rect 10590 32902 10592 32954
rect 10536 32900 10592 32902
rect 10640 32954 10696 32956
rect 10640 32902 10642 32954
rect 10642 32902 10694 32954
rect 10694 32902 10696 32954
rect 10640 32900 10696 32902
rect 10744 32954 10800 32956
rect 10744 32902 10746 32954
rect 10746 32902 10798 32954
rect 10798 32902 10800 32954
rect 10744 32900 10800 32902
rect 5874 32170 5930 32172
rect 5874 32118 5876 32170
rect 5876 32118 5928 32170
rect 5928 32118 5930 32170
rect 5874 32116 5930 32118
rect 5978 32170 6034 32172
rect 5978 32118 5980 32170
rect 5980 32118 6032 32170
rect 6032 32118 6034 32170
rect 5978 32116 6034 32118
rect 6082 32170 6138 32172
rect 6082 32118 6084 32170
rect 6084 32118 6136 32170
rect 6136 32118 6138 32170
rect 6082 32116 6138 32118
rect 10536 31386 10592 31388
rect 10536 31334 10538 31386
rect 10538 31334 10590 31386
rect 10590 31334 10592 31386
rect 10536 31332 10592 31334
rect 10640 31386 10696 31388
rect 10640 31334 10642 31386
rect 10642 31334 10694 31386
rect 10694 31334 10696 31386
rect 10640 31332 10696 31334
rect 10744 31386 10800 31388
rect 10744 31334 10746 31386
rect 10746 31334 10798 31386
rect 10798 31334 10800 31386
rect 10744 31332 10800 31334
rect 5874 30602 5930 30604
rect 5874 30550 5876 30602
rect 5876 30550 5928 30602
rect 5928 30550 5930 30602
rect 5874 30548 5930 30550
rect 5978 30602 6034 30604
rect 5978 30550 5980 30602
rect 5980 30550 6032 30602
rect 6032 30550 6034 30602
rect 5978 30548 6034 30550
rect 6082 30602 6138 30604
rect 6082 30550 6084 30602
rect 6084 30550 6136 30602
rect 6136 30550 6138 30602
rect 6082 30548 6138 30550
rect 10536 29818 10592 29820
rect 10536 29766 10538 29818
rect 10538 29766 10590 29818
rect 10590 29766 10592 29818
rect 10536 29764 10592 29766
rect 10640 29818 10696 29820
rect 10640 29766 10642 29818
rect 10642 29766 10694 29818
rect 10694 29766 10696 29818
rect 10640 29764 10696 29766
rect 10744 29818 10800 29820
rect 10744 29766 10746 29818
rect 10746 29766 10798 29818
rect 10798 29766 10800 29818
rect 10744 29764 10800 29766
rect 5874 29034 5930 29036
rect 5874 28982 5876 29034
rect 5876 28982 5928 29034
rect 5928 28982 5930 29034
rect 5874 28980 5930 28982
rect 5978 29034 6034 29036
rect 5978 28982 5980 29034
rect 5980 28982 6032 29034
rect 6032 28982 6034 29034
rect 5978 28980 6034 28982
rect 6082 29034 6138 29036
rect 6082 28982 6084 29034
rect 6084 28982 6136 29034
rect 6136 28982 6138 29034
rect 6082 28980 6138 28982
rect 10536 28250 10592 28252
rect 10536 28198 10538 28250
rect 10538 28198 10590 28250
rect 10590 28198 10592 28250
rect 10536 28196 10592 28198
rect 10640 28250 10696 28252
rect 10640 28198 10642 28250
rect 10642 28198 10694 28250
rect 10694 28198 10696 28250
rect 10640 28196 10696 28198
rect 10744 28250 10800 28252
rect 10744 28198 10746 28250
rect 10746 28198 10798 28250
rect 10798 28198 10800 28250
rect 10744 28196 10800 28198
rect 5874 27466 5930 27468
rect 5874 27414 5876 27466
rect 5876 27414 5928 27466
rect 5928 27414 5930 27466
rect 5874 27412 5930 27414
rect 5978 27466 6034 27468
rect 5978 27414 5980 27466
rect 5980 27414 6032 27466
rect 6032 27414 6034 27466
rect 5978 27412 6034 27414
rect 6082 27466 6138 27468
rect 6082 27414 6084 27466
rect 6084 27414 6136 27466
rect 6136 27414 6138 27466
rect 6082 27412 6138 27414
rect 1820 26796 1876 26852
rect 1820 26236 1876 26292
rect 1708 25564 1764 25620
rect 2492 26796 2548 26852
rect 10536 26682 10592 26684
rect 10536 26630 10538 26682
rect 10538 26630 10590 26682
rect 10590 26630 10592 26682
rect 10536 26628 10592 26630
rect 10640 26682 10696 26684
rect 10640 26630 10642 26682
rect 10642 26630 10694 26682
rect 10694 26630 10696 26682
rect 10640 26628 10696 26630
rect 10744 26682 10800 26684
rect 10744 26630 10746 26682
rect 10746 26630 10798 26682
rect 10798 26630 10800 26682
rect 10744 26628 10800 26630
rect 1820 24892 1876 24948
rect 1708 24220 1764 24276
rect 1708 23714 1764 23716
rect 1708 23662 1710 23714
rect 1710 23662 1762 23714
rect 1762 23662 1764 23714
rect 1708 23660 1764 23662
rect 1708 22876 1764 22932
rect 1708 22258 1764 22260
rect 1708 22206 1710 22258
rect 1710 22206 1762 22258
rect 1762 22206 1764 22258
rect 1708 22204 1764 22206
rect 2492 24892 2548 24948
rect 2044 23154 2100 23156
rect 2044 23102 2046 23154
rect 2046 23102 2098 23154
rect 2098 23102 2100 23154
rect 2044 23100 2100 23102
rect 2044 22258 2100 22260
rect 2044 22206 2046 22258
rect 2046 22206 2098 22258
rect 2098 22206 2100 22258
rect 2044 22204 2100 22206
rect 2044 21586 2100 21588
rect 2044 21534 2046 21586
rect 2046 21534 2098 21586
rect 2098 21534 2100 21586
rect 2044 21532 2100 21534
rect 1932 21308 1988 21364
rect 1708 20860 1764 20916
rect 1708 20578 1764 20580
rect 1708 20526 1710 20578
rect 1710 20526 1762 20578
rect 1762 20526 1764 20578
rect 1708 20524 1764 20526
rect 2380 21756 2436 21812
rect 2492 20860 2548 20916
rect 2156 20636 2212 20692
rect 2044 20188 2100 20244
rect 2716 20972 2772 21028
rect 2604 20076 2660 20132
rect 2044 20018 2100 20020
rect 2044 19966 2046 20018
rect 2046 19966 2098 20018
rect 2098 19966 2100 20018
rect 2044 19964 2100 19966
rect 1708 19516 1764 19572
rect 2044 19404 2100 19460
rect 5874 25898 5930 25900
rect 5874 25846 5876 25898
rect 5876 25846 5928 25898
rect 5928 25846 5930 25898
rect 5874 25844 5930 25846
rect 5978 25898 6034 25900
rect 5978 25846 5980 25898
rect 5980 25846 6032 25898
rect 6032 25846 6034 25898
rect 5978 25844 6034 25846
rect 6082 25898 6138 25900
rect 6082 25846 6084 25898
rect 6084 25846 6136 25898
rect 6136 25846 6138 25898
rect 6082 25844 6138 25846
rect 10536 25114 10592 25116
rect 10536 25062 10538 25114
rect 10538 25062 10590 25114
rect 10590 25062 10592 25114
rect 10536 25060 10592 25062
rect 10640 25114 10696 25116
rect 10640 25062 10642 25114
rect 10642 25062 10694 25114
rect 10694 25062 10696 25114
rect 10640 25060 10696 25062
rect 10744 25114 10800 25116
rect 10744 25062 10746 25114
rect 10746 25062 10798 25114
rect 10798 25062 10800 25114
rect 10744 25060 10800 25062
rect 5874 24330 5930 24332
rect 5874 24278 5876 24330
rect 5876 24278 5928 24330
rect 5928 24278 5930 24330
rect 5874 24276 5930 24278
rect 5978 24330 6034 24332
rect 5978 24278 5980 24330
rect 5980 24278 6032 24330
rect 6032 24278 6034 24330
rect 5978 24276 6034 24278
rect 6082 24330 6138 24332
rect 6082 24278 6084 24330
rect 6084 24278 6136 24330
rect 6136 24278 6138 24330
rect 6082 24276 6138 24278
rect 15198 35306 15254 35308
rect 15198 35254 15200 35306
rect 15200 35254 15252 35306
rect 15252 35254 15254 35306
rect 15198 35252 15254 35254
rect 15302 35306 15358 35308
rect 15302 35254 15304 35306
rect 15304 35254 15356 35306
rect 15356 35254 15358 35306
rect 15302 35252 15358 35254
rect 15406 35306 15462 35308
rect 15406 35254 15408 35306
rect 15408 35254 15460 35306
rect 15460 35254 15462 35306
rect 15406 35252 15462 35254
rect 15198 33738 15254 33740
rect 15198 33686 15200 33738
rect 15200 33686 15252 33738
rect 15252 33686 15254 33738
rect 15198 33684 15254 33686
rect 15302 33738 15358 33740
rect 15302 33686 15304 33738
rect 15304 33686 15356 33738
rect 15356 33686 15358 33738
rect 15302 33684 15358 33686
rect 15406 33738 15462 33740
rect 15406 33686 15408 33738
rect 15408 33686 15460 33738
rect 15460 33686 15462 33738
rect 15406 33684 15462 33686
rect 15198 32170 15254 32172
rect 15198 32118 15200 32170
rect 15200 32118 15252 32170
rect 15252 32118 15254 32170
rect 15198 32116 15254 32118
rect 15302 32170 15358 32172
rect 15302 32118 15304 32170
rect 15304 32118 15356 32170
rect 15356 32118 15358 32170
rect 15302 32116 15358 32118
rect 15406 32170 15462 32172
rect 15406 32118 15408 32170
rect 15408 32118 15460 32170
rect 15460 32118 15462 32170
rect 15406 32116 15462 32118
rect 15198 30602 15254 30604
rect 15198 30550 15200 30602
rect 15200 30550 15252 30602
rect 15252 30550 15254 30602
rect 15198 30548 15254 30550
rect 15302 30602 15358 30604
rect 15302 30550 15304 30602
rect 15304 30550 15356 30602
rect 15356 30550 15358 30602
rect 15302 30548 15358 30550
rect 15406 30602 15462 30604
rect 15406 30550 15408 30602
rect 15408 30550 15460 30602
rect 15460 30550 15462 30602
rect 15406 30548 15462 30550
rect 15198 29034 15254 29036
rect 15198 28982 15200 29034
rect 15200 28982 15252 29034
rect 15252 28982 15254 29034
rect 15198 28980 15254 28982
rect 15302 29034 15358 29036
rect 15302 28982 15304 29034
rect 15304 28982 15356 29034
rect 15356 28982 15358 29034
rect 15302 28980 15358 28982
rect 15406 29034 15462 29036
rect 15406 28982 15408 29034
rect 15408 28982 15460 29034
rect 15460 28982 15462 29034
rect 15406 28980 15462 28982
rect 16044 35308 16100 35364
rect 15708 28588 15764 28644
rect 15198 27466 15254 27468
rect 15198 27414 15200 27466
rect 15200 27414 15252 27466
rect 15252 27414 15254 27466
rect 15198 27412 15254 27414
rect 15302 27466 15358 27468
rect 15302 27414 15304 27466
rect 15304 27414 15356 27466
rect 15356 27414 15358 27466
rect 15302 27412 15358 27414
rect 15406 27466 15462 27468
rect 15406 27414 15408 27466
rect 15408 27414 15460 27466
rect 15460 27414 15462 27466
rect 15406 27412 15462 27414
rect 15198 25898 15254 25900
rect 15198 25846 15200 25898
rect 15200 25846 15252 25898
rect 15252 25846 15254 25898
rect 15198 25844 15254 25846
rect 15302 25898 15358 25900
rect 15302 25846 15304 25898
rect 15304 25846 15356 25898
rect 15356 25846 15358 25898
rect 15302 25844 15358 25846
rect 15406 25898 15462 25900
rect 15406 25846 15408 25898
rect 15408 25846 15460 25898
rect 15460 25846 15462 25898
rect 15406 25844 15462 25846
rect 15198 24330 15254 24332
rect 15198 24278 15200 24330
rect 15200 24278 15252 24330
rect 15252 24278 15254 24330
rect 15198 24276 15254 24278
rect 15302 24330 15358 24332
rect 15302 24278 15304 24330
rect 15304 24278 15356 24330
rect 15356 24278 15358 24330
rect 15302 24276 15358 24278
rect 15406 24330 15462 24332
rect 15406 24278 15408 24330
rect 15408 24278 15460 24330
rect 15460 24278 15462 24330
rect 15406 24276 15462 24278
rect 15036 23996 15092 24052
rect 16604 24050 16660 24052
rect 16604 23998 16606 24050
rect 16606 23998 16658 24050
rect 16658 23998 16660 24050
rect 16604 23996 16660 23998
rect 17276 35308 17332 35364
rect 17612 28588 17668 28644
rect 17612 24444 17668 24500
rect 10536 23546 10592 23548
rect 10536 23494 10538 23546
rect 10538 23494 10590 23546
rect 10590 23494 10592 23546
rect 10536 23492 10592 23494
rect 10640 23546 10696 23548
rect 10640 23494 10642 23546
rect 10642 23494 10694 23546
rect 10694 23494 10696 23546
rect 10640 23492 10696 23494
rect 10744 23546 10800 23548
rect 10744 23494 10746 23546
rect 10746 23494 10798 23546
rect 10798 23494 10800 23546
rect 10744 23492 10800 23494
rect 15596 23100 15652 23156
rect 5874 22762 5930 22764
rect 5874 22710 5876 22762
rect 5876 22710 5928 22762
rect 5928 22710 5930 22762
rect 5874 22708 5930 22710
rect 5978 22762 6034 22764
rect 5978 22710 5980 22762
rect 5980 22710 6032 22762
rect 6032 22710 6034 22762
rect 5978 22708 6034 22710
rect 6082 22762 6138 22764
rect 6082 22710 6084 22762
rect 6084 22710 6136 22762
rect 6136 22710 6138 22762
rect 6082 22708 6138 22710
rect 15198 22762 15254 22764
rect 15198 22710 15200 22762
rect 15200 22710 15252 22762
rect 15252 22710 15254 22762
rect 15198 22708 15254 22710
rect 15302 22762 15358 22764
rect 15302 22710 15304 22762
rect 15304 22710 15356 22762
rect 15356 22710 15358 22762
rect 15302 22708 15358 22710
rect 15406 22762 15462 22764
rect 15406 22710 15408 22762
rect 15408 22710 15460 22762
rect 15460 22710 15462 22762
rect 15406 22708 15462 22710
rect 14700 22204 14756 22260
rect 10536 21978 10592 21980
rect 10536 21926 10538 21978
rect 10538 21926 10590 21978
rect 10590 21926 10592 21978
rect 10536 21924 10592 21926
rect 10640 21978 10696 21980
rect 10640 21926 10642 21978
rect 10642 21926 10694 21978
rect 10694 21926 10696 21978
rect 10640 21924 10696 21926
rect 10744 21978 10800 21980
rect 10744 21926 10746 21978
rect 10746 21926 10798 21978
rect 10798 21926 10800 21978
rect 10744 21924 10800 21926
rect 17052 23884 17108 23940
rect 17388 24050 17444 24052
rect 17388 23998 17390 24050
rect 17390 23998 17442 24050
rect 17442 23998 17444 24050
rect 17388 23996 17444 23998
rect 16716 22540 16772 22596
rect 17164 22428 17220 22484
rect 17388 22540 17444 22596
rect 17612 22370 17668 22372
rect 17612 22318 17614 22370
rect 17614 22318 17666 22370
rect 17666 22318 17668 22370
rect 17612 22316 17668 22318
rect 18508 33964 18564 34020
rect 19068 31948 19124 32004
rect 19068 30044 19124 30100
rect 19292 33964 19348 34020
rect 19292 25452 19348 25508
rect 19180 25282 19236 25284
rect 19180 25230 19182 25282
rect 19182 25230 19234 25282
rect 19234 25230 19236 25282
rect 19180 25228 19236 25230
rect 19404 25228 19460 25284
rect 18396 24780 18452 24836
rect 19860 36090 19916 36092
rect 19860 36038 19862 36090
rect 19862 36038 19914 36090
rect 19914 36038 19916 36090
rect 19860 36036 19916 36038
rect 19964 36090 20020 36092
rect 19964 36038 19966 36090
rect 19966 36038 20018 36090
rect 20018 36038 20020 36090
rect 19964 36036 20020 36038
rect 20068 36090 20124 36092
rect 20068 36038 20070 36090
rect 20070 36038 20122 36090
rect 20122 36038 20124 36090
rect 20068 36036 20124 36038
rect 19860 34522 19916 34524
rect 19860 34470 19862 34522
rect 19862 34470 19914 34522
rect 19914 34470 19916 34522
rect 19860 34468 19916 34470
rect 19964 34522 20020 34524
rect 19964 34470 19966 34522
rect 19966 34470 20018 34522
rect 20018 34470 20020 34522
rect 19964 34468 20020 34470
rect 20068 34522 20124 34524
rect 20068 34470 20070 34522
rect 20070 34470 20122 34522
rect 20122 34470 20124 34522
rect 20068 34468 20124 34470
rect 19860 32954 19916 32956
rect 19860 32902 19862 32954
rect 19862 32902 19914 32954
rect 19914 32902 19916 32954
rect 19860 32900 19916 32902
rect 19964 32954 20020 32956
rect 19964 32902 19966 32954
rect 19966 32902 20018 32954
rect 20018 32902 20020 32954
rect 19964 32900 20020 32902
rect 20068 32954 20124 32956
rect 20068 32902 20070 32954
rect 20070 32902 20122 32954
rect 20122 32902 20124 32954
rect 20068 32900 20124 32902
rect 19740 31948 19796 32004
rect 19860 31386 19916 31388
rect 19860 31334 19862 31386
rect 19862 31334 19914 31386
rect 19914 31334 19916 31386
rect 19860 31332 19916 31334
rect 19964 31386 20020 31388
rect 19964 31334 19966 31386
rect 19966 31334 20018 31386
rect 20018 31334 20020 31386
rect 19964 31332 20020 31334
rect 20068 31386 20124 31388
rect 20068 31334 20070 31386
rect 20070 31334 20122 31386
rect 20122 31334 20124 31386
rect 20068 31332 20124 31334
rect 20188 30044 20244 30100
rect 19860 29818 19916 29820
rect 19860 29766 19862 29818
rect 19862 29766 19914 29818
rect 19914 29766 19916 29818
rect 19860 29764 19916 29766
rect 19964 29818 20020 29820
rect 19964 29766 19966 29818
rect 19966 29766 20018 29818
rect 20018 29766 20020 29818
rect 19964 29764 20020 29766
rect 20068 29818 20124 29820
rect 20068 29766 20070 29818
rect 20070 29766 20122 29818
rect 20122 29766 20124 29818
rect 20068 29764 20124 29766
rect 19860 28250 19916 28252
rect 19860 28198 19862 28250
rect 19862 28198 19914 28250
rect 19914 28198 19916 28250
rect 19860 28196 19916 28198
rect 19964 28250 20020 28252
rect 19964 28198 19966 28250
rect 19966 28198 20018 28250
rect 20018 28198 20020 28250
rect 19964 28196 20020 28198
rect 20068 28250 20124 28252
rect 20068 28198 20070 28250
rect 20070 28198 20122 28250
rect 20122 28198 20124 28250
rect 20068 28196 20124 28198
rect 19860 26682 19916 26684
rect 19860 26630 19862 26682
rect 19862 26630 19914 26682
rect 19914 26630 19916 26682
rect 19860 26628 19916 26630
rect 19964 26682 20020 26684
rect 19964 26630 19966 26682
rect 19966 26630 20018 26682
rect 20018 26630 20020 26682
rect 19964 26628 20020 26630
rect 20068 26682 20124 26684
rect 20068 26630 20070 26682
rect 20070 26630 20122 26682
rect 20122 26630 20124 26682
rect 20068 26628 20124 26630
rect 19852 25506 19908 25508
rect 19852 25454 19854 25506
rect 19854 25454 19906 25506
rect 19906 25454 19908 25506
rect 19852 25452 19908 25454
rect 19740 25228 19796 25284
rect 18620 24498 18676 24500
rect 18620 24446 18622 24498
rect 18622 24446 18674 24498
rect 18674 24446 18676 24498
rect 18620 24444 18676 24446
rect 19516 24498 19572 24500
rect 19516 24446 19518 24498
rect 19518 24446 19570 24498
rect 19570 24446 19572 24498
rect 19516 24444 19572 24446
rect 18844 23938 18900 23940
rect 18844 23886 18846 23938
rect 18846 23886 18898 23938
rect 18898 23886 18900 23938
rect 18844 23884 18900 23886
rect 18844 22482 18900 22484
rect 18844 22430 18846 22482
rect 18846 22430 18898 22482
rect 18898 22430 18900 22482
rect 18844 22428 18900 22430
rect 18620 22370 18676 22372
rect 18620 22318 18622 22370
rect 18622 22318 18674 22370
rect 18674 22318 18676 22370
rect 18620 22316 18676 22318
rect 12348 21698 12404 21700
rect 12348 21646 12350 21698
rect 12350 21646 12402 21698
rect 12402 21646 12404 21698
rect 12348 21644 12404 21646
rect 10332 21308 10388 21364
rect 5874 21194 5930 21196
rect 5874 21142 5876 21194
rect 5876 21142 5928 21194
rect 5928 21142 5930 21194
rect 5874 21140 5930 21142
rect 5978 21194 6034 21196
rect 5978 21142 5980 21194
rect 5980 21142 6032 21194
rect 6032 21142 6034 21194
rect 5978 21140 6034 21142
rect 6082 21194 6138 21196
rect 6082 21142 6084 21194
rect 6084 21142 6136 21194
rect 6136 21142 6138 21194
rect 6082 21140 6138 21142
rect 15198 21194 15254 21196
rect 15198 21142 15200 21194
rect 15200 21142 15252 21194
rect 15252 21142 15254 21194
rect 15198 21140 15254 21142
rect 15302 21194 15358 21196
rect 15302 21142 15304 21194
rect 15304 21142 15356 21194
rect 15356 21142 15358 21194
rect 15302 21140 15358 21142
rect 15406 21194 15462 21196
rect 15406 21142 15408 21194
rect 15408 21142 15460 21194
rect 15460 21142 15462 21194
rect 15406 21140 15462 21142
rect 11116 20690 11172 20692
rect 11116 20638 11118 20690
rect 11118 20638 11170 20690
rect 11170 20638 11172 20690
rect 11116 20636 11172 20638
rect 10780 20578 10836 20580
rect 10780 20526 10782 20578
rect 10782 20526 10834 20578
rect 10834 20526 10836 20578
rect 10780 20524 10836 20526
rect 5874 19626 5930 19628
rect 5874 19574 5876 19626
rect 5876 19574 5928 19626
rect 5928 19574 5930 19626
rect 5874 19572 5930 19574
rect 5978 19626 6034 19628
rect 5978 19574 5980 19626
rect 5980 19574 6032 19626
rect 6032 19574 6034 19626
rect 5978 19572 6034 19574
rect 6082 19626 6138 19628
rect 6082 19574 6084 19626
rect 6084 19574 6136 19626
rect 6136 19574 6138 19626
rect 6082 19572 6138 19574
rect 2828 19180 2884 19236
rect 1708 19010 1764 19012
rect 1708 18958 1710 19010
rect 1710 18958 1762 19010
rect 1762 18958 1764 19010
rect 1708 18956 1764 18958
rect 2044 18450 2100 18452
rect 2044 18398 2046 18450
rect 2046 18398 2098 18450
rect 2098 18398 2100 18450
rect 2044 18396 2100 18398
rect 10536 20410 10592 20412
rect 10536 20358 10538 20410
rect 10538 20358 10590 20410
rect 10590 20358 10592 20410
rect 10536 20356 10592 20358
rect 10640 20410 10696 20412
rect 10640 20358 10642 20410
rect 10642 20358 10694 20410
rect 10694 20358 10696 20410
rect 10640 20356 10696 20358
rect 10744 20410 10800 20412
rect 10744 20358 10746 20410
rect 10746 20358 10798 20410
rect 10798 20358 10800 20410
rect 10744 20356 10800 20358
rect 11788 20524 11844 20580
rect 11788 20188 11844 20244
rect 10780 20130 10836 20132
rect 10780 20078 10782 20130
rect 10782 20078 10834 20130
rect 10834 20078 10836 20130
rect 10780 20076 10836 20078
rect 11676 20076 11732 20132
rect 10536 18842 10592 18844
rect 10536 18790 10538 18842
rect 10538 18790 10590 18842
rect 10590 18790 10592 18842
rect 10536 18788 10592 18790
rect 10640 18842 10696 18844
rect 10640 18790 10642 18842
rect 10642 18790 10694 18842
rect 10694 18790 10696 18842
rect 10640 18788 10696 18790
rect 10744 18842 10800 18844
rect 10744 18790 10746 18842
rect 10746 18790 10798 18842
rect 10798 18790 10800 18842
rect 10744 18788 10800 18790
rect 1708 18172 1764 18228
rect 5874 18058 5930 18060
rect 5874 18006 5876 18058
rect 5876 18006 5928 18058
rect 5928 18006 5930 18058
rect 5874 18004 5930 18006
rect 5978 18058 6034 18060
rect 5978 18006 5980 18058
rect 5980 18006 6032 18058
rect 6032 18006 6034 18058
rect 5978 18004 6034 18006
rect 6082 18058 6138 18060
rect 6082 18006 6084 18058
rect 6084 18006 6136 18058
rect 6136 18006 6138 18058
rect 6082 18004 6138 18006
rect 2044 17836 2100 17892
rect 1708 17554 1764 17556
rect 1708 17502 1710 17554
rect 1710 17502 1762 17554
rect 1762 17502 1764 17554
rect 1708 17500 1764 17502
rect 1708 16156 1764 16212
rect 2716 17666 2772 17668
rect 2716 17614 2718 17666
rect 2718 17614 2770 17666
rect 2770 17614 2772 17666
rect 2716 17612 2772 17614
rect 10892 17612 10948 17668
rect 3164 17554 3220 17556
rect 3164 17502 3166 17554
rect 3166 17502 3218 17554
rect 3218 17502 3220 17554
rect 3164 17500 3220 17502
rect 2044 17442 2100 17444
rect 2044 17390 2046 17442
rect 2046 17390 2098 17442
rect 2098 17390 2100 17442
rect 2044 17388 2100 17390
rect 11676 19292 11732 19348
rect 11900 19794 11956 19796
rect 11900 19742 11902 19794
rect 11902 19742 11954 19794
rect 11954 19742 11956 19794
rect 11900 19740 11956 19742
rect 12012 20524 12068 20580
rect 14700 20748 14756 20804
rect 13580 20578 13636 20580
rect 13580 20526 13582 20578
rect 13582 20526 13634 20578
rect 13634 20526 13636 20578
rect 13580 20524 13636 20526
rect 14140 20690 14196 20692
rect 14140 20638 14142 20690
rect 14142 20638 14194 20690
rect 14194 20638 14196 20690
rect 14140 20636 14196 20638
rect 12124 20076 12180 20132
rect 14252 20130 14308 20132
rect 14252 20078 14254 20130
rect 14254 20078 14306 20130
rect 14306 20078 14308 20130
rect 14252 20076 14308 20078
rect 16828 20972 16884 21028
rect 15596 20748 15652 20804
rect 15260 20636 15316 20692
rect 16268 20690 16324 20692
rect 16268 20638 16270 20690
rect 16270 20638 16322 20690
rect 16322 20638 16324 20690
rect 16268 20636 16324 20638
rect 15372 20188 15428 20244
rect 17948 20860 18004 20916
rect 16156 20242 16212 20244
rect 16156 20190 16158 20242
rect 16158 20190 16210 20242
rect 16210 20190 16212 20242
rect 16156 20188 16212 20190
rect 19180 21586 19236 21588
rect 19180 21534 19182 21586
rect 19182 21534 19234 21586
rect 19234 21534 19236 21586
rect 19180 21532 19236 21534
rect 18844 20690 18900 20692
rect 18844 20638 18846 20690
rect 18846 20638 18898 20690
rect 18898 20638 18900 20690
rect 18844 20636 18900 20638
rect 19068 20524 19124 20580
rect 19860 25114 19916 25116
rect 19860 25062 19862 25114
rect 19862 25062 19914 25114
rect 19914 25062 19916 25114
rect 19860 25060 19916 25062
rect 19964 25114 20020 25116
rect 19964 25062 19966 25114
rect 19966 25062 20018 25114
rect 20018 25062 20020 25114
rect 19964 25060 20020 25062
rect 20068 25114 20124 25116
rect 20068 25062 20070 25114
rect 20070 25062 20122 25114
rect 20122 25062 20124 25114
rect 20068 25060 20124 25062
rect 19852 24722 19908 24724
rect 19852 24670 19854 24722
rect 19854 24670 19906 24722
rect 19906 24670 19908 24722
rect 19852 24668 19908 24670
rect 20300 24780 20356 24836
rect 19860 23546 19916 23548
rect 19860 23494 19862 23546
rect 19862 23494 19914 23546
rect 19914 23494 19916 23546
rect 19860 23492 19916 23494
rect 19964 23546 20020 23548
rect 19964 23494 19966 23546
rect 19966 23494 20018 23546
rect 20018 23494 20020 23546
rect 19964 23492 20020 23494
rect 20068 23546 20124 23548
rect 20068 23494 20070 23546
rect 20070 23494 20122 23546
rect 20122 23494 20124 23546
rect 20068 23492 20124 23494
rect 19740 23266 19796 23268
rect 19740 23214 19742 23266
rect 19742 23214 19794 23266
rect 19794 23214 19796 23266
rect 19740 23212 19796 23214
rect 19628 22370 19684 22372
rect 19628 22318 19630 22370
rect 19630 22318 19682 22370
rect 19682 22318 19684 22370
rect 19628 22316 19684 22318
rect 19964 22540 20020 22596
rect 19860 21978 19916 21980
rect 19860 21926 19862 21978
rect 19862 21926 19914 21978
rect 19914 21926 19916 21978
rect 19860 21924 19916 21926
rect 19964 21978 20020 21980
rect 19964 21926 19966 21978
rect 19966 21926 20018 21978
rect 20018 21926 20020 21978
rect 19964 21924 20020 21926
rect 20068 21978 20124 21980
rect 20068 21926 20070 21978
rect 20070 21926 20122 21978
rect 20122 21926 20124 21978
rect 20068 21924 20124 21926
rect 19740 21474 19796 21476
rect 19740 21422 19742 21474
rect 19742 21422 19794 21474
rect 19794 21422 19796 21474
rect 19740 21420 19796 21422
rect 20524 24722 20580 24724
rect 20524 24670 20526 24722
rect 20526 24670 20578 24722
rect 20578 24670 20580 24722
rect 20524 24668 20580 24670
rect 20636 23884 20692 23940
rect 20636 23548 20692 23604
rect 20412 23100 20468 23156
rect 20300 22540 20356 22596
rect 20300 22204 20356 22260
rect 21420 26460 21476 26516
rect 22092 25506 22148 25508
rect 22092 25454 22094 25506
rect 22094 25454 22146 25506
rect 22146 25454 22148 25506
rect 22092 25452 22148 25454
rect 21420 25228 21476 25284
rect 21084 24834 21140 24836
rect 21084 24782 21086 24834
rect 21086 24782 21138 24834
rect 21138 24782 21140 24834
rect 21084 24780 21140 24782
rect 20860 23324 20916 23380
rect 21084 23266 21140 23268
rect 21084 23214 21086 23266
rect 21086 23214 21138 23266
rect 21138 23214 21140 23266
rect 21084 23212 21140 23214
rect 21756 25340 21812 25396
rect 22316 26514 22372 26516
rect 22316 26462 22318 26514
rect 22318 26462 22370 26514
rect 22370 26462 22372 26514
rect 22316 26460 22372 26462
rect 22428 25394 22484 25396
rect 22428 25342 22430 25394
rect 22430 25342 22482 25394
rect 22482 25342 22484 25394
rect 22428 25340 22484 25342
rect 24522 36874 24578 36876
rect 24522 36822 24524 36874
rect 24524 36822 24576 36874
rect 24576 36822 24578 36874
rect 24522 36820 24578 36822
rect 24626 36874 24682 36876
rect 24626 36822 24628 36874
rect 24628 36822 24680 36874
rect 24680 36822 24682 36874
rect 24626 36820 24682 36822
rect 24730 36874 24786 36876
rect 24730 36822 24732 36874
rect 24732 36822 24784 36874
rect 24784 36822 24786 36874
rect 24730 36820 24786 36822
rect 24220 36652 24276 36708
rect 23324 36316 23380 36372
rect 23100 25506 23156 25508
rect 23100 25454 23102 25506
rect 23102 25454 23154 25506
rect 23154 25454 23156 25506
rect 23100 25452 23156 25454
rect 33846 36874 33902 36876
rect 33846 36822 33848 36874
rect 33848 36822 33900 36874
rect 33900 36822 33902 36874
rect 33846 36820 33902 36822
rect 33950 36874 34006 36876
rect 33950 36822 33952 36874
rect 33952 36822 34004 36874
rect 34004 36822 34006 36874
rect 33950 36820 34006 36822
rect 34054 36874 34110 36876
rect 34054 36822 34056 36874
rect 34056 36822 34108 36874
rect 34108 36822 34110 36874
rect 34054 36820 34110 36822
rect 37548 36876 37604 36932
rect 24892 36428 24948 36484
rect 25228 36652 25284 36708
rect 25676 36428 25732 36484
rect 25564 36370 25620 36372
rect 25564 36318 25566 36370
rect 25566 36318 25618 36370
rect 25618 36318 25620 36370
rect 25564 36316 25620 36318
rect 26124 36482 26180 36484
rect 26124 36430 26126 36482
rect 26126 36430 26178 36482
rect 26178 36430 26180 36482
rect 26124 36428 26180 36430
rect 23996 31500 24052 31556
rect 22204 24780 22260 24836
rect 22764 24108 22820 24164
rect 21196 23100 21252 23156
rect 20412 21532 20468 21588
rect 20300 21420 20356 21476
rect 20188 20748 20244 20804
rect 19628 20578 19684 20580
rect 19628 20526 19630 20578
rect 19630 20526 19682 20578
rect 19682 20526 19684 20578
rect 19628 20524 19684 20526
rect 19860 20410 19916 20412
rect 19860 20358 19862 20410
rect 19862 20358 19914 20410
rect 19914 20358 19916 20410
rect 19860 20356 19916 20358
rect 19964 20410 20020 20412
rect 19964 20358 19966 20410
rect 19966 20358 20018 20410
rect 20018 20358 20020 20410
rect 19964 20356 20020 20358
rect 20068 20410 20124 20412
rect 20068 20358 20070 20410
rect 20070 20358 20122 20410
rect 20122 20358 20124 20410
rect 20068 20356 20124 20358
rect 13580 19906 13636 19908
rect 13580 19854 13582 19906
rect 13582 19854 13634 19906
rect 13634 19854 13636 19906
rect 13580 19852 13636 19854
rect 12796 19794 12852 19796
rect 12796 19742 12798 19794
rect 12798 19742 12850 19794
rect 12850 19742 12852 19794
rect 12796 19740 12852 19742
rect 12124 18450 12180 18452
rect 12124 18398 12126 18450
rect 12126 18398 12178 18450
rect 12178 18398 12180 18450
rect 12124 18396 12180 18398
rect 11900 18226 11956 18228
rect 11900 18174 11902 18226
rect 11902 18174 11954 18226
rect 11954 18174 11956 18226
rect 11900 18172 11956 18174
rect 12796 18226 12852 18228
rect 12796 18174 12798 18226
rect 12798 18174 12850 18226
rect 12850 18174 12852 18226
rect 12796 18172 12852 18174
rect 15820 19964 15876 20020
rect 14924 19852 14980 19908
rect 15198 19626 15254 19628
rect 15198 19574 15200 19626
rect 15200 19574 15252 19626
rect 15252 19574 15254 19626
rect 15198 19572 15254 19574
rect 15302 19626 15358 19628
rect 15302 19574 15304 19626
rect 15304 19574 15356 19626
rect 15356 19574 15358 19626
rect 15302 19572 15358 19574
rect 15406 19626 15462 19628
rect 15406 19574 15408 19626
rect 15408 19574 15460 19626
rect 15460 19574 15462 19626
rect 15406 19572 15462 19574
rect 13580 19346 13636 19348
rect 13580 19294 13582 19346
rect 13582 19294 13634 19346
rect 13634 19294 13636 19346
rect 13580 19292 13636 19294
rect 14028 19292 14084 19348
rect 14924 19180 14980 19236
rect 14588 19068 14644 19124
rect 13804 18396 13860 18452
rect 12572 17836 12628 17892
rect 12908 17554 12964 17556
rect 12908 17502 12910 17554
rect 12910 17502 12962 17554
rect 12962 17502 12964 17554
rect 12908 17500 12964 17502
rect 10536 17274 10592 17276
rect 10536 17222 10538 17274
rect 10538 17222 10590 17274
rect 10590 17222 10592 17274
rect 10536 17220 10592 17222
rect 10640 17274 10696 17276
rect 10640 17222 10642 17274
rect 10642 17222 10694 17274
rect 10694 17222 10696 17274
rect 10640 17220 10696 17222
rect 10744 17274 10800 17276
rect 10744 17222 10746 17274
rect 10746 17222 10798 17274
rect 10798 17222 10800 17274
rect 10744 17220 10800 17222
rect 2380 17052 2436 17108
rect 2268 16940 2324 16996
rect 2044 16882 2100 16884
rect 2044 16830 2046 16882
rect 2046 16830 2098 16882
rect 2098 16830 2100 16882
rect 2044 16828 2100 16830
rect 1708 15874 1764 15876
rect 1708 15822 1710 15874
rect 1710 15822 1762 15874
rect 1762 15822 1764 15874
rect 1708 15820 1764 15822
rect 2044 15314 2100 15316
rect 2044 15262 2046 15314
rect 2046 15262 2098 15314
rect 2098 15262 2100 15314
rect 2044 15260 2100 15262
rect 1708 14812 1764 14868
rect 2156 15148 2212 15204
rect 2044 14306 2100 14308
rect 2044 14254 2046 14306
rect 2046 14254 2098 14306
rect 2098 14254 2100 14306
rect 2044 14252 2100 14254
rect 1708 14140 1764 14196
rect 1708 13468 1764 13524
rect 1708 12850 1764 12852
rect 1708 12798 1710 12850
rect 1710 12798 1762 12850
rect 1762 12798 1764 12850
rect 1708 12796 1764 12798
rect 11340 16940 11396 16996
rect 5874 16490 5930 16492
rect 5874 16438 5876 16490
rect 5876 16438 5928 16490
rect 5928 16438 5930 16490
rect 5874 16436 5930 16438
rect 5978 16490 6034 16492
rect 5978 16438 5980 16490
rect 5980 16438 6032 16490
rect 6032 16438 6034 16490
rect 5978 16436 6034 16438
rect 6082 16490 6138 16492
rect 6082 16438 6084 16490
rect 6084 16438 6136 16490
rect 6136 16438 6138 16490
rect 6082 16436 6138 16438
rect 10536 15706 10592 15708
rect 10536 15654 10538 15706
rect 10538 15654 10590 15706
rect 10590 15654 10592 15706
rect 10536 15652 10592 15654
rect 10640 15706 10696 15708
rect 10640 15654 10642 15706
rect 10642 15654 10694 15706
rect 10694 15654 10696 15706
rect 10640 15652 10696 15654
rect 10744 15706 10800 15708
rect 10744 15654 10746 15706
rect 10746 15654 10798 15706
rect 10798 15654 10800 15706
rect 10744 15652 10800 15654
rect 14028 18450 14084 18452
rect 14028 18398 14030 18450
rect 14030 18398 14082 18450
rect 14082 18398 14084 18450
rect 14028 18396 14084 18398
rect 13692 17500 13748 17556
rect 12908 16994 12964 16996
rect 12908 16942 12910 16994
rect 12910 16942 12962 16994
rect 12962 16942 12964 16994
rect 12908 16940 12964 16942
rect 12572 16828 12628 16884
rect 15932 19122 15988 19124
rect 15932 19070 15934 19122
rect 15934 19070 15986 19122
rect 15986 19070 15988 19122
rect 15932 19068 15988 19070
rect 15820 18508 15876 18564
rect 15372 18396 15428 18452
rect 14140 17836 14196 17892
rect 14924 18284 14980 18340
rect 14588 17666 14644 17668
rect 14588 17614 14590 17666
rect 14590 17614 14642 17666
rect 14642 17614 14644 17666
rect 14588 17612 14644 17614
rect 15198 18058 15254 18060
rect 15198 18006 15200 18058
rect 15200 18006 15252 18058
rect 15252 18006 15254 18058
rect 15198 18004 15254 18006
rect 15302 18058 15358 18060
rect 15302 18006 15304 18058
rect 15304 18006 15356 18058
rect 15356 18006 15358 18058
rect 15302 18004 15358 18006
rect 15406 18058 15462 18060
rect 15406 18006 15408 18058
rect 15408 18006 15460 18058
rect 15460 18006 15462 18058
rect 15406 18004 15462 18006
rect 15148 17666 15204 17668
rect 15148 17614 15150 17666
rect 15150 17614 15202 17666
rect 15202 17614 15204 17666
rect 15148 17612 15204 17614
rect 15036 17388 15092 17444
rect 14364 16994 14420 16996
rect 14364 16942 14366 16994
rect 14366 16942 14418 16994
rect 14418 16942 14420 16994
rect 14364 16940 14420 16942
rect 15198 16490 15254 16492
rect 15198 16438 15200 16490
rect 15200 16438 15252 16490
rect 15252 16438 15254 16490
rect 15198 16436 15254 16438
rect 15302 16490 15358 16492
rect 15302 16438 15304 16490
rect 15304 16438 15356 16490
rect 15356 16438 15358 16490
rect 15302 16436 15358 16438
rect 15406 16490 15462 16492
rect 15406 16438 15408 16490
rect 15408 16438 15460 16490
rect 15460 16438 15462 16490
rect 15406 16436 15462 16438
rect 14252 15932 14308 15988
rect 12124 15260 12180 15316
rect 5874 14922 5930 14924
rect 5874 14870 5876 14922
rect 5876 14870 5928 14922
rect 5928 14870 5930 14922
rect 5874 14868 5930 14870
rect 5978 14922 6034 14924
rect 5978 14870 5980 14922
rect 5980 14870 6032 14922
rect 6032 14870 6034 14922
rect 5978 14868 6034 14870
rect 6082 14922 6138 14924
rect 6082 14870 6084 14922
rect 6084 14870 6136 14922
rect 6136 14870 6138 14922
rect 6082 14868 6138 14870
rect 14700 15202 14756 15204
rect 14700 15150 14702 15202
rect 14702 15150 14754 15202
rect 14754 15150 14756 15202
rect 14700 15148 14756 15150
rect 15596 15148 15652 15204
rect 15198 14922 15254 14924
rect 15198 14870 15200 14922
rect 15200 14870 15252 14922
rect 15252 14870 15254 14922
rect 15198 14868 15254 14870
rect 15302 14922 15358 14924
rect 15302 14870 15304 14922
rect 15304 14870 15356 14922
rect 15356 14870 15358 14922
rect 15302 14868 15358 14870
rect 15406 14922 15462 14924
rect 15406 14870 15408 14922
rect 15408 14870 15460 14922
rect 15460 14870 15462 14922
rect 15406 14868 15462 14870
rect 15708 14476 15764 14532
rect 14924 14252 14980 14308
rect 15484 14252 15540 14308
rect 2492 14140 2548 14196
rect 10536 14138 10592 14140
rect 10536 14086 10538 14138
rect 10538 14086 10590 14138
rect 10590 14086 10592 14138
rect 10536 14084 10592 14086
rect 10640 14138 10696 14140
rect 10640 14086 10642 14138
rect 10642 14086 10694 14138
rect 10694 14086 10696 14138
rect 10640 14084 10696 14086
rect 10744 14138 10800 14140
rect 10744 14086 10746 14138
rect 10746 14086 10798 14138
rect 10798 14086 10800 14138
rect 10744 14084 10800 14086
rect 2492 13468 2548 13524
rect 14812 13580 14868 13636
rect 5874 13354 5930 13356
rect 5874 13302 5876 13354
rect 5876 13302 5928 13354
rect 5928 13302 5930 13354
rect 5874 13300 5930 13302
rect 5978 13354 6034 13356
rect 5978 13302 5980 13354
rect 5980 13302 6032 13354
rect 6032 13302 6034 13354
rect 5978 13300 6034 13302
rect 6082 13354 6138 13356
rect 6082 13302 6084 13354
rect 6084 13302 6136 13354
rect 6136 13302 6138 13354
rect 6082 13300 6138 13302
rect 2492 12850 2548 12852
rect 2492 12798 2494 12850
rect 2494 12798 2546 12850
rect 2546 12798 2548 12850
rect 2492 12796 2548 12798
rect 10536 12570 10592 12572
rect 10536 12518 10538 12570
rect 10538 12518 10590 12570
rect 10590 12518 10592 12570
rect 10536 12516 10592 12518
rect 10640 12570 10696 12572
rect 10640 12518 10642 12570
rect 10642 12518 10694 12570
rect 10694 12518 10696 12570
rect 10640 12516 10696 12518
rect 10744 12570 10800 12572
rect 10744 12518 10746 12570
rect 10746 12518 10798 12570
rect 10798 12518 10800 12570
rect 10744 12516 10800 12518
rect 5874 11786 5930 11788
rect 5874 11734 5876 11786
rect 5876 11734 5928 11786
rect 5928 11734 5930 11786
rect 5874 11732 5930 11734
rect 5978 11786 6034 11788
rect 5978 11734 5980 11786
rect 5980 11734 6032 11786
rect 6032 11734 6034 11786
rect 5978 11732 6034 11734
rect 6082 11786 6138 11788
rect 6082 11734 6084 11786
rect 6084 11734 6136 11786
rect 6136 11734 6138 11786
rect 6082 11732 6138 11734
rect 10536 11002 10592 11004
rect 10536 10950 10538 11002
rect 10538 10950 10590 11002
rect 10590 10950 10592 11002
rect 10536 10948 10592 10950
rect 10640 11002 10696 11004
rect 10640 10950 10642 11002
rect 10642 10950 10694 11002
rect 10694 10950 10696 11002
rect 10640 10948 10696 10950
rect 10744 11002 10800 11004
rect 10744 10950 10746 11002
rect 10746 10950 10798 11002
rect 10798 10950 10800 11002
rect 10744 10948 10800 10950
rect 5874 10218 5930 10220
rect 5874 10166 5876 10218
rect 5876 10166 5928 10218
rect 5928 10166 5930 10218
rect 5874 10164 5930 10166
rect 5978 10218 6034 10220
rect 5978 10166 5980 10218
rect 5980 10166 6032 10218
rect 6032 10166 6034 10218
rect 5978 10164 6034 10166
rect 6082 10218 6138 10220
rect 6082 10166 6084 10218
rect 6084 10166 6136 10218
rect 6136 10166 6138 10218
rect 6082 10164 6138 10166
rect 10536 9434 10592 9436
rect 10536 9382 10538 9434
rect 10538 9382 10590 9434
rect 10590 9382 10592 9434
rect 10536 9380 10592 9382
rect 10640 9434 10696 9436
rect 10640 9382 10642 9434
rect 10642 9382 10694 9434
rect 10694 9382 10696 9434
rect 10640 9380 10696 9382
rect 10744 9434 10800 9436
rect 10744 9382 10746 9434
rect 10746 9382 10798 9434
rect 10798 9382 10800 9434
rect 10744 9380 10800 9382
rect 5874 8650 5930 8652
rect 5874 8598 5876 8650
rect 5876 8598 5928 8650
rect 5928 8598 5930 8650
rect 5874 8596 5930 8598
rect 5978 8650 6034 8652
rect 5978 8598 5980 8650
rect 5980 8598 6032 8650
rect 6032 8598 6034 8650
rect 5978 8596 6034 8598
rect 6082 8650 6138 8652
rect 6082 8598 6084 8650
rect 6084 8598 6136 8650
rect 6136 8598 6138 8650
rect 6082 8596 6138 8598
rect 10536 7866 10592 7868
rect 10536 7814 10538 7866
rect 10538 7814 10590 7866
rect 10590 7814 10592 7866
rect 10536 7812 10592 7814
rect 10640 7866 10696 7868
rect 10640 7814 10642 7866
rect 10642 7814 10694 7866
rect 10694 7814 10696 7866
rect 10640 7812 10696 7814
rect 10744 7866 10800 7868
rect 10744 7814 10746 7866
rect 10746 7814 10798 7866
rect 10798 7814 10800 7866
rect 10744 7812 10800 7814
rect 5874 7082 5930 7084
rect 5874 7030 5876 7082
rect 5876 7030 5928 7082
rect 5928 7030 5930 7082
rect 5874 7028 5930 7030
rect 5978 7082 6034 7084
rect 5978 7030 5980 7082
rect 5980 7030 6032 7082
rect 6032 7030 6034 7082
rect 5978 7028 6034 7030
rect 6082 7082 6138 7084
rect 6082 7030 6084 7082
rect 6084 7030 6136 7082
rect 6136 7030 6138 7082
rect 6082 7028 6138 7030
rect 10536 6298 10592 6300
rect 10536 6246 10538 6298
rect 10538 6246 10590 6298
rect 10590 6246 10592 6298
rect 10536 6244 10592 6246
rect 10640 6298 10696 6300
rect 10640 6246 10642 6298
rect 10642 6246 10694 6298
rect 10694 6246 10696 6298
rect 10640 6244 10696 6246
rect 10744 6298 10800 6300
rect 10744 6246 10746 6298
rect 10746 6246 10798 6298
rect 10798 6246 10800 6298
rect 10744 6244 10800 6246
rect 5874 5514 5930 5516
rect 5874 5462 5876 5514
rect 5876 5462 5928 5514
rect 5928 5462 5930 5514
rect 5874 5460 5930 5462
rect 5978 5514 6034 5516
rect 5978 5462 5980 5514
rect 5980 5462 6032 5514
rect 6032 5462 6034 5514
rect 5978 5460 6034 5462
rect 6082 5514 6138 5516
rect 6082 5462 6084 5514
rect 6084 5462 6136 5514
rect 6136 5462 6138 5514
rect 6082 5460 6138 5462
rect 10536 4730 10592 4732
rect 10536 4678 10538 4730
rect 10538 4678 10590 4730
rect 10590 4678 10592 4730
rect 10536 4676 10592 4678
rect 10640 4730 10696 4732
rect 10640 4678 10642 4730
rect 10642 4678 10694 4730
rect 10694 4678 10696 4730
rect 10640 4676 10696 4678
rect 10744 4730 10800 4732
rect 10744 4678 10746 4730
rect 10746 4678 10798 4730
rect 10798 4678 10800 4730
rect 10744 4676 10800 4678
rect 5874 3946 5930 3948
rect 5874 3894 5876 3946
rect 5876 3894 5928 3946
rect 5928 3894 5930 3946
rect 5874 3892 5930 3894
rect 5978 3946 6034 3948
rect 5978 3894 5980 3946
rect 5980 3894 6032 3946
rect 6032 3894 6034 3946
rect 5978 3892 6034 3894
rect 6082 3946 6138 3948
rect 6082 3894 6084 3946
rect 6084 3894 6136 3946
rect 6136 3894 6138 3946
rect 6082 3892 6138 3894
rect 10536 3162 10592 3164
rect 10536 3110 10538 3162
rect 10538 3110 10590 3162
rect 10590 3110 10592 3162
rect 10536 3108 10592 3110
rect 10640 3162 10696 3164
rect 10640 3110 10642 3162
rect 10642 3110 10694 3162
rect 10694 3110 10696 3162
rect 10640 3108 10696 3110
rect 10744 3162 10800 3164
rect 10744 3110 10746 3162
rect 10746 3110 10798 3162
rect 10798 3110 10800 3162
rect 10744 3108 10800 3110
rect 15198 13354 15254 13356
rect 15198 13302 15200 13354
rect 15200 13302 15252 13354
rect 15252 13302 15254 13354
rect 15198 13300 15254 13302
rect 15302 13354 15358 13356
rect 15302 13302 15304 13354
rect 15304 13302 15356 13354
rect 15356 13302 15358 13354
rect 15302 13300 15358 13302
rect 15406 13354 15462 13356
rect 15406 13302 15408 13354
rect 15408 13302 15460 13354
rect 15460 13302 15462 13354
rect 15406 13300 15462 13302
rect 15198 11786 15254 11788
rect 15198 11734 15200 11786
rect 15200 11734 15252 11786
rect 15252 11734 15254 11786
rect 15198 11732 15254 11734
rect 15302 11786 15358 11788
rect 15302 11734 15304 11786
rect 15304 11734 15356 11786
rect 15356 11734 15358 11786
rect 15302 11732 15358 11734
rect 15406 11786 15462 11788
rect 15406 11734 15408 11786
rect 15408 11734 15460 11786
rect 15460 11734 15462 11786
rect 15406 11732 15462 11734
rect 15198 10218 15254 10220
rect 15198 10166 15200 10218
rect 15200 10166 15252 10218
rect 15252 10166 15254 10218
rect 15198 10164 15254 10166
rect 15302 10218 15358 10220
rect 15302 10166 15304 10218
rect 15304 10166 15356 10218
rect 15356 10166 15358 10218
rect 15302 10164 15358 10166
rect 15406 10218 15462 10220
rect 15406 10166 15408 10218
rect 15408 10166 15460 10218
rect 15460 10166 15462 10218
rect 15406 10164 15462 10166
rect 15198 8650 15254 8652
rect 15198 8598 15200 8650
rect 15200 8598 15252 8650
rect 15252 8598 15254 8650
rect 15198 8596 15254 8598
rect 15302 8650 15358 8652
rect 15302 8598 15304 8650
rect 15304 8598 15356 8650
rect 15356 8598 15358 8650
rect 15302 8596 15358 8598
rect 15406 8650 15462 8652
rect 15406 8598 15408 8650
rect 15408 8598 15460 8650
rect 15460 8598 15462 8650
rect 15406 8596 15462 8598
rect 15198 7082 15254 7084
rect 15198 7030 15200 7082
rect 15200 7030 15252 7082
rect 15252 7030 15254 7082
rect 15198 7028 15254 7030
rect 15302 7082 15358 7084
rect 15302 7030 15304 7082
rect 15304 7030 15356 7082
rect 15356 7030 15358 7082
rect 15302 7028 15358 7030
rect 15406 7082 15462 7084
rect 15406 7030 15408 7082
rect 15408 7030 15460 7082
rect 15460 7030 15462 7082
rect 15406 7028 15462 7030
rect 15198 5514 15254 5516
rect 15198 5462 15200 5514
rect 15200 5462 15252 5514
rect 15252 5462 15254 5514
rect 15198 5460 15254 5462
rect 15302 5514 15358 5516
rect 15302 5462 15304 5514
rect 15304 5462 15356 5514
rect 15356 5462 15358 5514
rect 15302 5460 15358 5462
rect 15406 5514 15462 5516
rect 15406 5462 15408 5514
rect 15408 5462 15460 5514
rect 15460 5462 15462 5514
rect 15406 5460 15462 5462
rect 15198 3946 15254 3948
rect 15198 3894 15200 3946
rect 15200 3894 15252 3946
rect 15252 3894 15254 3946
rect 15198 3892 15254 3894
rect 15302 3946 15358 3948
rect 15302 3894 15304 3946
rect 15304 3894 15356 3946
rect 15356 3894 15358 3946
rect 15302 3892 15358 3894
rect 15406 3946 15462 3948
rect 15406 3894 15408 3946
rect 15408 3894 15460 3946
rect 15460 3894 15462 3946
rect 15406 3892 15462 3894
rect 16044 18450 16100 18452
rect 16044 18398 16046 18450
rect 16046 18398 16098 18450
rect 16098 18398 16100 18450
rect 16044 18396 16100 18398
rect 15932 18284 15988 18340
rect 16268 17836 16324 17892
rect 16380 18450 16436 18452
rect 16380 18398 16382 18450
rect 16382 18398 16434 18450
rect 16434 18398 16436 18450
rect 16380 18396 16436 18398
rect 16940 19010 16996 19012
rect 16940 18958 16942 19010
rect 16942 18958 16994 19010
rect 16994 18958 16996 19010
rect 16940 18956 16996 18958
rect 17612 19794 17668 19796
rect 17612 19742 17614 19794
rect 17614 19742 17666 19794
rect 17666 19742 17668 19794
rect 17612 19740 17668 19742
rect 18172 19740 18228 19796
rect 17500 18396 17556 18452
rect 17836 18450 17892 18452
rect 17836 18398 17838 18450
rect 17838 18398 17890 18450
rect 17890 18398 17892 18450
rect 17836 18396 17892 18398
rect 16492 18284 16548 18340
rect 17724 18338 17780 18340
rect 17724 18286 17726 18338
rect 17726 18286 17778 18338
rect 17778 18286 17780 18338
rect 17724 18284 17780 18286
rect 16828 18172 16884 18228
rect 16380 17388 16436 17444
rect 18172 17836 18228 17892
rect 18396 19964 18452 20020
rect 19964 20130 20020 20132
rect 19964 20078 19966 20130
rect 19966 20078 20018 20130
rect 20018 20078 20020 20130
rect 19964 20076 20020 20078
rect 19628 20018 19684 20020
rect 19628 19966 19630 20018
rect 19630 19966 19682 20018
rect 19682 19966 19684 20018
rect 19628 19964 19684 19966
rect 19516 19628 19572 19684
rect 18396 18508 18452 18564
rect 18508 18450 18564 18452
rect 18508 18398 18510 18450
rect 18510 18398 18562 18450
rect 18562 18398 18564 18450
rect 18508 18396 18564 18398
rect 19740 19122 19796 19124
rect 19740 19070 19742 19122
rect 19742 19070 19794 19122
rect 19794 19070 19796 19122
rect 19740 19068 19796 19070
rect 19860 18842 19916 18844
rect 19860 18790 19862 18842
rect 19862 18790 19914 18842
rect 19914 18790 19916 18842
rect 19860 18788 19916 18790
rect 19964 18842 20020 18844
rect 19964 18790 19966 18842
rect 19966 18790 20018 18842
rect 20018 18790 20020 18842
rect 19964 18788 20020 18790
rect 20068 18842 20124 18844
rect 20068 18790 20070 18842
rect 20070 18790 20122 18842
rect 20122 18790 20124 18842
rect 20068 18788 20124 18790
rect 19068 18508 19124 18564
rect 19516 18450 19572 18452
rect 19516 18398 19518 18450
rect 19518 18398 19570 18450
rect 19570 18398 19572 18450
rect 19516 18396 19572 18398
rect 18844 18284 18900 18340
rect 19852 18172 19908 18228
rect 20188 18396 20244 18452
rect 16604 17388 16660 17444
rect 15932 16882 15988 16884
rect 15932 16830 15934 16882
rect 15934 16830 15986 16882
rect 15986 16830 15988 16882
rect 15932 16828 15988 16830
rect 16716 16882 16772 16884
rect 16716 16830 16718 16882
rect 16718 16830 16770 16882
rect 16770 16830 16772 16882
rect 16716 16828 16772 16830
rect 16716 15986 16772 15988
rect 16716 15934 16718 15986
rect 16718 15934 16770 15986
rect 16770 15934 16772 15986
rect 16716 15932 16772 15934
rect 16828 14700 16884 14756
rect 17052 14364 17108 14420
rect 16156 14252 16212 14308
rect 16828 13634 16884 13636
rect 16828 13582 16830 13634
rect 16830 13582 16882 13634
rect 16882 13582 16884 13634
rect 16828 13580 16884 13582
rect 17388 13580 17444 13636
rect 18284 17442 18340 17444
rect 18284 17390 18286 17442
rect 18286 17390 18338 17442
rect 18338 17390 18340 17442
rect 18284 17388 18340 17390
rect 18284 17052 18340 17108
rect 17612 16882 17668 16884
rect 17612 16830 17614 16882
rect 17614 16830 17666 16882
rect 17666 16830 17668 16882
rect 17612 16828 17668 16830
rect 18620 16268 18676 16324
rect 18396 16098 18452 16100
rect 18396 16046 18398 16098
rect 18398 16046 18450 16098
rect 18450 16046 18452 16098
rect 18396 16044 18452 16046
rect 18508 15932 18564 15988
rect 18284 14754 18340 14756
rect 18284 14702 18286 14754
rect 18286 14702 18338 14754
rect 18338 14702 18340 14754
rect 18284 14700 18340 14702
rect 18060 14364 18116 14420
rect 17612 13804 17668 13860
rect 17612 13634 17668 13636
rect 17612 13582 17614 13634
rect 17614 13582 17666 13634
rect 17666 13582 17668 13634
rect 17612 13580 17668 13582
rect 17612 13356 17668 13412
rect 16604 12684 16660 12740
rect 17388 12738 17444 12740
rect 17388 12686 17390 12738
rect 17390 12686 17442 12738
rect 17442 12686 17444 12738
rect 17388 12684 17444 12686
rect 18732 15932 18788 15988
rect 18284 13692 18340 13748
rect 18508 13804 18564 13860
rect 18060 13580 18116 13636
rect 17948 11788 18004 11844
rect 18956 15820 19012 15876
rect 19404 16828 19460 16884
rect 19860 17274 19916 17276
rect 19860 17222 19862 17274
rect 19862 17222 19914 17274
rect 19914 17222 19916 17274
rect 19860 17220 19916 17222
rect 19964 17274 20020 17276
rect 19964 17222 19966 17274
rect 19966 17222 20018 17274
rect 20018 17222 20020 17274
rect 19964 17220 20020 17222
rect 20068 17274 20124 17276
rect 20068 17222 20070 17274
rect 20070 17222 20122 17274
rect 20122 17222 20124 17274
rect 20068 17220 20124 17222
rect 20636 20748 20692 20804
rect 20748 20578 20804 20580
rect 20748 20526 20750 20578
rect 20750 20526 20802 20578
rect 20802 20526 20804 20578
rect 20748 20524 20804 20526
rect 20636 19852 20692 19908
rect 21756 23436 21812 23492
rect 21420 22428 21476 22484
rect 21532 22204 21588 22260
rect 21420 21532 21476 21588
rect 21420 19964 21476 20020
rect 23772 24108 23828 24164
rect 24522 35306 24578 35308
rect 24522 35254 24524 35306
rect 24524 35254 24576 35306
rect 24576 35254 24578 35306
rect 24522 35252 24578 35254
rect 24626 35306 24682 35308
rect 24626 35254 24628 35306
rect 24628 35254 24680 35306
rect 24680 35254 24682 35306
rect 24626 35252 24682 35254
rect 24730 35306 24786 35308
rect 24730 35254 24732 35306
rect 24732 35254 24784 35306
rect 24784 35254 24786 35306
rect 24730 35252 24786 35254
rect 24522 33738 24578 33740
rect 24522 33686 24524 33738
rect 24524 33686 24576 33738
rect 24576 33686 24578 33738
rect 24522 33684 24578 33686
rect 24626 33738 24682 33740
rect 24626 33686 24628 33738
rect 24628 33686 24680 33738
rect 24680 33686 24682 33738
rect 24626 33684 24682 33686
rect 24730 33738 24786 33740
rect 24730 33686 24732 33738
rect 24732 33686 24784 33738
rect 24784 33686 24786 33738
rect 24730 33684 24786 33686
rect 24522 32170 24578 32172
rect 24522 32118 24524 32170
rect 24524 32118 24576 32170
rect 24576 32118 24578 32170
rect 24522 32116 24578 32118
rect 24626 32170 24682 32172
rect 24626 32118 24628 32170
rect 24628 32118 24680 32170
rect 24680 32118 24682 32170
rect 24626 32116 24682 32118
rect 24730 32170 24786 32172
rect 24730 32118 24732 32170
rect 24732 32118 24784 32170
rect 24784 32118 24786 32170
rect 24730 32116 24786 32118
rect 24522 30602 24578 30604
rect 24522 30550 24524 30602
rect 24524 30550 24576 30602
rect 24576 30550 24578 30602
rect 24522 30548 24578 30550
rect 24626 30602 24682 30604
rect 24626 30550 24628 30602
rect 24628 30550 24680 30602
rect 24680 30550 24682 30602
rect 24626 30548 24682 30550
rect 24730 30602 24786 30604
rect 24730 30550 24732 30602
rect 24732 30550 24784 30602
rect 24784 30550 24786 30602
rect 24730 30548 24786 30550
rect 24522 29034 24578 29036
rect 24522 28982 24524 29034
rect 24524 28982 24576 29034
rect 24576 28982 24578 29034
rect 24522 28980 24578 28982
rect 24626 29034 24682 29036
rect 24626 28982 24628 29034
rect 24628 28982 24680 29034
rect 24680 28982 24682 29034
rect 24626 28980 24682 28982
rect 24730 29034 24786 29036
rect 24730 28982 24732 29034
rect 24732 28982 24784 29034
rect 24784 28982 24786 29034
rect 24730 28980 24786 28982
rect 24522 27466 24578 27468
rect 24522 27414 24524 27466
rect 24524 27414 24576 27466
rect 24576 27414 24578 27466
rect 24522 27412 24578 27414
rect 24626 27466 24682 27468
rect 24626 27414 24628 27466
rect 24628 27414 24680 27466
rect 24680 27414 24682 27466
rect 24626 27412 24682 27414
rect 24730 27466 24786 27468
rect 24730 27414 24732 27466
rect 24732 27414 24784 27466
rect 24784 27414 24786 27466
rect 24730 27412 24786 27414
rect 36316 36258 36372 36260
rect 36316 36206 36318 36258
rect 36318 36206 36370 36258
rect 36370 36206 36372 36258
rect 36316 36204 36372 36206
rect 29184 36090 29240 36092
rect 29184 36038 29186 36090
rect 29186 36038 29238 36090
rect 29238 36038 29240 36090
rect 29184 36036 29240 36038
rect 29288 36090 29344 36092
rect 29288 36038 29290 36090
rect 29290 36038 29342 36090
rect 29342 36038 29344 36090
rect 29288 36036 29344 36038
rect 29392 36090 29448 36092
rect 29392 36038 29394 36090
rect 29394 36038 29446 36090
rect 29446 36038 29448 36090
rect 29392 36036 29448 36038
rect 33846 35306 33902 35308
rect 33846 35254 33848 35306
rect 33848 35254 33900 35306
rect 33900 35254 33902 35306
rect 33846 35252 33902 35254
rect 33950 35306 34006 35308
rect 33950 35254 33952 35306
rect 33952 35254 34004 35306
rect 34004 35254 34006 35306
rect 33950 35252 34006 35254
rect 34054 35306 34110 35308
rect 34054 35254 34056 35306
rect 34056 35254 34108 35306
rect 34108 35254 34110 35306
rect 34054 35252 34110 35254
rect 29184 34522 29240 34524
rect 29184 34470 29186 34522
rect 29186 34470 29238 34522
rect 29238 34470 29240 34522
rect 29184 34468 29240 34470
rect 29288 34522 29344 34524
rect 29288 34470 29290 34522
rect 29290 34470 29342 34522
rect 29342 34470 29344 34522
rect 29288 34468 29344 34470
rect 29392 34522 29448 34524
rect 29392 34470 29394 34522
rect 29394 34470 29446 34522
rect 29446 34470 29448 34522
rect 29392 34468 29448 34470
rect 33846 33738 33902 33740
rect 33846 33686 33848 33738
rect 33848 33686 33900 33738
rect 33900 33686 33902 33738
rect 33846 33684 33902 33686
rect 33950 33738 34006 33740
rect 33950 33686 33952 33738
rect 33952 33686 34004 33738
rect 34004 33686 34006 33738
rect 33950 33684 34006 33686
rect 34054 33738 34110 33740
rect 34054 33686 34056 33738
rect 34056 33686 34108 33738
rect 34108 33686 34110 33738
rect 34054 33684 34110 33686
rect 28588 33180 28644 33236
rect 25900 26460 25956 26516
rect 27020 30828 27076 30884
rect 24522 25898 24578 25900
rect 24522 25846 24524 25898
rect 24524 25846 24576 25898
rect 24576 25846 24578 25898
rect 24522 25844 24578 25846
rect 24626 25898 24682 25900
rect 24626 25846 24628 25898
rect 24628 25846 24680 25898
rect 24680 25846 24682 25898
rect 24626 25844 24682 25846
rect 24730 25898 24786 25900
rect 24730 25846 24732 25898
rect 24732 25846 24784 25898
rect 24784 25846 24786 25898
rect 24730 25844 24786 25846
rect 26012 25452 26068 25508
rect 26684 25394 26740 25396
rect 26684 25342 26686 25394
rect 26686 25342 26738 25394
rect 26738 25342 26740 25394
rect 26684 25340 26740 25342
rect 26124 24722 26180 24724
rect 26124 24670 26126 24722
rect 26126 24670 26178 24722
rect 26178 24670 26180 24722
rect 26124 24668 26180 24670
rect 24522 24330 24578 24332
rect 24522 24278 24524 24330
rect 24524 24278 24576 24330
rect 24576 24278 24578 24330
rect 24522 24276 24578 24278
rect 24626 24330 24682 24332
rect 24626 24278 24628 24330
rect 24628 24278 24680 24330
rect 24680 24278 24682 24330
rect 24626 24276 24682 24278
rect 24730 24330 24786 24332
rect 24730 24278 24732 24330
rect 24732 24278 24784 24330
rect 24784 24278 24786 24330
rect 24730 24276 24786 24278
rect 24668 24162 24724 24164
rect 24668 24110 24670 24162
rect 24670 24110 24722 24162
rect 24722 24110 24724 24162
rect 24668 24108 24724 24110
rect 24892 23772 24948 23828
rect 25452 24108 25508 24164
rect 25340 23826 25396 23828
rect 25340 23774 25342 23826
rect 25342 23774 25394 23826
rect 25394 23774 25396 23826
rect 25340 23772 25396 23774
rect 25228 23436 25284 23492
rect 23884 23378 23940 23380
rect 23884 23326 23886 23378
rect 23886 23326 23938 23378
rect 23938 23326 23940 23378
rect 23884 23324 23940 23326
rect 22092 23266 22148 23268
rect 22092 23214 22094 23266
rect 22094 23214 22146 23266
rect 22146 23214 22148 23266
rect 22092 23212 22148 23214
rect 21980 23154 22036 23156
rect 21980 23102 21982 23154
rect 21982 23102 22034 23154
rect 22034 23102 22036 23154
rect 21980 23100 22036 23102
rect 23212 22540 23268 22596
rect 21084 19740 21140 19796
rect 22428 22204 22484 22260
rect 24522 22762 24578 22764
rect 24522 22710 24524 22762
rect 24524 22710 24576 22762
rect 24576 22710 24578 22762
rect 24522 22708 24578 22710
rect 24626 22762 24682 22764
rect 24626 22710 24628 22762
rect 24628 22710 24680 22762
rect 24680 22710 24682 22762
rect 24626 22708 24682 22710
rect 24730 22762 24786 22764
rect 24730 22710 24732 22762
rect 24732 22710 24784 22762
rect 24784 22710 24786 22762
rect 24730 22708 24786 22710
rect 25788 23938 25844 23940
rect 25788 23886 25790 23938
rect 25790 23886 25842 23938
rect 25842 23886 25844 23938
rect 25788 23884 25844 23886
rect 26236 23884 26292 23940
rect 26012 23436 26068 23492
rect 23548 22204 23604 22260
rect 23100 21810 23156 21812
rect 23100 21758 23102 21810
rect 23102 21758 23154 21810
rect 23154 21758 23156 21810
rect 23100 21756 23156 21758
rect 21644 20636 21700 20692
rect 24444 21698 24500 21700
rect 24444 21646 24446 21698
rect 24446 21646 24498 21698
rect 24498 21646 24500 21698
rect 24444 21644 24500 21646
rect 23660 21532 23716 21588
rect 23548 20860 23604 20916
rect 22540 20690 22596 20692
rect 22540 20638 22542 20690
rect 22542 20638 22594 20690
rect 22594 20638 22596 20690
rect 22540 20636 22596 20638
rect 21756 20524 21812 20580
rect 24332 21586 24388 21588
rect 24332 21534 24334 21586
rect 24334 21534 24386 21586
rect 24386 21534 24388 21586
rect 24332 21532 24388 21534
rect 25228 21644 25284 21700
rect 24668 21308 24724 21364
rect 24522 21194 24578 21196
rect 24522 21142 24524 21194
rect 24524 21142 24576 21194
rect 24576 21142 24578 21194
rect 24522 21140 24578 21142
rect 24626 21194 24682 21196
rect 24626 21142 24628 21194
rect 24628 21142 24680 21194
rect 24680 21142 24682 21194
rect 24626 21140 24682 21142
rect 24730 21194 24786 21196
rect 24730 21142 24732 21194
rect 24732 21142 24784 21194
rect 24784 21142 24786 21194
rect 24730 21140 24786 21142
rect 25564 21532 25620 21588
rect 25452 21308 25508 21364
rect 24444 20972 24500 21028
rect 25340 20690 25396 20692
rect 25340 20638 25342 20690
rect 25342 20638 25394 20690
rect 25394 20638 25396 20690
rect 25340 20636 25396 20638
rect 22092 20076 22148 20132
rect 23996 20130 24052 20132
rect 23996 20078 23998 20130
rect 23998 20078 24050 20130
rect 24050 20078 24052 20130
rect 23996 20076 24052 20078
rect 22652 20018 22708 20020
rect 22652 19966 22654 20018
rect 22654 19966 22706 20018
rect 22706 19966 22708 20018
rect 22652 19964 22708 19966
rect 21532 19292 21588 19348
rect 22428 19628 22484 19684
rect 21868 19180 21924 19236
rect 21084 19068 21140 19124
rect 20300 18172 20356 18228
rect 21084 18450 21140 18452
rect 21084 18398 21086 18450
rect 21086 18398 21138 18450
rect 21138 18398 21140 18450
rect 21084 18396 21140 18398
rect 21756 18396 21812 18452
rect 20860 18284 20916 18340
rect 21980 18338 22036 18340
rect 21980 18286 21982 18338
rect 21982 18286 22034 18338
rect 22034 18286 22036 18338
rect 21980 18284 22036 18286
rect 20748 17442 20804 17444
rect 20748 17390 20750 17442
rect 20750 17390 20802 17442
rect 20802 17390 20804 17442
rect 20748 17388 20804 17390
rect 20300 16940 20356 16996
rect 21084 16994 21140 16996
rect 21084 16942 21086 16994
rect 21086 16942 21138 16994
rect 21138 16942 21140 16994
rect 21084 16940 21140 16942
rect 22092 17500 22148 17556
rect 21532 16940 21588 16996
rect 20412 16882 20468 16884
rect 20412 16830 20414 16882
rect 20414 16830 20466 16882
rect 20466 16830 20468 16882
rect 20412 16828 20468 16830
rect 19516 16322 19572 16324
rect 19516 16270 19518 16322
rect 19518 16270 19570 16322
rect 19570 16270 19572 16322
rect 19516 16268 19572 16270
rect 20524 16268 20580 16324
rect 19068 15036 19124 15092
rect 19068 14476 19124 14532
rect 19404 14700 19460 14756
rect 19180 14418 19236 14420
rect 19180 14366 19182 14418
rect 19182 14366 19234 14418
rect 19234 14366 19236 14418
rect 19180 14364 19236 14366
rect 19068 14306 19124 14308
rect 19068 14254 19070 14306
rect 19070 14254 19122 14306
rect 19122 14254 19124 14306
rect 19068 14252 19124 14254
rect 18844 11788 18900 11844
rect 20188 16044 20244 16100
rect 20076 15932 20132 15988
rect 19860 15706 19916 15708
rect 19860 15654 19862 15706
rect 19862 15654 19914 15706
rect 19914 15654 19916 15706
rect 19860 15652 19916 15654
rect 19964 15706 20020 15708
rect 19964 15654 19966 15706
rect 19966 15654 20018 15706
rect 20018 15654 20020 15706
rect 19964 15652 20020 15654
rect 20068 15706 20124 15708
rect 20068 15654 20070 15706
rect 20070 15654 20122 15706
rect 20122 15654 20124 15706
rect 20068 15652 20124 15654
rect 20412 15874 20468 15876
rect 20412 15822 20414 15874
rect 20414 15822 20466 15874
rect 20466 15822 20468 15874
rect 20412 15820 20468 15822
rect 20188 15426 20244 15428
rect 20188 15374 20190 15426
rect 20190 15374 20242 15426
rect 20242 15374 20244 15426
rect 20188 15372 20244 15374
rect 19740 15036 19796 15092
rect 21308 16210 21364 16212
rect 21308 16158 21310 16210
rect 21310 16158 21362 16210
rect 21362 16158 21364 16210
rect 21308 16156 21364 16158
rect 21532 16322 21588 16324
rect 21532 16270 21534 16322
rect 21534 16270 21586 16322
rect 21586 16270 21588 16322
rect 21532 16268 21588 16270
rect 21868 15874 21924 15876
rect 21868 15822 21870 15874
rect 21870 15822 21922 15874
rect 21922 15822 21924 15874
rect 21868 15820 21924 15822
rect 21868 15372 21924 15428
rect 19860 14138 19916 14140
rect 19860 14086 19862 14138
rect 19862 14086 19914 14138
rect 19914 14086 19916 14138
rect 19860 14084 19916 14086
rect 19964 14138 20020 14140
rect 19964 14086 19966 14138
rect 19966 14086 20018 14138
rect 20018 14086 20020 14138
rect 19964 14084 20020 14086
rect 20068 14138 20124 14140
rect 20068 14086 20070 14138
rect 20070 14086 20122 14138
rect 20122 14086 20124 14138
rect 20068 14084 20124 14086
rect 19964 13858 20020 13860
rect 19964 13806 19966 13858
rect 19966 13806 20018 13858
rect 20018 13806 20020 13858
rect 19964 13804 20020 13806
rect 20636 12908 20692 12964
rect 22540 19346 22596 19348
rect 22540 19294 22542 19346
rect 22542 19294 22594 19346
rect 22594 19294 22596 19346
rect 22540 19292 22596 19294
rect 22988 19292 23044 19348
rect 22764 18338 22820 18340
rect 22764 18286 22766 18338
rect 22766 18286 22818 18338
rect 22818 18286 22820 18338
rect 22764 18284 22820 18286
rect 24522 19626 24578 19628
rect 24522 19574 24524 19626
rect 24524 19574 24576 19626
rect 24576 19574 24578 19626
rect 24522 19572 24578 19574
rect 24626 19626 24682 19628
rect 24626 19574 24628 19626
rect 24628 19574 24680 19626
rect 24680 19574 24682 19626
rect 24626 19572 24682 19574
rect 24730 19626 24786 19628
rect 24730 19574 24732 19626
rect 24732 19574 24784 19626
rect 24784 19574 24786 19626
rect 24730 19572 24786 19574
rect 23436 19292 23492 19348
rect 23100 19122 23156 19124
rect 23100 19070 23102 19122
rect 23102 19070 23154 19122
rect 23154 19070 23156 19122
rect 23100 19068 23156 19070
rect 23996 19122 24052 19124
rect 23996 19070 23998 19122
rect 23998 19070 24050 19122
rect 24050 19070 24052 19122
rect 23996 19068 24052 19070
rect 26124 23100 26180 23156
rect 27804 27132 27860 27188
rect 27132 24946 27188 24948
rect 27132 24894 27134 24946
rect 27134 24894 27186 24946
rect 27186 24894 27188 24946
rect 27132 24892 27188 24894
rect 27244 24668 27300 24724
rect 27580 24444 27636 24500
rect 27132 23660 27188 23716
rect 27356 23772 27412 23828
rect 27356 23212 27412 23268
rect 26348 21644 26404 21700
rect 25788 20636 25844 20692
rect 29184 32954 29240 32956
rect 29184 32902 29186 32954
rect 29186 32902 29238 32954
rect 29238 32902 29240 32954
rect 29184 32900 29240 32902
rect 29288 32954 29344 32956
rect 29288 32902 29290 32954
rect 29290 32902 29342 32954
rect 29342 32902 29344 32954
rect 29288 32900 29344 32902
rect 29392 32954 29448 32956
rect 29392 32902 29394 32954
rect 29394 32902 29446 32954
rect 29446 32902 29448 32954
rect 29392 32900 29448 32902
rect 33846 32170 33902 32172
rect 33846 32118 33848 32170
rect 33848 32118 33900 32170
rect 33900 32118 33902 32170
rect 33846 32116 33902 32118
rect 33950 32170 34006 32172
rect 33950 32118 33952 32170
rect 33952 32118 34004 32170
rect 34004 32118 34006 32170
rect 33950 32116 34006 32118
rect 34054 32170 34110 32172
rect 34054 32118 34056 32170
rect 34056 32118 34108 32170
rect 34108 32118 34110 32170
rect 34054 32116 34110 32118
rect 36876 36370 36932 36372
rect 36876 36318 36878 36370
rect 36878 36318 36930 36370
rect 36930 36318 36932 36370
rect 36876 36316 36932 36318
rect 37100 35698 37156 35700
rect 37100 35646 37102 35698
rect 37102 35646 37154 35698
rect 37154 35646 37156 35698
rect 37100 35644 37156 35646
rect 37212 35196 37268 35252
rect 38220 36258 38276 36260
rect 38220 36206 38222 36258
rect 38222 36206 38274 36258
rect 38274 36206 38276 36258
rect 38220 36204 38276 36206
rect 37996 35698 38052 35700
rect 37996 35646 37998 35698
rect 37998 35646 38050 35698
rect 38050 35646 38052 35698
rect 37996 35644 38052 35646
rect 29184 31386 29240 31388
rect 29184 31334 29186 31386
rect 29186 31334 29238 31386
rect 29238 31334 29240 31386
rect 29184 31332 29240 31334
rect 29288 31386 29344 31388
rect 29288 31334 29290 31386
rect 29290 31334 29342 31386
rect 29342 31334 29344 31386
rect 29288 31332 29344 31334
rect 29392 31386 29448 31388
rect 29392 31334 29394 31386
rect 29394 31334 29446 31386
rect 29446 31334 29448 31386
rect 29392 31332 29448 31334
rect 33846 30602 33902 30604
rect 33846 30550 33848 30602
rect 33848 30550 33900 30602
rect 33900 30550 33902 30602
rect 33846 30548 33902 30550
rect 33950 30602 34006 30604
rect 33950 30550 33952 30602
rect 33952 30550 34004 30602
rect 34004 30550 34006 30602
rect 33950 30548 34006 30550
rect 34054 30602 34110 30604
rect 34054 30550 34056 30602
rect 34056 30550 34108 30602
rect 34108 30550 34110 30602
rect 34054 30548 34110 30550
rect 29184 29818 29240 29820
rect 29184 29766 29186 29818
rect 29186 29766 29238 29818
rect 29238 29766 29240 29818
rect 29184 29764 29240 29766
rect 29288 29818 29344 29820
rect 29288 29766 29290 29818
rect 29290 29766 29342 29818
rect 29342 29766 29344 29818
rect 29288 29764 29344 29766
rect 29392 29818 29448 29820
rect 29392 29766 29394 29818
rect 29394 29766 29446 29818
rect 29446 29766 29448 29818
rect 29392 29764 29448 29766
rect 33846 29034 33902 29036
rect 33846 28982 33848 29034
rect 33848 28982 33900 29034
rect 33900 28982 33902 29034
rect 33846 28980 33902 28982
rect 33950 29034 34006 29036
rect 33950 28982 33952 29034
rect 33952 28982 34004 29034
rect 34004 28982 34006 29034
rect 33950 28980 34006 28982
rect 34054 29034 34110 29036
rect 34054 28982 34056 29034
rect 34056 28982 34108 29034
rect 34108 28982 34110 29034
rect 34054 28980 34110 28982
rect 29184 28250 29240 28252
rect 29184 28198 29186 28250
rect 29186 28198 29238 28250
rect 29238 28198 29240 28250
rect 29184 28196 29240 28198
rect 29288 28250 29344 28252
rect 29288 28198 29290 28250
rect 29290 28198 29342 28250
rect 29342 28198 29344 28250
rect 29288 28196 29344 28198
rect 29392 28250 29448 28252
rect 29392 28198 29394 28250
rect 29394 28198 29446 28250
rect 29446 28198 29448 28250
rect 29392 28196 29448 28198
rect 30380 27804 30436 27860
rect 29184 26682 29240 26684
rect 29184 26630 29186 26682
rect 29186 26630 29238 26682
rect 29238 26630 29240 26682
rect 29184 26628 29240 26630
rect 29288 26682 29344 26684
rect 29288 26630 29290 26682
rect 29290 26630 29342 26682
rect 29342 26630 29344 26682
rect 29288 26628 29344 26630
rect 29392 26682 29448 26684
rect 29392 26630 29394 26682
rect 29394 26630 29446 26682
rect 29446 26630 29448 26682
rect 29392 26628 29448 26630
rect 28700 24892 28756 24948
rect 29484 25394 29540 25396
rect 29484 25342 29486 25394
rect 29486 25342 29538 25394
rect 29538 25342 29540 25394
rect 29484 25340 29540 25342
rect 29184 25114 29240 25116
rect 29184 25062 29186 25114
rect 29186 25062 29238 25114
rect 29238 25062 29240 25114
rect 29184 25060 29240 25062
rect 29288 25114 29344 25116
rect 29288 25062 29290 25114
rect 29290 25062 29342 25114
rect 29342 25062 29344 25114
rect 29288 25060 29344 25062
rect 29392 25114 29448 25116
rect 29392 25062 29394 25114
rect 29394 25062 29446 25114
rect 29446 25062 29448 25114
rect 29392 25060 29448 25062
rect 27804 24722 27860 24724
rect 27804 24670 27806 24722
rect 27806 24670 27858 24722
rect 27858 24670 27860 24722
rect 27804 24668 27860 24670
rect 28588 24668 28644 24724
rect 28028 24498 28084 24500
rect 28028 24446 28030 24498
rect 28030 24446 28082 24498
rect 28082 24446 28084 24498
rect 28028 24444 28084 24446
rect 28364 24444 28420 24500
rect 30156 24946 30212 24948
rect 30156 24894 30158 24946
rect 30158 24894 30210 24946
rect 30210 24894 30212 24946
rect 30156 24892 30212 24894
rect 29708 24722 29764 24724
rect 29708 24670 29710 24722
rect 29710 24670 29762 24722
rect 29762 24670 29764 24722
rect 29708 24668 29764 24670
rect 28924 24498 28980 24500
rect 28924 24446 28926 24498
rect 28926 24446 28978 24498
rect 28978 24446 28980 24498
rect 28924 24444 28980 24446
rect 28812 24108 28868 24164
rect 28588 23826 28644 23828
rect 28588 23774 28590 23826
rect 28590 23774 28642 23826
rect 28642 23774 28644 23826
rect 28588 23772 28644 23774
rect 28476 23212 28532 23268
rect 26796 21698 26852 21700
rect 26796 21646 26798 21698
rect 26798 21646 26850 21698
rect 26850 21646 26852 21698
rect 26796 21644 26852 21646
rect 26572 21532 26628 21588
rect 27468 21698 27524 21700
rect 27468 21646 27470 21698
rect 27470 21646 27522 21698
rect 27522 21646 27524 21698
rect 27468 21644 27524 21646
rect 27244 21308 27300 21364
rect 27356 21586 27412 21588
rect 27356 21534 27358 21586
rect 27358 21534 27410 21586
rect 27410 21534 27412 21586
rect 27356 21532 27412 21534
rect 26684 20578 26740 20580
rect 26684 20526 26686 20578
rect 26686 20526 26738 20578
rect 26738 20526 26740 20578
rect 26684 20524 26740 20526
rect 26012 19852 26068 19908
rect 26012 19292 26068 19348
rect 24332 19122 24388 19124
rect 24332 19070 24334 19122
rect 24334 19070 24386 19122
rect 24386 19070 24388 19122
rect 24332 19068 24388 19070
rect 25340 19122 25396 19124
rect 25340 19070 25342 19122
rect 25342 19070 25394 19122
rect 25394 19070 25396 19122
rect 25340 19068 25396 19070
rect 22988 18172 23044 18228
rect 22652 17554 22708 17556
rect 22652 17502 22654 17554
rect 22654 17502 22706 17554
rect 22706 17502 22708 17554
rect 22652 17500 22708 17502
rect 23100 17554 23156 17556
rect 23100 17502 23102 17554
rect 23102 17502 23154 17554
rect 23154 17502 23156 17554
rect 23100 17500 23156 17502
rect 24444 18172 24500 18228
rect 24522 18058 24578 18060
rect 24522 18006 24524 18058
rect 24524 18006 24576 18058
rect 24576 18006 24578 18058
rect 24522 18004 24578 18006
rect 24626 18058 24682 18060
rect 24626 18006 24628 18058
rect 24628 18006 24680 18058
rect 24680 18006 24682 18058
rect 24626 18004 24682 18006
rect 24730 18058 24786 18060
rect 24730 18006 24732 18058
rect 24732 18006 24784 18058
rect 24784 18006 24786 18058
rect 24730 18004 24786 18006
rect 22876 16882 22932 16884
rect 22876 16830 22878 16882
rect 22878 16830 22930 16882
rect 22930 16830 22932 16882
rect 22876 16828 22932 16830
rect 23324 16882 23380 16884
rect 23324 16830 23326 16882
rect 23326 16830 23378 16882
rect 23378 16830 23380 16882
rect 23324 16828 23380 16830
rect 23100 16156 23156 16212
rect 22764 16044 22820 16100
rect 23660 17500 23716 17556
rect 23548 16044 23604 16100
rect 23212 15148 23268 15204
rect 21868 13634 21924 13636
rect 21868 13582 21870 13634
rect 21870 13582 21922 13634
rect 21922 13582 21924 13634
rect 21868 13580 21924 13582
rect 22316 13634 22372 13636
rect 22316 13582 22318 13634
rect 22318 13582 22370 13634
rect 22370 13582 22372 13634
rect 22316 13580 22372 13582
rect 22764 13634 22820 13636
rect 22764 13582 22766 13634
rect 22766 13582 22818 13634
rect 22818 13582 22820 13634
rect 22764 13580 22820 13582
rect 20188 12684 20244 12740
rect 21420 12738 21476 12740
rect 21420 12686 21422 12738
rect 21422 12686 21474 12738
rect 21474 12686 21476 12738
rect 21420 12684 21476 12686
rect 19860 12570 19916 12572
rect 19860 12518 19862 12570
rect 19862 12518 19914 12570
rect 19914 12518 19916 12570
rect 19860 12516 19916 12518
rect 19964 12570 20020 12572
rect 19964 12518 19966 12570
rect 19966 12518 20018 12570
rect 20018 12518 20020 12570
rect 19964 12516 20020 12518
rect 20068 12570 20124 12572
rect 20068 12518 20070 12570
rect 20070 12518 20122 12570
rect 20122 12518 20124 12570
rect 20068 12516 20124 12518
rect 19860 11002 19916 11004
rect 19860 10950 19862 11002
rect 19862 10950 19914 11002
rect 19914 10950 19916 11002
rect 19860 10948 19916 10950
rect 19964 11002 20020 11004
rect 19964 10950 19966 11002
rect 19966 10950 20018 11002
rect 20018 10950 20020 11002
rect 19964 10948 20020 10950
rect 20068 11002 20124 11004
rect 20068 10950 20070 11002
rect 20070 10950 20122 11002
rect 20122 10950 20124 11002
rect 20068 10948 20124 10950
rect 19860 9434 19916 9436
rect 19860 9382 19862 9434
rect 19862 9382 19914 9434
rect 19914 9382 19916 9434
rect 19860 9380 19916 9382
rect 19964 9434 20020 9436
rect 19964 9382 19966 9434
rect 19966 9382 20018 9434
rect 20018 9382 20020 9434
rect 19964 9380 20020 9382
rect 20068 9434 20124 9436
rect 20068 9382 20070 9434
rect 20070 9382 20122 9434
rect 20122 9382 20124 9434
rect 20068 9380 20124 9382
rect 19860 7866 19916 7868
rect 19860 7814 19862 7866
rect 19862 7814 19914 7866
rect 19914 7814 19916 7866
rect 19860 7812 19916 7814
rect 19964 7866 20020 7868
rect 19964 7814 19966 7866
rect 19966 7814 20018 7866
rect 20018 7814 20020 7866
rect 19964 7812 20020 7814
rect 20068 7866 20124 7868
rect 20068 7814 20070 7866
rect 20070 7814 20122 7866
rect 20122 7814 20124 7866
rect 20068 7812 20124 7814
rect 19860 6298 19916 6300
rect 19860 6246 19862 6298
rect 19862 6246 19914 6298
rect 19914 6246 19916 6298
rect 19860 6244 19916 6246
rect 19964 6298 20020 6300
rect 19964 6246 19966 6298
rect 19966 6246 20018 6298
rect 20018 6246 20020 6298
rect 19964 6244 20020 6246
rect 20068 6298 20124 6300
rect 20068 6246 20070 6298
rect 20070 6246 20122 6298
rect 20122 6246 20124 6298
rect 20068 6244 20124 6246
rect 19860 4730 19916 4732
rect 19860 4678 19862 4730
rect 19862 4678 19914 4730
rect 19914 4678 19916 4730
rect 19860 4676 19916 4678
rect 19964 4730 20020 4732
rect 19964 4678 19966 4730
rect 19966 4678 20018 4730
rect 20018 4678 20020 4730
rect 19964 4676 20020 4678
rect 20068 4730 20124 4732
rect 20068 4678 20070 4730
rect 20070 4678 20122 4730
rect 20122 4678 20124 4730
rect 20068 4676 20124 4678
rect 21980 12962 22036 12964
rect 21980 12910 21982 12962
rect 21982 12910 22034 12962
rect 22034 12910 22036 12962
rect 21980 12908 22036 12910
rect 22764 11788 22820 11844
rect 23548 13804 23604 13860
rect 23324 13692 23380 13748
rect 24332 17554 24388 17556
rect 24332 17502 24334 17554
rect 24334 17502 24386 17554
rect 24386 17502 24388 17554
rect 24332 17500 24388 17502
rect 24780 17500 24836 17556
rect 24220 16604 24276 16660
rect 24522 16490 24578 16492
rect 24522 16438 24524 16490
rect 24524 16438 24576 16490
rect 24576 16438 24578 16490
rect 24522 16436 24578 16438
rect 24626 16490 24682 16492
rect 24626 16438 24628 16490
rect 24628 16438 24680 16490
rect 24680 16438 24682 16490
rect 24626 16436 24682 16438
rect 24730 16490 24786 16492
rect 24730 16438 24732 16490
rect 24732 16438 24784 16490
rect 24784 16438 24786 16490
rect 24730 16436 24786 16438
rect 24220 16210 24276 16212
rect 24220 16158 24222 16210
rect 24222 16158 24274 16210
rect 24274 16158 24276 16210
rect 24220 16156 24276 16158
rect 24444 16098 24500 16100
rect 24444 16046 24446 16098
rect 24446 16046 24498 16098
rect 24498 16046 24500 16098
rect 24444 16044 24500 16046
rect 24780 15986 24836 15988
rect 24780 15934 24782 15986
rect 24782 15934 24834 15986
rect 24834 15934 24836 15986
rect 24780 15932 24836 15934
rect 24332 15820 24388 15876
rect 23772 15314 23828 15316
rect 23772 15262 23774 15314
rect 23774 15262 23826 15314
rect 23826 15262 23828 15314
rect 23772 15260 23828 15262
rect 23884 13746 23940 13748
rect 23884 13694 23886 13746
rect 23886 13694 23938 13746
rect 23938 13694 23940 13746
rect 23884 13692 23940 13694
rect 23660 12684 23716 12740
rect 24220 15148 24276 15204
rect 24220 13746 24276 13748
rect 24220 13694 24222 13746
rect 24222 13694 24274 13746
rect 24274 13694 24276 13746
rect 24220 13692 24276 13694
rect 24108 11788 24164 11844
rect 23548 4956 23604 5012
rect 24108 3500 24164 3556
rect 19860 3162 19916 3164
rect 19860 3110 19862 3162
rect 19862 3110 19914 3162
rect 19914 3110 19916 3162
rect 19860 3108 19916 3110
rect 19964 3162 20020 3164
rect 19964 3110 19966 3162
rect 19966 3110 20018 3162
rect 20018 3110 20020 3162
rect 19964 3108 20020 3110
rect 20068 3162 20124 3164
rect 20068 3110 20070 3162
rect 20070 3110 20122 3162
rect 20122 3110 20124 3162
rect 20068 3108 20124 3110
rect 24220 3388 24276 3444
rect 24522 14922 24578 14924
rect 24522 14870 24524 14922
rect 24524 14870 24576 14922
rect 24576 14870 24578 14922
rect 24522 14868 24578 14870
rect 24626 14922 24682 14924
rect 24626 14870 24628 14922
rect 24628 14870 24680 14922
rect 24680 14870 24682 14922
rect 24626 14868 24682 14870
rect 24730 14922 24786 14924
rect 24730 14870 24732 14922
rect 24732 14870 24784 14922
rect 24784 14870 24786 14922
rect 24730 14868 24786 14870
rect 24668 13634 24724 13636
rect 24668 13582 24670 13634
rect 24670 13582 24722 13634
rect 24722 13582 24724 13634
rect 24668 13580 24724 13582
rect 24522 13354 24578 13356
rect 24522 13302 24524 13354
rect 24524 13302 24576 13354
rect 24576 13302 24578 13354
rect 24522 13300 24578 13302
rect 24626 13354 24682 13356
rect 24626 13302 24628 13354
rect 24628 13302 24680 13354
rect 24680 13302 24682 13354
rect 24626 13300 24682 13302
rect 24730 13354 24786 13356
rect 24730 13302 24732 13354
rect 24732 13302 24784 13354
rect 24784 13302 24786 13354
rect 24730 13300 24786 13302
rect 24444 12738 24500 12740
rect 24444 12686 24446 12738
rect 24446 12686 24498 12738
rect 24498 12686 24500 12738
rect 24444 12684 24500 12686
rect 24522 11786 24578 11788
rect 24522 11734 24524 11786
rect 24524 11734 24576 11786
rect 24576 11734 24578 11786
rect 24522 11732 24578 11734
rect 24626 11786 24682 11788
rect 24626 11734 24628 11786
rect 24628 11734 24680 11786
rect 24680 11734 24682 11786
rect 24626 11732 24682 11734
rect 24730 11786 24786 11788
rect 24730 11734 24732 11786
rect 24732 11734 24784 11786
rect 24784 11734 24786 11786
rect 24730 11732 24786 11734
rect 24522 10218 24578 10220
rect 24522 10166 24524 10218
rect 24524 10166 24576 10218
rect 24576 10166 24578 10218
rect 24522 10164 24578 10166
rect 24626 10218 24682 10220
rect 24626 10166 24628 10218
rect 24628 10166 24680 10218
rect 24680 10166 24682 10218
rect 24626 10164 24682 10166
rect 24730 10218 24786 10220
rect 24730 10166 24732 10218
rect 24732 10166 24784 10218
rect 24784 10166 24786 10218
rect 24730 10164 24786 10166
rect 24522 8650 24578 8652
rect 24522 8598 24524 8650
rect 24524 8598 24576 8650
rect 24576 8598 24578 8650
rect 24522 8596 24578 8598
rect 24626 8650 24682 8652
rect 24626 8598 24628 8650
rect 24628 8598 24680 8650
rect 24680 8598 24682 8650
rect 24626 8596 24682 8598
rect 24730 8650 24786 8652
rect 24730 8598 24732 8650
rect 24732 8598 24784 8650
rect 24784 8598 24786 8650
rect 24730 8596 24786 8598
rect 25676 19010 25732 19012
rect 25676 18958 25678 19010
rect 25678 18958 25730 19010
rect 25730 18958 25732 19010
rect 25676 18956 25732 18958
rect 26348 19010 26404 19012
rect 26348 18958 26350 19010
rect 26350 18958 26402 19010
rect 26402 18958 26404 19010
rect 26348 18956 26404 18958
rect 28140 20690 28196 20692
rect 28140 20638 28142 20690
rect 28142 20638 28194 20690
rect 28194 20638 28196 20690
rect 28140 20636 28196 20638
rect 26908 19852 26964 19908
rect 26684 19740 26740 19796
rect 28252 19964 28308 20020
rect 29148 24108 29204 24164
rect 29184 23546 29240 23548
rect 29184 23494 29186 23546
rect 29186 23494 29238 23546
rect 29238 23494 29240 23546
rect 29184 23492 29240 23494
rect 29288 23546 29344 23548
rect 29288 23494 29290 23546
rect 29290 23494 29342 23546
rect 29342 23494 29344 23546
rect 29288 23492 29344 23494
rect 29392 23546 29448 23548
rect 29392 23494 29394 23546
rect 29394 23494 29446 23546
rect 29446 23494 29448 23546
rect 29392 23492 29448 23494
rect 33846 27466 33902 27468
rect 33846 27414 33848 27466
rect 33848 27414 33900 27466
rect 33900 27414 33902 27466
rect 33846 27412 33902 27414
rect 33950 27466 34006 27468
rect 33950 27414 33952 27466
rect 33952 27414 34004 27466
rect 34004 27414 34006 27466
rect 33950 27412 34006 27414
rect 34054 27466 34110 27468
rect 34054 27414 34056 27466
rect 34056 27414 34108 27466
rect 34108 27414 34110 27466
rect 34054 27412 34110 27414
rect 33846 25898 33902 25900
rect 33846 25846 33848 25898
rect 33848 25846 33900 25898
rect 33900 25846 33902 25898
rect 33846 25844 33902 25846
rect 33950 25898 34006 25900
rect 33950 25846 33952 25898
rect 33952 25846 34004 25898
rect 34004 25846 34006 25898
rect 33950 25844 34006 25846
rect 34054 25898 34110 25900
rect 34054 25846 34056 25898
rect 34056 25846 34108 25898
rect 34108 25846 34110 25898
rect 34054 25844 34110 25846
rect 33846 24330 33902 24332
rect 33846 24278 33848 24330
rect 33848 24278 33900 24330
rect 33900 24278 33902 24330
rect 33846 24276 33902 24278
rect 33950 24330 34006 24332
rect 33950 24278 33952 24330
rect 33952 24278 34004 24330
rect 34004 24278 34006 24330
rect 33950 24276 34006 24278
rect 34054 24330 34110 24332
rect 34054 24278 34056 24330
rect 34056 24278 34108 24330
rect 34108 24278 34110 24330
rect 34054 24276 34110 24278
rect 28924 23266 28980 23268
rect 28924 23214 28926 23266
rect 28926 23214 28978 23266
rect 28978 23214 28980 23266
rect 28924 23212 28980 23214
rect 29260 22258 29316 22260
rect 29260 22206 29262 22258
rect 29262 22206 29314 22258
rect 29314 22206 29316 22258
rect 29260 22204 29316 22206
rect 31276 23436 31332 23492
rect 30492 22316 30548 22372
rect 29184 21978 29240 21980
rect 29184 21926 29186 21978
rect 29186 21926 29238 21978
rect 29238 21926 29240 21978
rect 29184 21924 29240 21926
rect 29288 21978 29344 21980
rect 29288 21926 29290 21978
rect 29290 21926 29342 21978
rect 29342 21926 29344 21978
rect 29288 21924 29344 21926
rect 29392 21978 29448 21980
rect 29392 21926 29394 21978
rect 29394 21926 29446 21978
rect 29446 21926 29448 21978
rect 29392 21924 29448 21926
rect 29596 21868 29652 21924
rect 29148 21698 29204 21700
rect 29148 21646 29150 21698
rect 29150 21646 29202 21698
rect 29202 21646 29204 21698
rect 29148 21644 29204 21646
rect 29820 22204 29876 22260
rect 30268 21980 30324 22036
rect 29708 21644 29764 21700
rect 29036 21532 29092 21588
rect 28700 21420 28756 21476
rect 29260 21084 29316 21140
rect 29260 20802 29316 20804
rect 29260 20750 29262 20802
rect 29262 20750 29314 20802
rect 29314 20750 29316 20802
rect 29260 20748 29316 20750
rect 30380 21420 30436 21476
rect 29184 20410 29240 20412
rect 29184 20358 29186 20410
rect 29186 20358 29238 20410
rect 29238 20358 29240 20410
rect 29184 20356 29240 20358
rect 29288 20410 29344 20412
rect 29288 20358 29290 20410
rect 29290 20358 29342 20410
rect 29342 20358 29344 20410
rect 29288 20356 29344 20358
rect 29392 20410 29448 20412
rect 29392 20358 29394 20410
rect 29394 20358 29446 20410
rect 29446 20358 29448 20410
rect 29392 20356 29448 20358
rect 28924 20130 28980 20132
rect 28924 20078 28926 20130
rect 28926 20078 28978 20130
rect 28978 20078 28980 20130
rect 28924 20076 28980 20078
rect 30604 22258 30660 22260
rect 30604 22206 30606 22258
rect 30606 22206 30658 22258
rect 30658 22206 30660 22258
rect 30604 22204 30660 22206
rect 33846 22762 33902 22764
rect 33846 22710 33848 22762
rect 33848 22710 33900 22762
rect 33900 22710 33902 22762
rect 33846 22708 33902 22710
rect 33950 22762 34006 22764
rect 33950 22710 33952 22762
rect 33952 22710 34004 22762
rect 34004 22710 34006 22762
rect 33950 22708 34006 22710
rect 34054 22762 34110 22764
rect 34054 22710 34056 22762
rect 34056 22710 34108 22762
rect 34108 22710 34110 22762
rect 34054 22708 34110 22710
rect 36540 31554 36596 31556
rect 36540 31502 36542 31554
rect 36542 31502 36594 31554
rect 36594 31502 36596 31554
rect 36540 31500 36596 31502
rect 38508 36090 38564 36092
rect 38508 36038 38510 36090
rect 38510 36038 38562 36090
rect 38562 36038 38564 36090
rect 38508 36036 38564 36038
rect 38612 36090 38668 36092
rect 38612 36038 38614 36090
rect 38614 36038 38666 36090
rect 38666 36038 38668 36090
rect 38612 36036 38668 36038
rect 38716 36090 38772 36092
rect 38716 36038 38718 36090
rect 38718 36038 38770 36090
rect 38770 36038 38772 36090
rect 38716 36036 38772 36038
rect 38332 35644 38388 35700
rect 39116 35196 39172 35252
rect 38220 34972 38276 35028
rect 38508 34522 38564 34524
rect 38508 34470 38510 34522
rect 38510 34470 38562 34522
rect 38562 34470 38564 34522
rect 38508 34468 38564 34470
rect 38612 34522 38668 34524
rect 38612 34470 38614 34522
rect 38614 34470 38666 34522
rect 38666 34470 38668 34522
rect 38612 34468 38668 34470
rect 38716 34522 38772 34524
rect 38716 34470 38718 34522
rect 38718 34470 38770 34522
rect 38770 34470 38772 34522
rect 38716 34468 38772 34470
rect 38444 34300 38500 34356
rect 38220 33628 38276 33684
rect 37884 33234 37940 33236
rect 37884 33182 37886 33234
rect 37886 33182 37938 33234
rect 37938 33182 37940 33234
rect 37884 33180 37940 33182
rect 38220 33122 38276 33124
rect 38220 33070 38222 33122
rect 38222 33070 38274 33122
rect 38274 33070 38276 33122
rect 38220 33068 38276 33070
rect 38508 32954 38564 32956
rect 38508 32902 38510 32954
rect 38510 32902 38562 32954
rect 38562 32902 38564 32954
rect 38508 32900 38564 32902
rect 38612 32954 38668 32956
rect 38612 32902 38614 32954
rect 38614 32902 38666 32954
rect 38666 32902 38668 32954
rect 38612 32900 38668 32902
rect 38716 32954 38772 32956
rect 38716 32902 38718 32954
rect 38718 32902 38770 32954
rect 38770 32902 38772 32954
rect 38716 32900 38772 32902
rect 37212 32284 37268 32340
rect 38220 32284 38276 32340
rect 37212 31500 37268 31556
rect 37212 27132 37268 27188
rect 37100 25340 37156 25396
rect 37212 26572 37268 26628
rect 36988 24892 37044 24948
rect 37548 31666 37604 31668
rect 37548 31614 37550 31666
rect 37550 31614 37602 31666
rect 37602 31614 37604 31666
rect 37548 31612 37604 31614
rect 37548 30882 37604 30884
rect 37548 30830 37550 30882
rect 37550 30830 37602 30882
rect 37602 30830 37604 30882
rect 37548 30828 37604 30830
rect 38508 31386 38564 31388
rect 38508 31334 38510 31386
rect 38510 31334 38562 31386
rect 38562 31334 38564 31386
rect 38508 31332 38564 31334
rect 38612 31386 38668 31388
rect 38612 31334 38614 31386
rect 38614 31334 38666 31386
rect 38666 31334 38668 31386
rect 38612 31332 38668 31334
rect 38716 31386 38772 31388
rect 38716 31334 38718 31386
rect 38718 31334 38770 31386
rect 38770 31334 38772 31386
rect 38716 31332 38772 31334
rect 38444 30940 38500 30996
rect 38220 30268 38276 30324
rect 38220 29708 38276 29764
rect 38508 29818 38564 29820
rect 38508 29766 38510 29818
rect 38510 29766 38562 29818
rect 38562 29766 38564 29818
rect 38508 29764 38564 29766
rect 38612 29818 38668 29820
rect 38612 29766 38614 29818
rect 38614 29766 38666 29818
rect 38666 29766 38668 29818
rect 38612 29764 38668 29766
rect 38716 29818 38772 29820
rect 38716 29766 38718 29818
rect 38718 29766 38770 29818
rect 38770 29766 38772 29818
rect 38716 29764 38772 29766
rect 37324 25452 37380 25508
rect 37324 24108 37380 24164
rect 37548 27020 37604 27076
rect 37884 27858 37940 27860
rect 37884 27806 37886 27858
rect 37886 27806 37938 27858
rect 37938 27806 37940 27858
rect 37884 27804 37940 27806
rect 38220 28924 38276 28980
rect 38220 28418 38276 28420
rect 38220 28366 38222 28418
rect 38222 28366 38274 28418
rect 38274 28366 38276 28418
rect 38220 28364 38276 28366
rect 38508 28250 38564 28252
rect 38508 28198 38510 28250
rect 38510 28198 38562 28250
rect 38562 28198 38564 28250
rect 38508 28196 38564 28198
rect 38612 28250 38668 28252
rect 38612 28198 38614 28250
rect 38614 28198 38666 28250
rect 38666 28198 38668 28250
rect 38612 28196 38668 28198
rect 38716 28250 38772 28252
rect 38716 28198 38718 28250
rect 38718 28198 38770 28250
rect 38770 28198 38772 28250
rect 38716 28196 38772 28198
rect 38220 27580 38276 27636
rect 37660 26572 37716 26628
rect 37660 26178 37716 26180
rect 37660 26126 37662 26178
rect 37662 26126 37714 26178
rect 37714 26126 37716 26178
rect 37660 26124 37716 26126
rect 37548 23436 37604 23492
rect 37436 23324 37492 23380
rect 36428 22204 36484 22260
rect 30940 21868 30996 21924
rect 37100 21756 37156 21812
rect 33846 21194 33902 21196
rect 33846 21142 33848 21194
rect 33848 21142 33900 21194
rect 33900 21142 33902 21194
rect 33846 21140 33902 21142
rect 33950 21194 34006 21196
rect 33950 21142 33952 21194
rect 33952 21142 34004 21194
rect 34004 21142 34006 21194
rect 33950 21140 34006 21142
rect 34054 21194 34110 21196
rect 34054 21142 34056 21194
rect 34056 21142 34108 21194
rect 34108 21142 34110 21194
rect 34054 21140 34110 21142
rect 37548 21532 37604 21588
rect 38508 26682 38564 26684
rect 38508 26630 38510 26682
rect 38510 26630 38562 26682
rect 38562 26630 38564 26682
rect 38508 26628 38564 26630
rect 38612 26682 38668 26684
rect 38612 26630 38614 26682
rect 38614 26630 38666 26682
rect 38666 26630 38668 26682
rect 38612 26628 38668 26630
rect 38716 26682 38772 26684
rect 38716 26630 38718 26682
rect 38718 26630 38770 26682
rect 38770 26630 38772 26682
rect 38716 26628 38772 26630
rect 38108 26348 38164 26404
rect 38220 26124 38276 26180
rect 38220 25564 38276 25620
rect 38220 25004 38276 25060
rect 38508 25114 38564 25116
rect 38508 25062 38510 25114
rect 38510 25062 38562 25114
rect 38562 25062 38564 25114
rect 38508 25060 38564 25062
rect 38612 25114 38668 25116
rect 38612 25062 38614 25114
rect 38614 25062 38666 25114
rect 38666 25062 38668 25114
rect 38612 25060 38668 25062
rect 38716 25114 38772 25116
rect 38716 25062 38718 25114
rect 38718 25062 38770 25114
rect 38770 25062 38772 25114
rect 38716 25060 38772 25062
rect 37884 23154 37940 23156
rect 37884 23102 37886 23154
rect 37886 23102 37938 23154
rect 37938 23102 37940 23154
rect 37884 23100 37940 23102
rect 37772 22540 37828 22596
rect 37996 22316 38052 22372
rect 37884 21980 37940 22036
rect 37660 20972 37716 21028
rect 37212 20860 37268 20916
rect 37884 20524 37940 20580
rect 37884 20130 37940 20132
rect 37884 20078 37886 20130
rect 37886 20078 37938 20130
rect 37938 20078 37940 20130
rect 37884 20076 37940 20078
rect 28364 19404 28420 19460
rect 27244 19122 27300 19124
rect 27244 19070 27246 19122
rect 27246 19070 27298 19122
rect 27298 19070 27300 19122
rect 27244 19068 27300 19070
rect 26572 18562 26628 18564
rect 26572 18510 26574 18562
rect 26574 18510 26626 18562
rect 26626 18510 26628 18562
rect 26572 18508 26628 18510
rect 27356 18508 27412 18564
rect 26460 18450 26516 18452
rect 26460 18398 26462 18450
rect 26462 18398 26514 18450
rect 26514 18398 26516 18450
rect 26460 18396 26516 18398
rect 25452 17052 25508 17108
rect 26572 17052 26628 17108
rect 26460 16882 26516 16884
rect 26460 16830 26462 16882
rect 26462 16830 26514 16882
rect 26514 16830 26516 16882
rect 26460 16828 26516 16830
rect 25564 16716 25620 16772
rect 26236 16770 26292 16772
rect 26236 16718 26238 16770
rect 26238 16718 26290 16770
rect 26290 16718 26292 16770
rect 26236 16716 26292 16718
rect 25116 15986 25172 15988
rect 25116 15934 25118 15986
rect 25118 15934 25170 15986
rect 25170 15934 25172 15986
rect 25116 15932 25172 15934
rect 25900 16210 25956 16212
rect 25900 16158 25902 16210
rect 25902 16158 25954 16210
rect 25954 16158 25956 16210
rect 25900 16156 25956 16158
rect 24892 7980 24948 8036
rect 24522 7082 24578 7084
rect 24522 7030 24524 7082
rect 24524 7030 24576 7082
rect 24576 7030 24578 7082
rect 24522 7028 24578 7030
rect 24626 7082 24682 7084
rect 24626 7030 24628 7082
rect 24628 7030 24680 7082
rect 24680 7030 24682 7082
rect 24626 7028 24682 7030
rect 24730 7082 24786 7084
rect 24730 7030 24732 7082
rect 24732 7030 24784 7082
rect 24784 7030 24786 7082
rect 24730 7028 24786 7030
rect 24522 5514 24578 5516
rect 24522 5462 24524 5514
rect 24524 5462 24576 5514
rect 24576 5462 24578 5514
rect 24522 5460 24578 5462
rect 24626 5514 24682 5516
rect 24626 5462 24628 5514
rect 24628 5462 24680 5514
rect 24680 5462 24682 5514
rect 24626 5460 24682 5462
rect 24730 5514 24786 5516
rect 24730 5462 24732 5514
rect 24732 5462 24784 5514
rect 24784 5462 24786 5514
rect 24730 5460 24786 5462
rect 25228 15314 25284 15316
rect 25228 15262 25230 15314
rect 25230 15262 25282 15314
rect 25282 15262 25284 15314
rect 25228 15260 25284 15262
rect 25228 13746 25284 13748
rect 25228 13694 25230 13746
rect 25230 13694 25282 13746
rect 25282 13694 25284 13746
rect 25228 13692 25284 13694
rect 25564 14476 25620 14532
rect 25452 11228 25508 11284
rect 25004 4172 25060 4228
rect 24522 3946 24578 3948
rect 24522 3894 24524 3946
rect 24524 3894 24576 3946
rect 24576 3894 24578 3946
rect 24522 3892 24578 3894
rect 24626 3946 24682 3948
rect 24626 3894 24628 3946
rect 24628 3894 24680 3946
rect 24680 3894 24682 3946
rect 24626 3892 24682 3894
rect 24730 3946 24786 3948
rect 24730 3894 24732 3946
rect 24732 3894 24784 3946
rect 24784 3894 24786 3946
rect 24730 3892 24786 3894
rect 24892 3612 24948 3668
rect 24780 3554 24836 3556
rect 24780 3502 24782 3554
rect 24782 3502 24834 3554
rect 24834 3502 24836 3554
rect 24780 3500 24836 3502
rect 25900 13580 25956 13636
rect 25676 3612 25732 3668
rect 25228 3442 25284 3444
rect 25228 3390 25230 3442
rect 25230 3390 25282 3442
rect 25282 3390 25284 3442
rect 25228 3388 25284 3390
rect 26572 12684 26628 12740
rect 26124 3612 26180 3668
rect 26124 3388 26180 3444
rect 26908 16828 26964 16884
rect 28364 19068 28420 19124
rect 27468 18396 27524 18452
rect 27916 18620 27972 18676
rect 28364 18508 28420 18564
rect 38220 24220 38276 24276
rect 38220 23714 38276 23716
rect 38220 23662 38222 23714
rect 38222 23662 38274 23714
rect 38274 23662 38276 23714
rect 38220 23660 38276 23662
rect 38508 23546 38564 23548
rect 38508 23494 38510 23546
rect 38510 23494 38562 23546
rect 38562 23494 38564 23546
rect 38508 23492 38564 23494
rect 38612 23546 38668 23548
rect 38612 23494 38614 23546
rect 38614 23494 38666 23546
rect 38666 23494 38668 23546
rect 38612 23492 38668 23494
rect 38716 23546 38772 23548
rect 38716 23494 38718 23546
rect 38718 23494 38770 23546
rect 38770 23494 38772 23546
rect 38716 23492 38772 23494
rect 39116 25340 39172 25396
rect 39116 24668 39172 24724
rect 39004 23772 39060 23828
rect 38892 23212 38948 23268
rect 38220 22876 38276 22932
rect 38220 22258 38276 22260
rect 38220 22206 38222 22258
rect 38222 22206 38274 22258
rect 38274 22206 38276 22258
rect 38220 22204 38276 22206
rect 38508 21978 38564 21980
rect 38508 21926 38510 21978
rect 38510 21926 38562 21978
rect 38562 21926 38564 21978
rect 38508 21924 38564 21926
rect 38612 21978 38668 21980
rect 38612 21926 38614 21978
rect 38614 21926 38666 21978
rect 38666 21926 38668 21978
rect 38612 21924 38668 21926
rect 38716 21978 38772 21980
rect 38716 21926 38718 21978
rect 38718 21926 38770 21978
rect 38770 21926 38772 21978
rect 38716 21924 38772 21926
rect 38220 20860 38276 20916
rect 38108 20636 38164 20692
rect 38508 20410 38564 20412
rect 38508 20358 38510 20410
rect 38510 20358 38562 20410
rect 38562 20358 38564 20410
rect 38508 20356 38564 20358
rect 38612 20410 38668 20412
rect 38612 20358 38614 20410
rect 38614 20358 38666 20410
rect 38666 20358 38668 20410
rect 38612 20356 38668 20358
rect 38716 20410 38772 20412
rect 38716 20358 38718 20410
rect 38718 20358 38770 20410
rect 38770 20358 38772 20410
rect 38716 20356 38772 20358
rect 38444 20188 38500 20244
rect 37996 19964 38052 20020
rect 29036 19068 29092 19124
rect 28700 18956 28756 19012
rect 28588 18620 28644 18676
rect 28924 18732 28980 18788
rect 29596 19122 29652 19124
rect 29596 19070 29598 19122
rect 29598 19070 29650 19122
rect 29650 19070 29652 19122
rect 29596 19068 29652 19070
rect 29484 18956 29540 19012
rect 29184 18842 29240 18844
rect 29184 18790 29186 18842
rect 29186 18790 29238 18842
rect 29238 18790 29240 18842
rect 29184 18788 29240 18790
rect 29288 18842 29344 18844
rect 29288 18790 29290 18842
rect 29290 18790 29342 18842
rect 29342 18790 29344 18842
rect 29288 18788 29344 18790
rect 29392 18842 29448 18844
rect 29392 18790 29394 18842
rect 29394 18790 29446 18842
rect 29446 18790 29448 18842
rect 29392 18788 29448 18790
rect 30156 19068 30212 19124
rect 29596 18508 29652 18564
rect 30044 18956 30100 19012
rect 30268 18508 30324 18564
rect 28364 18338 28420 18340
rect 28364 18286 28366 18338
rect 28366 18286 28418 18338
rect 28418 18286 28420 18338
rect 28364 18284 28420 18286
rect 27132 17388 27188 17444
rect 28476 17388 28532 17444
rect 27020 16716 27076 16772
rect 27132 15314 27188 15316
rect 27132 15262 27134 15314
rect 27134 15262 27186 15314
rect 27186 15262 27188 15314
rect 27132 15260 27188 15262
rect 27468 16770 27524 16772
rect 27468 16718 27470 16770
rect 27470 16718 27522 16770
rect 27522 16718 27524 16770
rect 27468 16716 27524 16718
rect 27356 15202 27412 15204
rect 27356 15150 27358 15202
rect 27358 15150 27410 15202
rect 27410 15150 27412 15202
rect 27356 15148 27412 15150
rect 27468 14418 27524 14420
rect 27468 14366 27470 14418
rect 27470 14366 27522 14418
rect 27522 14366 27524 14418
rect 27468 14364 27524 14366
rect 28028 15314 28084 15316
rect 28028 15262 28030 15314
rect 28030 15262 28082 15314
rect 28082 15262 28084 15314
rect 28028 15260 28084 15262
rect 28476 15260 28532 15316
rect 28140 13692 28196 13748
rect 27916 10556 27972 10612
rect 29932 18284 29988 18340
rect 29260 17442 29316 17444
rect 29260 17390 29262 17442
rect 29262 17390 29314 17442
rect 29314 17390 29316 17442
rect 29260 17388 29316 17390
rect 29184 17274 29240 17276
rect 29184 17222 29186 17274
rect 29186 17222 29238 17274
rect 29238 17222 29240 17274
rect 29184 17220 29240 17222
rect 29288 17274 29344 17276
rect 29288 17222 29290 17274
rect 29290 17222 29342 17274
rect 29342 17222 29344 17274
rect 29288 17220 29344 17222
rect 29392 17274 29448 17276
rect 29392 17222 29394 17274
rect 29394 17222 29446 17274
rect 29446 17222 29448 17274
rect 29392 17220 29448 17222
rect 29820 16882 29876 16884
rect 29820 16830 29822 16882
rect 29822 16830 29874 16882
rect 29874 16830 29876 16882
rect 29820 16828 29876 16830
rect 29148 16604 29204 16660
rect 29184 15706 29240 15708
rect 29184 15654 29186 15706
rect 29186 15654 29238 15706
rect 29238 15654 29240 15706
rect 29184 15652 29240 15654
rect 29288 15706 29344 15708
rect 29288 15654 29290 15706
rect 29290 15654 29342 15706
rect 29342 15654 29344 15706
rect 29288 15652 29344 15654
rect 29392 15706 29448 15708
rect 29392 15654 29394 15706
rect 29394 15654 29446 15706
rect 29446 15654 29448 15706
rect 29392 15652 29448 15654
rect 29820 15314 29876 15316
rect 29820 15262 29822 15314
rect 29822 15262 29874 15314
rect 29874 15262 29876 15314
rect 29820 15260 29876 15262
rect 28924 15202 28980 15204
rect 28924 15150 28926 15202
rect 28926 15150 28978 15202
rect 28978 15150 28980 15202
rect 28924 15148 28980 15150
rect 29820 14306 29876 14308
rect 29820 14254 29822 14306
rect 29822 14254 29874 14306
rect 29874 14254 29876 14306
rect 29820 14252 29876 14254
rect 29184 14138 29240 14140
rect 29184 14086 29186 14138
rect 29186 14086 29238 14138
rect 29238 14086 29240 14138
rect 29184 14084 29240 14086
rect 29288 14138 29344 14140
rect 29288 14086 29290 14138
rect 29290 14086 29342 14138
rect 29342 14086 29344 14138
rect 29288 14084 29344 14086
rect 29392 14138 29448 14140
rect 29392 14086 29394 14138
rect 29394 14086 29446 14138
rect 29446 14086 29448 14138
rect 29392 14084 29448 14086
rect 29184 12570 29240 12572
rect 29184 12518 29186 12570
rect 29186 12518 29238 12570
rect 29238 12518 29240 12570
rect 29184 12516 29240 12518
rect 29288 12570 29344 12572
rect 29288 12518 29290 12570
rect 29290 12518 29342 12570
rect 29342 12518 29344 12570
rect 29288 12516 29344 12518
rect 29392 12570 29448 12572
rect 29392 12518 29394 12570
rect 29394 12518 29446 12570
rect 29446 12518 29448 12570
rect 29392 12516 29448 12518
rect 29184 11002 29240 11004
rect 29184 10950 29186 11002
rect 29186 10950 29238 11002
rect 29238 10950 29240 11002
rect 29184 10948 29240 10950
rect 29288 11002 29344 11004
rect 29288 10950 29290 11002
rect 29290 10950 29342 11002
rect 29342 10950 29344 11002
rect 29288 10948 29344 10950
rect 29392 11002 29448 11004
rect 29392 10950 29394 11002
rect 29394 10950 29446 11002
rect 29446 10950 29448 11002
rect 29392 10948 29448 10950
rect 29184 9434 29240 9436
rect 29184 9382 29186 9434
rect 29186 9382 29238 9434
rect 29238 9382 29240 9434
rect 29184 9380 29240 9382
rect 29288 9434 29344 9436
rect 29288 9382 29290 9434
rect 29290 9382 29342 9434
rect 29342 9382 29344 9434
rect 29288 9380 29344 9382
rect 29392 9434 29448 9436
rect 29392 9382 29394 9434
rect 29394 9382 29446 9434
rect 29446 9382 29448 9434
rect 29392 9380 29448 9382
rect 29184 7866 29240 7868
rect 29184 7814 29186 7866
rect 29186 7814 29238 7866
rect 29238 7814 29240 7866
rect 29184 7812 29240 7814
rect 29288 7866 29344 7868
rect 29288 7814 29290 7866
rect 29290 7814 29342 7866
rect 29342 7814 29344 7866
rect 29288 7812 29344 7814
rect 29392 7866 29448 7868
rect 29392 7814 29394 7866
rect 29394 7814 29446 7866
rect 29446 7814 29448 7866
rect 29392 7812 29448 7814
rect 28588 7308 28644 7364
rect 26684 6524 26740 6580
rect 29184 6298 29240 6300
rect 29184 6246 29186 6298
rect 29186 6246 29238 6298
rect 29238 6246 29240 6298
rect 29184 6244 29240 6246
rect 29288 6298 29344 6300
rect 29288 6246 29290 6298
rect 29290 6246 29342 6298
rect 29342 6246 29344 6298
rect 29288 6244 29344 6246
rect 29392 6298 29448 6300
rect 29392 6246 29394 6298
rect 29394 6246 29446 6298
rect 29446 6246 29448 6298
rect 29392 6244 29448 6246
rect 30044 16658 30100 16660
rect 30044 16606 30046 16658
rect 30046 16606 30098 16658
rect 30098 16606 30100 16658
rect 30044 16604 30100 16606
rect 30716 19122 30772 19124
rect 30716 19070 30718 19122
rect 30718 19070 30770 19122
rect 30770 19070 30772 19122
rect 30716 19068 30772 19070
rect 30604 18956 30660 19012
rect 33846 19626 33902 19628
rect 33846 19574 33848 19626
rect 33848 19574 33900 19626
rect 33900 19574 33902 19626
rect 33846 19572 33902 19574
rect 33950 19626 34006 19628
rect 33950 19574 33952 19626
rect 33952 19574 34004 19626
rect 34004 19574 34006 19626
rect 33950 19572 34006 19574
rect 34054 19626 34110 19628
rect 34054 19574 34056 19626
rect 34056 19574 34108 19626
rect 34108 19574 34110 19626
rect 34054 19572 34110 19574
rect 38220 19516 38276 19572
rect 37884 19234 37940 19236
rect 37884 19182 37886 19234
rect 37886 19182 37938 19234
rect 37938 19182 37940 19234
rect 37884 19180 37940 19182
rect 30940 18620 30996 18676
rect 30380 17388 30436 17444
rect 30492 18284 30548 18340
rect 30492 16828 30548 16884
rect 30716 17388 30772 17444
rect 31724 18338 31780 18340
rect 31724 18286 31726 18338
rect 31726 18286 31778 18338
rect 31778 18286 31780 18338
rect 31724 18284 31780 18286
rect 30716 16882 30772 16884
rect 30716 16830 30718 16882
rect 30718 16830 30770 16882
rect 30770 16830 30772 16882
rect 30716 16828 30772 16830
rect 30940 16658 30996 16660
rect 30940 16606 30942 16658
rect 30942 16606 30994 16658
rect 30994 16606 30996 16658
rect 30940 16604 30996 16606
rect 30156 15260 30212 15316
rect 31052 12796 31108 12852
rect 30828 10892 30884 10948
rect 31500 15314 31556 15316
rect 31500 15262 31502 15314
rect 31502 15262 31554 15314
rect 31554 15262 31556 15314
rect 31500 15260 31556 15262
rect 29932 5740 29988 5796
rect 31276 5068 31332 5124
rect 27468 4956 27524 5012
rect 29184 4730 29240 4732
rect 29184 4678 29186 4730
rect 29186 4678 29238 4730
rect 29238 4678 29240 4730
rect 29184 4676 29240 4678
rect 29288 4730 29344 4732
rect 29288 4678 29290 4730
rect 29290 4678 29342 4730
rect 29342 4678 29344 4730
rect 29288 4676 29344 4678
rect 29392 4730 29448 4732
rect 29392 4678 29394 4730
rect 29394 4678 29446 4730
rect 29446 4678 29448 4730
rect 29392 4676 29448 4678
rect 27244 3442 27300 3444
rect 27244 3390 27246 3442
rect 27246 3390 27298 3442
rect 27298 3390 27300 3442
rect 27244 3388 27300 3390
rect 38220 19010 38276 19012
rect 38220 18958 38222 19010
rect 38222 18958 38274 19010
rect 38274 18958 38276 19010
rect 38220 18956 38276 18958
rect 38508 18842 38564 18844
rect 38508 18790 38510 18842
rect 38510 18790 38562 18842
rect 38562 18790 38564 18842
rect 38508 18788 38564 18790
rect 38612 18842 38668 18844
rect 38612 18790 38614 18842
rect 38614 18790 38666 18842
rect 38666 18790 38668 18842
rect 38612 18788 38668 18790
rect 38716 18842 38772 18844
rect 38716 18790 38718 18842
rect 38718 18790 38770 18842
rect 38770 18790 38772 18842
rect 38716 18788 38772 18790
rect 37884 18450 37940 18452
rect 37884 18398 37886 18450
rect 37886 18398 37938 18450
rect 37938 18398 37940 18450
rect 37884 18396 37940 18398
rect 37436 18284 37492 18340
rect 33846 18058 33902 18060
rect 33846 18006 33848 18058
rect 33848 18006 33900 18058
rect 33900 18006 33902 18058
rect 33846 18004 33902 18006
rect 33950 18058 34006 18060
rect 33950 18006 33952 18058
rect 33952 18006 34004 18058
rect 34004 18006 34006 18058
rect 33950 18004 34006 18006
rect 34054 18058 34110 18060
rect 34054 18006 34056 18058
rect 34056 18006 34108 18058
rect 34108 18006 34110 18058
rect 34054 18004 34110 18006
rect 37212 17554 37268 17556
rect 37212 17502 37214 17554
rect 37214 17502 37266 17554
rect 37266 17502 37268 17554
rect 37212 17500 37268 17502
rect 32396 16882 32452 16884
rect 32396 16830 32398 16882
rect 32398 16830 32450 16882
rect 32450 16830 32452 16882
rect 32396 16828 32452 16830
rect 37100 16828 37156 16884
rect 33846 16490 33902 16492
rect 33846 16438 33848 16490
rect 33848 16438 33900 16490
rect 33900 16438 33902 16490
rect 33846 16436 33902 16438
rect 33950 16490 34006 16492
rect 33950 16438 33952 16490
rect 33952 16438 34004 16490
rect 34004 16438 34006 16490
rect 33950 16436 34006 16438
rect 34054 16490 34110 16492
rect 34054 16438 34056 16490
rect 34056 16438 34108 16490
rect 34108 16438 34110 16490
rect 34054 16436 34110 16438
rect 31948 16044 32004 16100
rect 33846 14922 33902 14924
rect 33846 14870 33848 14922
rect 33848 14870 33900 14922
rect 33900 14870 33902 14922
rect 33846 14868 33902 14870
rect 33950 14922 34006 14924
rect 33950 14870 33952 14922
rect 33952 14870 34004 14922
rect 34004 14870 34006 14922
rect 33950 14868 34006 14870
rect 34054 14922 34110 14924
rect 34054 14870 34056 14922
rect 34056 14870 34108 14922
rect 34108 14870 34110 14922
rect 34054 14868 34110 14870
rect 33846 13354 33902 13356
rect 33846 13302 33848 13354
rect 33848 13302 33900 13354
rect 33900 13302 33902 13354
rect 33846 13300 33902 13302
rect 33950 13354 34006 13356
rect 33950 13302 33952 13354
rect 33952 13302 34004 13354
rect 34004 13302 34006 13354
rect 33950 13300 34006 13302
rect 34054 13354 34110 13356
rect 34054 13302 34056 13354
rect 34056 13302 34108 13354
rect 34108 13302 34110 13354
rect 34054 13300 34110 13302
rect 33846 11786 33902 11788
rect 33846 11734 33848 11786
rect 33848 11734 33900 11786
rect 33900 11734 33902 11786
rect 33846 11732 33902 11734
rect 33950 11786 34006 11788
rect 33950 11734 33952 11786
rect 33952 11734 34004 11786
rect 34004 11734 34006 11786
rect 33950 11732 34006 11734
rect 34054 11786 34110 11788
rect 34054 11734 34056 11786
rect 34056 11734 34108 11786
rect 34108 11734 34110 11786
rect 34054 11732 34110 11734
rect 33846 10218 33902 10220
rect 33846 10166 33848 10218
rect 33848 10166 33900 10218
rect 33900 10166 33902 10218
rect 33846 10164 33902 10166
rect 33950 10218 34006 10220
rect 33950 10166 33952 10218
rect 33952 10166 34004 10218
rect 34004 10166 34006 10218
rect 33950 10164 34006 10166
rect 34054 10218 34110 10220
rect 34054 10166 34056 10218
rect 34056 10166 34108 10218
rect 34108 10166 34110 10218
rect 34054 10164 34110 10166
rect 33846 8650 33902 8652
rect 33846 8598 33848 8650
rect 33848 8598 33900 8650
rect 33900 8598 33902 8650
rect 33846 8596 33902 8598
rect 33950 8650 34006 8652
rect 33950 8598 33952 8650
rect 33952 8598 34004 8650
rect 34004 8598 34006 8650
rect 33950 8596 34006 8598
rect 34054 8650 34110 8652
rect 34054 8598 34056 8650
rect 34056 8598 34108 8650
rect 34108 8598 34110 8650
rect 34054 8596 34110 8598
rect 36428 8034 36484 8036
rect 36428 7982 36430 8034
rect 36430 7982 36482 8034
rect 36482 7982 36484 8034
rect 36428 7980 36484 7982
rect 33846 7082 33902 7084
rect 33846 7030 33848 7082
rect 33848 7030 33900 7082
rect 33900 7030 33902 7082
rect 33846 7028 33902 7030
rect 33950 7082 34006 7084
rect 33950 7030 33952 7082
rect 33952 7030 34004 7082
rect 34004 7030 34006 7082
rect 33950 7028 34006 7030
rect 34054 7082 34110 7084
rect 34054 7030 34056 7082
rect 34056 7030 34108 7082
rect 34108 7030 34110 7082
rect 34054 7028 34110 7030
rect 33846 5514 33902 5516
rect 33846 5462 33848 5514
rect 33848 5462 33900 5514
rect 33900 5462 33902 5514
rect 33846 5460 33902 5462
rect 33950 5514 34006 5516
rect 33950 5462 33952 5514
rect 33952 5462 34004 5514
rect 34004 5462 34006 5514
rect 33950 5460 34006 5462
rect 34054 5514 34110 5516
rect 34054 5462 34056 5514
rect 34056 5462 34108 5514
rect 34108 5462 34110 5514
rect 34054 5460 34110 5462
rect 33846 3946 33902 3948
rect 33846 3894 33848 3946
rect 33848 3894 33900 3946
rect 33900 3894 33902 3946
rect 33846 3892 33902 3894
rect 33950 3946 34006 3948
rect 33950 3894 33952 3946
rect 33952 3894 34004 3946
rect 34004 3894 34006 3946
rect 33950 3892 34006 3894
rect 34054 3946 34110 3948
rect 34054 3894 34056 3946
rect 34056 3894 34108 3946
rect 34108 3894 34110 3946
rect 34054 3892 34110 3894
rect 31836 3388 31892 3444
rect 36428 3442 36484 3444
rect 36428 3390 36430 3442
rect 36430 3390 36482 3442
rect 36482 3390 36484 3442
rect 36428 3388 36484 3390
rect 37212 14476 37268 14532
rect 37324 10892 37380 10948
rect 38220 18172 38276 18228
rect 37884 17666 37940 17668
rect 37884 17614 37886 17666
rect 37886 17614 37938 17666
rect 37938 17614 37940 17666
rect 37884 17612 37940 17614
rect 38220 17554 38276 17556
rect 38220 17502 38222 17554
rect 38222 17502 38274 17554
rect 38274 17502 38276 17554
rect 38220 17500 38276 17502
rect 38508 17274 38564 17276
rect 38508 17222 38510 17274
rect 38510 17222 38562 17274
rect 38562 17222 38564 17274
rect 38508 17220 38564 17222
rect 38612 17274 38668 17276
rect 38612 17222 38614 17274
rect 38614 17222 38666 17274
rect 38666 17222 38668 17274
rect 38612 17220 38668 17222
rect 38716 17274 38772 17276
rect 38716 17222 38718 17274
rect 38718 17222 38770 17274
rect 38770 17222 38772 17274
rect 38716 17220 38772 17222
rect 37884 16994 37940 16996
rect 37884 16942 37886 16994
rect 37886 16942 37938 16994
rect 37938 16942 37940 16994
rect 37884 16940 37940 16942
rect 37548 16828 37604 16884
rect 38220 16156 38276 16212
rect 37884 16098 37940 16100
rect 37884 16046 37886 16098
rect 37886 16046 37938 16098
rect 37938 16046 37940 16098
rect 37884 16044 37940 16046
rect 38508 15706 38564 15708
rect 38508 15654 38510 15706
rect 38510 15654 38562 15706
rect 38562 15654 38564 15706
rect 38508 15652 38564 15654
rect 38612 15706 38668 15708
rect 38612 15654 38614 15706
rect 38614 15654 38666 15706
rect 38666 15654 38668 15706
rect 38612 15652 38668 15654
rect 38716 15706 38772 15708
rect 38716 15654 38718 15706
rect 38718 15654 38770 15706
rect 38770 15654 38772 15706
rect 38716 15652 38772 15654
rect 38444 15484 38500 15540
rect 37772 15148 37828 15204
rect 37884 14588 37940 14644
rect 37996 15260 38052 15316
rect 37884 14418 37940 14420
rect 37884 14366 37886 14418
rect 37886 14366 37938 14418
rect 37938 14366 37940 14418
rect 37884 14364 37940 14366
rect 37884 13746 37940 13748
rect 37884 13694 37886 13746
rect 37886 13694 37938 13746
rect 37938 13694 37940 13746
rect 37884 13692 37940 13694
rect 37884 12850 37940 12852
rect 37884 12798 37886 12850
rect 37886 12798 37938 12850
rect 37938 12798 37940 12850
rect 37884 12796 37940 12798
rect 37548 12236 37604 12292
rect 37660 12178 37716 12180
rect 37660 12126 37662 12178
rect 37662 12126 37714 12178
rect 37714 12126 37716 12178
rect 37660 12124 37716 12126
rect 37884 11282 37940 11284
rect 37884 11230 37886 11282
rect 37886 11230 37938 11282
rect 37938 11230 37940 11282
rect 37884 11228 37940 11230
rect 37884 10610 37940 10612
rect 37884 10558 37886 10610
rect 37886 10558 37938 10610
rect 37938 10558 37940 10610
rect 37884 10556 37940 10558
rect 37660 9602 37716 9604
rect 37660 9550 37662 9602
rect 37662 9550 37714 9602
rect 37714 9550 37716 9602
rect 37660 9548 37716 9550
rect 38220 14812 38276 14868
rect 38220 14306 38276 14308
rect 38220 14254 38222 14306
rect 38222 14254 38274 14306
rect 38274 14254 38276 14306
rect 38220 14252 38276 14254
rect 38508 14138 38564 14140
rect 38508 14086 38510 14138
rect 38510 14086 38562 14138
rect 38562 14086 38564 14138
rect 38508 14084 38564 14086
rect 38612 14138 38668 14140
rect 38612 14086 38614 14138
rect 38614 14086 38666 14138
rect 38666 14086 38668 14138
rect 38612 14084 38668 14086
rect 38716 14138 38772 14140
rect 38716 14086 38718 14138
rect 38718 14086 38770 14138
rect 38770 14086 38772 14138
rect 38716 14084 38772 14086
rect 38220 13468 38276 13524
rect 38220 12850 38276 12852
rect 38220 12798 38222 12850
rect 38222 12798 38274 12850
rect 38274 12798 38276 12850
rect 38220 12796 38276 12798
rect 38508 12570 38564 12572
rect 38508 12518 38510 12570
rect 38510 12518 38562 12570
rect 38562 12518 38564 12570
rect 38508 12516 38564 12518
rect 38612 12570 38668 12572
rect 38612 12518 38614 12570
rect 38614 12518 38666 12570
rect 38666 12518 38668 12570
rect 38612 12516 38668 12518
rect 38716 12570 38772 12572
rect 38716 12518 38718 12570
rect 38718 12518 38770 12570
rect 38770 12518 38772 12570
rect 38716 12516 38772 12518
rect 38220 12178 38276 12180
rect 38220 12126 38222 12178
rect 38222 12126 38274 12178
rect 38274 12126 38276 12178
rect 38220 12124 38276 12126
rect 38220 11452 38276 11508
rect 38508 11002 38564 11004
rect 38508 10950 38510 11002
rect 38510 10950 38562 11002
rect 38562 10950 38564 11002
rect 38508 10948 38564 10950
rect 38612 11002 38668 11004
rect 38612 10950 38614 11002
rect 38614 10950 38666 11002
rect 38666 10950 38668 11002
rect 38612 10948 38668 10950
rect 38716 11002 38772 11004
rect 38716 10950 38718 11002
rect 38718 10950 38770 11002
rect 38770 10950 38772 11002
rect 38716 10948 38772 10950
rect 38444 10780 38500 10836
rect 38220 10108 38276 10164
rect 38220 9548 38276 9604
rect 38508 9434 38564 9436
rect 38508 9382 38510 9434
rect 38510 9382 38562 9434
rect 38562 9382 38564 9434
rect 38508 9380 38564 9382
rect 38612 9434 38668 9436
rect 38612 9382 38614 9434
rect 38614 9382 38666 9434
rect 38666 9382 38668 9434
rect 38612 9380 38668 9382
rect 38716 9434 38772 9436
rect 38716 9382 38718 9434
rect 38718 9382 38770 9434
rect 38770 9382 38772 9434
rect 38716 9380 38772 9382
rect 38220 8764 38276 8820
rect 37660 8092 37716 8148
rect 37212 7980 37268 8036
rect 38220 8146 38276 8148
rect 38220 8094 38222 8146
rect 38222 8094 38274 8146
rect 38274 8094 38276 8146
rect 38220 8092 38276 8094
rect 38508 7866 38564 7868
rect 38508 7814 38510 7866
rect 38510 7814 38562 7866
rect 38562 7814 38564 7866
rect 38508 7812 38564 7814
rect 38612 7866 38668 7868
rect 38612 7814 38614 7866
rect 38614 7814 38666 7866
rect 38666 7814 38668 7866
rect 38612 7812 38668 7814
rect 38716 7866 38772 7868
rect 38716 7814 38718 7866
rect 38718 7814 38770 7866
rect 38770 7814 38772 7866
rect 38716 7812 38772 7814
rect 37548 7420 37604 7476
rect 37212 7362 37268 7364
rect 37212 7310 37214 7362
rect 37214 7310 37266 7362
rect 37266 7310 37268 7362
rect 37212 7308 37268 7310
rect 37884 7308 37940 7364
rect 38220 6748 38276 6804
rect 37548 6578 37604 6580
rect 37548 6526 37550 6578
rect 37550 6526 37602 6578
rect 37602 6526 37604 6578
rect 37548 6524 37604 6526
rect 38220 6188 38276 6244
rect 38508 6298 38564 6300
rect 38508 6246 38510 6298
rect 38510 6246 38562 6298
rect 38562 6246 38564 6298
rect 38508 6244 38564 6246
rect 38612 6298 38668 6300
rect 38612 6246 38614 6298
rect 38614 6246 38666 6298
rect 38666 6246 38668 6298
rect 38612 6244 38668 6246
rect 38716 6298 38772 6300
rect 38716 6246 38718 6298
rect 38718 6246 38770 6298
rect 38770 6246 38772 6298
rect 38716 6244 38772 6246
rect 37660 5794 37716 5796
rect 37660 5742 37662 5794
rect 37662 5742 37714 5794
rect 37714 5742 37716 5794
rect 37660 5740 37716 5742
rect 38220 5404 38276 5460
rect 37548 5122 37604 5124
rect 37548 5070 37550 5122
rect 37550 5070 37602 5122
rect 37602 5070 37604 5122
rect 37548 5068 37604 5070
rect 37996 5122 38052 5124
rect 37996 5070 37998 5122
rect 37998 5070 38050 5122
rect 38050 5070 38052 5122
rect 37996 5068 38052 5070
rect 38220 4898 38276 4900
rect 38220 4846 38222 4898
rect 38222 4846 38274 4898
rect 38274 4846 38276 4898
rect 38220 4844 38276 4846
rect 38508 4730 38564 4732
rect 38508 4678 38510 4730
rect 38510 4678 38562 4730
rect 38562 4678 38564 4730
rect 38508 4676 38564 4678
rect 38612 4730 38668 4732
rect 38612 4678 38614 4730
rect 38614 4678 38666 4730
rect 38666 4678 38668 4730
rect 38612 4676 38668 4678
rect 38716 4730 38772 4732
rect 38716 4678 38718 4730
rect 38718 4678 38770 4730
rect 38770 4678 38772 4730
rect 38716 4676 38772 4678
rect 37660 4226 37716 4228
rect 37660 4174 37662 4226
rect 37662 4174 37714 4226
rect 37714 4174 37716 4226
rect 37660 4172 37716 4174
rect 38220 4060 38276 4116
rect 37884 3442 37940 3444
rect 37884 3390 37886 3442
rect 37886 3390 37938 3442
rect 37938 3390 37940 3442
rect 37884 3388 37940 3390
rect 38220 3442 38276 3444
rect 38220 3390 38222 3442
rect 38222 3390 38274 3442
rect 38274 3390 38276 3442
rect 38220 3388 38276 3390
rect 29184 3162 29240 3164
rect 29184 3110 29186 3162
rect 29186 3110 29238 3162
rect 29238 3110 29240 3162
rect 29184 3108 29240 3110
rect 29288 3162 29344 3164
rect 29288 3110 29290 3162
rect 29290 3110 29342 3162
rect 29342 3110 29344 3162
rect 29288 3108 29344 3110
rect 29392 3162 29448 3164
rect 29392 3110 29394 3162
rect 29394 3110 29446 3162
rect 29446 3110 29448 3162
rect 29392 3108 29448 3110
rect 38508 3162 38564 3164
rect 38508 3110 38510 3162
rect 38510 3110 38562 3162
rect 38562 3110 38564 3162
rect 38508 3108 38564 3110
rect 38612 3162 38668 3164
rect 38612 3110 38614 3162
rect 38614 3110 38666 3162
rect 38666 3110 38668 3162
rect 38612 3108 38668 3110
rect 38716 3162 38772 3164
rect 38716 3110 38718 3162
rect 38718 3110 38770 3162
rect 38770 3110 38772 3162
rect 38716 3108 38772 3110
rect 37548 2716 37604 2772
<< metal3 >>
rect 39200 37044 40000 37072
rect 37548 36988 40000 37044
rect 37548 36932 37604 36988
rect 39200 36960 40000 36988
rect 37538 36876 37548 36932
rect 37604 36876 37614 36932
rect 5864 36820 5874 36876
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 6138 36820 6148 36876
rect 15188 36820 15198 36876
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15462 36820 15472 36876
rect 24512 36820 24522 36876
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24786 36820 24796 36876
rect 33836 36820 33846 36876
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 34110 36820 34120 36876
rect 24210 36652 24220 36708
rect 24276 36652 25228 36708
rect 25284 36652 25294 36708
rect 24882 36428 24892 36484
rect 24948 36428 25676 36484
rect 25732 36428 26124 36484
rect 26180 36428 26190 36484
rect 39200 36372 40000 36400
rect 23314 36316 23324 36372
rect 23380 36316 25564 36372
rect 25620 36316 25630 36372
rect 36866 36316 36876 36372
rect 36932 36316 40000 36372
rect 39200 36288 40000 36316
rect 36306 36204 36316 36260
rect 36372 36204 38220 36260
rect 38276 36204 38286 36260
rect 10526 36036 10536 36092
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10800 36036 10810 36092
rect 19850 36036 19860 36092
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 20124 36036 20134 36092
rect 29174 36036 29184 36092
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29448 36036 29458 36092
rect 38498 36036 38508 36092
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38772 36036 38782 36092
rect 39200 35700 40000 35728
rect 37090 35644 37100 35700
rect 37156 35644 37996 35700
rect 38052 35644 38062 35700
rect 38322 35644 38332 35700
rect 38388 35644 40000 35700
rect 39200 35616 40000 35644
rect 16034 35308 16044 35364
rect 16100 35308 17276 35364
rect 17332 35308 17342 35364
rect 5864 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6148 35308
rect 15188 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15472 35308
rect 24512 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24796 35308
rect 33836 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34120 35308
rect 37202 35196 37212 35252
rect 37268 35196 39116 35252
rect 39172 35196 39182 35252
rect 39200 35028 40000 35056
rect 38210 34972 38220 35028
rect 38276 34972 40000 35028
rect 39200 34944 40000 34972
rect 10526 34468 10536 34524
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10800 34468 10810 34524
rect 19850 34468 19860 34524
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 20124 34468 20134 34524
rect 29174 34468 29184 34524
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29448 34468 29458 34524
rect 38498 34468 38508 34524
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38772 34468 38782 34524
rect 39200 34356 40000 34384
rect 38434 34300 38444 34356
rect 38500 34300 40000 34356
rect 39200 34272 40000 34300
rect 18498 33964 18508 34020
rect 18564 33964 19292 34020
rect 19348 33964 19358 34020
rect 5864 33684 5874 33740
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 6138 33684 6148 33740
rect 15188 33684 15198 33740
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15462 33684 15472 33740
rect 24512 33684 24522 33740
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24786 33684 24796 33740
rect 33836 33684 33846 33740
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 34110 33684 34120 33740
rect 39200 33684 40000 33712
rect 38210 33628 38220 33684
rect 38276 33628 40000 33684
rect 39200 33600 40000 33628
rect 28578 33180 28588 33236
rect 28644 33180 37884 33236
rect 37940 33180 37950 33236
rect 38210 33068 38220 33124
rect 38276 33068 38948 33124
rect 38892 33012 38948 33068
rect 39200 33012 40000 33040
rect 38892 32956 40000 33012
rect 10526 32900 10536 32956
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10800 32900 10810 32956
rect 19850 32900 19860 32956
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 20124 32900 20134 32956
rect 29174 32900 29184 32956
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29448 32900 29458 32956
rect 38498 32900 38508 32956
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38772 32900 38782 32956
rect 39200 32928 40000 32956
rect 39200 32340 40000 32368
rect 37202 32284 37212 32340
rect 37268 32284 38220 32340
rect 38276 32284 40000 32340
rect 39200 32256 40000 32284
rect 5864 32116 5874 32172
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 6138 32116 6148 32172
rect 15188 32116 15198 32172
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15462 32116 15472 32172
rect 24512 32116 24522 32172
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24786 32116 24796 32172
rect 33836 32116 33846 32172
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 34110 32116 34120 32172
rect 19058 31948 19068 32004
rect 19124 31948 19740 32004
rect 19796 31948 19806 32004
rect 39200 31668 40000 31696
rect 37538 31612 37548 31668
rect 37604 31612 40000 31668
rect 39200 31584 40000 31612
rect 23986 31500 23996 31556
rect 24052 31500 36540 31556
rect 36596 31500 37212 31556
rect 37268 31500 37278 31556
rect 10526 31332 10536 31388
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10800 31332 10810 31388
rect 19850 31332 19860 31388
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 20124 31332 20134 31388
rect 29174 31332 29184 31388
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29448 31332 29458 31388
rect 38498 31332 38508 31388
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38772 31332 38782 31388
rect 39200 30996 40000 31024
rect 38434 30940 38444 30996
rect 38500 30940 40000 30996
rect 39200 30912 40000 30940
rect 27010 30828 27020 30884
rect 27076 30828 37548 30884
rect 37604 30828 37614 30884
rect 5864 30548 5874 30604
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 6138 30548 6148 30604
rect 15188 30548 15198 30604
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15462 30548 15472 30604
rect 24512 30548 24522 30604
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24786 30548 24796 30604
rect 33836 30548 33846 30604
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 34110 30548 34120 30604
rect 39200 30324 40000 30352
rect 38210 30268 38220 30324
rect 38276 30268 40000 30324
rect 39200 30240 40000 30268
rect 19058 30044 19068 30100
rect 19124 30044 20188 30100
rect 20244 30044 20254 30100
rect 10526 29764 10536 29820
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10800 29764 10810 29820
rect 19850 29764 19860 29820
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 20124 29764 20134 29820
rect 29174 29764 29184 29820
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29448 29764 29458 29820
rect 38498 29764 38508 29820
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38772 29764 38782 29820
rect 38210 29708 38220 29764
rect 38276 29708 38286 29764
rect 38220 29652 38276 29708
rect 39200 29652 40000 29680
rect 38220 29596 40000 29652
rect 39200 29568 40000 29596
rect 5864 28980 5874 29036
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 6138 28980 6148 29036
rect 15188 28980 15198 29036
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15462 28980 15472 29036
rect 24512 28980 24522 29036
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24786 28980 24796 29036
rect 33836 28980 33846 29036
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 34110 28980 34120 29036
rect 39200 28980 40000 29008
rect 38210 28924 38220 28980
rect 38276 28924 40000 28980
rect 39200 28896 40000 28924
rect 15698 28588 15708 28644
rect 15764 28588 17612 28644
rect 17668 28588 17678 28644
rect 38210 28364 38220 28420
rect 38276 28364 38948 28420
rect 38892 28308 38948 28364
rect 39200 28308 40000 28336
rect 38892 28252 40000 28308
rect 10526 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10810 28252
rect 19850 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20134 28252
rect 29174 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29458 28252
rect 38498 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38782 28252
rect 39200 28224 40000 28252
rect 30370 27804 30380 27860
rect 30436 27804 37884 27860
rect 37940 27804 37950 27860
rect 39200 27636 40000 27664
rect 38210 27580 38220 27636
rect 38276 27580 40000 27636
rect 39200 27552 40000 27580
rect 5864 27412 5874 27468
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 6138 27412 6148 27468
rect 15188 27412 15198 27468
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15462 27412 15472 27468
rect 24512 27412 24522 27468
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24786 27412 24796 27468
rect 33836 27412 33846 27468
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 34110 27412 34120 27468
rect 27794 27132 27804 27188
rect 27860 27132 37212 27188
rect 37268 27132 37278 27188
rect 37538 27020 37548 27076
rect 37604 27020 39060 27076
rect 39004 26964 39060 27020
rect 39200 26964 40000 26992
rect 39004 26908 40000 26964
rect 39200 26880 40000 26908
rect 1810 26796 1820 26852
rect 1876 26796 2492 26852
rect 2548 26796 2558 26852
rect 10526 26628 10536 26684
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10800 26628 10810 26684
rect 19850 26628 19860 26684
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 20124 26628 20134 26684
rect 29174 26628 29184 26684
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29448 26628 29458 26684
rect 38498 26628 38508 26684
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38772 26628 38782 26684
rect 37202 26572 37212 26628
rect 37268 26572 37660 26628
rect 37716 26572 37726 26628
rect 21410 26460 21420 26516
rect 21476 26460 22316 26516
rect 22372 26460 25900 26516
rect 25956 26460 25966 26516
rect 38098 26348 38108 26404
rect 38164 26348 38174 26404
rect 0 26292 800 26320
rect 38108 26292 38164 26348
rect 39200 26292 40000 26320
rect 0 26236 1820 26292
rect 1876 26236 1886 26292
rect 38108 26236 40000 26292
rect 0 26208 800 26236
rect 39200 26208 40000 26236
rect 37650 26124 37660 26180
rect 37716 26124 38220 26180
rect 38276 26124 38286 26180
rect 5864 25844 5874 25900
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 6138 25844 6148 25900
rect 15188 25844 15198 25900
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15462 25844 15472 25900
rect 24512 25844 24522 25900
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24786 25844 24796 25900
rect 33836 25844 33846 25900
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 34110 25844 34120 25900
rect 0 25620 800 25648
rect 39200 25620 40000 25648
rect 0 25564 1708 25620
rect 1764 25564 1774 25620
rect 38210 25564 38220 25620
rect 38276 25564 40000 25620
rect 0 25536 800 25564
rect 39200 25536 40000 25564
rect 19282 25452 19292 25508
rect 19348 25452 19852 25508
rect 19908 25452 19918 25508
rect 22082 25452 22092 25508
rect 22148 25452 23100 25508
rect 23156 25452 23166 25508
rect 26002 25452 26012 25508
rect 26068 25452 37324 25508
rect 37380 25452 37390 25508
rect 21746 25340 21756 25396
rect 21812 25340 22428 25396
rect 22484 25340 22494 25396
rect 26674 25340 26684 25396
rect 26740 25340 26908 25396
rect 29474 25340 29484 25396
rect 29540 25340 37100 25396
rect 37156 25340 37166 25396
rect 37324 25340 39116 25396
rect 39172 25340 39182 25396
rect 26852 25284 26908 25340
rect 37324 25284 37380 25340
rect 19170 25228 19180 25284
rect 19236 25228 19246 25284
rect 19394 25228 19404 25284
rect 19460 25228 19740 25284
rect 19796 25228 21420 25284
rect 21476 25228 21486 25284
rect 26852 25228 37380 25284
rect 10526 25060 10536 25116
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10800 25060 10810 25116
rect 0 24948 800 24976
rect 0 24892 1820 24948
rect 1876 24892 2492 24948
rect 2548 24892 2558 24948
rect 0 24864 800 24892
rect 19180 24836 19236 25228
rect 19850 25060 19860 25116
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 20124 25060 20134 25116
rect 29174 25060 29184 25116
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29448 25060 29458 25116
rect 38498 25060 38508 25116
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38772 25060 38782 25116
rect 38210 25004 38220 25060
rect 38276 25004 38286 25060
rect 38220 24948 38276 25004
rect 39200 24948 40000 24976
rect 27122 24892 27132 24948
rect 27188 24892 28700 24948
rect 28756 24892 30156 24948
rect 30212 24892 36988 24948
rect 37044 24892 37054 24948
rect 38220 24892 40000 24948
rect 39200 24864 40000 24892
rect 18386 24780 18396 24836
rect 18452 24780 20300 24836
rect 20356 24780 21084 24836
rect 21140 24780 22204 24836
rect 22260 24780 22270 24836
rect 19842 24668 19852 24724
rect 19908 24668 20524 24724
rect 20580 24668 20590 24724
rect 26114 24668 26124 24724
rect 26180 24668 27244 24724
rect 27300 24668 27804 24724
rect 27860 24668 28588 24724
rect 28644 24668 29708 24724
rect 29764 24668 39116 24724
rect 39172 24668 39182 24724
rect 17602 24444 17612 24500
rect 17668 24444 18620 24500
rect 18676 24444 19516 24500
rect 19572 24444 19582 24500
rect 27570 24444 27580 24500
rect 27636 24444 28028 24500
rect 28084 24444 28364 24500
rect 28420 24444 28924 24500
rect 28980 24444 28990 24500
rect 0 24276 800 24304
rect 5864 24276 5874 24332
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 6138 24276 6148 24332
rect 15188 24276 15198 24332
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15462 24276 15472 24332
rect 24512 24276 24522 24332
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24786 24276 24796 24332
rect 33836 24276 33846 24332
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 34110 24276 34120 24332
rect 39200 24276 40000 24304
rect 0 24220 1708 24276
rect 1764 24220 1774 24276
rect 38210 24220 38220 24276
rect 38276 24220 40000 24276
rect 0 24192 800 24220
rect 39200 24192 40000 24220
rect 22754 24108 22764 24164
rect 22820 24108 23772 24164
rect 23828 24108 23838 24164
rect 24658 24108 24668 24164
rect 24724 24108 25452 24164
rect 25508 24108 25518 24164
rect 26852 24108 28812 24164
rect 28868 24108 29148 24164
rect 29204 24108 37324 24164
rect 37380 24108 37390 24164
rect 15026 23996 15036 24052
rect 15092 23996 16604 24052
rect 16660 23996 17388 24052
rect 17444 23996 17454 24052
rect 26852 23940 26908 24108
rect 17042 23884 17052 23940
rect 17108 23884 18844 23940
rect 18900 23884 20636 23940
rect 20692 23884 20702 23940
rect 25778 23884 25788 23940
rect 25844 23884 26236 23940
rect 26292 23884 26908 23940
rect 24882 23772 24892 23828
rect 24948 23772 25340 23828
rect 25396 23772 27356 23828
rect 27412 23772 27422 23828
rect 28578 23772 28588 23828
rect 28644 23772 39004 23828
rect 39060 23772 39070 23828
rect 1698 23660 1708 23716
rect 1764 23660 1774 23716
rect 26852 23660 27132 23716
rect 27188 23660 27198 23716
rect 38210 23660 38220 23716
rect 38276 23660 38948 23716
rect 0 23604 800 23632
rect 1708 23604 1764 23660
rect 0 23548 1764 23604
rect 20626 23548 20636 23604
rect 20692 23548 21812 23604
rect 0 23520 800 23548
rect 10526 23492 10536 23548
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10800 23492 10810 23548
rect 19850 23492 19860 23548
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 20124 23492 20134 23548
rect 21756 23492 21812 23548
rect 26852 23492 26908 23660
rect 38892 23604 38948 23660
rect 39200 23604 40000 23632
rect 38892 23548 40000 23604
rect 29174 23492 29184 23548
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29448 23492 29458 23548
rect 38498 23492 38508 23548
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38772 23492 38782 23548
rect 39200 23520 40000 23548
rect 21746 23436 21756 23492
rect 21812 23436 21822 23492
rect 25218 23436 25228 23492
rect 25284 23436 26012 23492
rect 26068 23436 26908 23492
rect 31266 23436 31276 23492
rect 31332 23436 37548 23492
rect 37604 23436 37614 23492
rect 19740 23324 20860 23380
rect 20916 23324 20926 23380
rect 23874 23324 23884 23380
rect 23940 23324 37436 23380
rect 37492 23324 37502 23380
rect 19740 23268 19796 23324
rect 19730 23212 19740 23268
rect 19796 23212 19806 23268
rect 21074 23212 21084 23268
rect 21140 23212 22092 23268
rect 22148 23212 22158 23268
rect 27346 23212 27356 23268
rect 27412 23212 28476 23268
rect 28532 23212 28924 23268
rect 28980 23212 38892 23268
rect 38948 23212 38958 23268
rect 2034 23100 2044 23156
rect 2100 23100 15596 23156
rect 15652 23100 15662 23156
rect 20402 23100 20412 23156
rect 20468 23100 21196 23156
rect 21252 23100 21980 23156
rect 22036 23100 22046 23156
rect 26114 23100 26124 23156
rect 26180 23100 37884 23156
rect 37940 23100 37950 23156
rect 0 22932 800 22960
rect 39200 22932 40000 22960
rect 0 22876 1708 22932
rect 1764 22876 1774 22932
rect 38210 22876 38220 22932
rect 38276 22876 40000 22932
rect 0 22848 800 22876
rect 39200 22848 40000 22876
rect 5864 22708 5874 22764
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 6138 22708 6148 22764
rect 15188 22708 15198 22764
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15462 22708 15472 22764
rect 24512 22708 24522 22764
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24786 22708 24796 22764
rect 33836 22708 33846 22764
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 34110 22708 34120 22764
rect 16706 22540 16716 22596
rect 16772 22540 17388 22596
rect 17444 22540 17454 22596
rect 19954 22540 19964 22596
rect 20020 22540 20300 22596
rect 20356 22540 20366 22596
rect 23202 22540 23212 22596
rect 23268 22540 37772 22596
rect 37828 22540 37838 22596
rect 17154 22428 17164 22484
rect 17220 22428 18844 22484
rect 18900 22428 21420 22484
rect 21476 22428 21486 22484
rect 17602 22316 17612 22372
rect 17668 22316 18620 22372
rect 18676 22316 19628 22372
rect 19684 22316 19694 22372
rect 30482 22316 30492 22372
rect 30548 22316 37996 22372
rect 38052 22316 38062 22372
rect 0 22260 800 22288
rect 39200 22260 40000 22288
rect 0 22204 1708 22260
rect 1764 22204 1774 22260
rect 2034 22204 2044 22260
rect 2100 22204 14700 22260
rect 14756 22204 14766 22260
rect 20290 22204 20300 22260
rect 20356 22204 21532 22260
rect 21588 22204 21598 22260
rect 22418 22204 22428 22260
rect 22484 22204 23548 22260
rect 23604 22204 23614 22260
rect 29250 22204 29260 22260
rect 29316 22204 29820 22260
rect 29876 22204 29886 22260
rect 30594 22204 30604 22260
rect 30660 22204 36428 22260
rect 36484 22204 36494 22260
rect 38210 22204 38220 22260
rect 38276 22204 40000 22260
rect 0 22176 800 22204
rect 39200 22176 40000 22204
rect 30258 21980 30268 22036
rect 30324 21980 37884 22036
rect 37940 21980 37950 22036
rect 10526 21924 10536 21980
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10800 21924 10810 21980
rect 19850 21924 19860 21980
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 20124 21924 20134 21980
rect 29174 21924 29184 21980
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29448 21924 29458 21980
rect 38498 21924 38508 21980
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38772 21924 38782 21980
rect 29586 21868 29596 21924
rect 29652 21868 30940 21924
rect 30996 21868 31006 21924
rect 924 21756 2380 21812
rect 2436 21756 2446 21812
rect 23090 21756 23100 21812
rect 23156 21756 37100 21812
rect 37156 21756 37166 21812
rect 0 21588 800 21616
rect 924 21588 980 21756
rect 8372 21644 12348 21700
rect 12404 21644 12414 21700
rect 24434 21644 24444 21700
rect 24500 21644 25228 21700
rect 25284 21644 26348 21700
rect 26404 21644 26414 21700
rect 26786 21644 26796 21700
rect 26852 21644 27468 21700
rect 27524 21644 29148 21700
rect 29204 21644 29708 21700
rect 29764 21644 29774 21700
rect 8372 21588 8428 21644
rect 39200 21588 40000 21616
rect 0 21532 980 21588
rect 2034 21532 2044 21588
rect 2100 21532 8428 21588
rect 19170 21532 19180 21588
rect 19236 21532 20412 21588
rect 20468 21532 21420 21588
rect 21476 21532 21486 21588
rect 23650 21532 23660 21588
rect 23716 21532 24332 21588
rect 24388 21532 25564 21588
rect 25620 21532 26572 21588
rect 26628 21532 26638 21588
rect 27346 21532 27356 21588
rect 27412 21532 29036 21588
rect 29092 21532 29102 21588
rect 37538 21532 37548 21588
rect 37604 21532 40000 21588
rect 0 21504 800 21532
rect 39200 21504 40000 21532
rect 19730 21420 19740 21476
rect 19796 21420 20300 21476
rect 20356 21420 20366 21476
rect 28690 21420 28700 21476
rect 28756 21420 30380 21476
rect 30436 21420 30446 21476
rect 1922 21308 1932 21364
rect 1988 21308 10332 21364
rect 10388 21308 10398 21364
rect 24658 21308 24668 21364
rect 24724 21308 25452 21364
rect 25508 21308 27244 21364
rect 27300 21308 27310 21364
rect 5864 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6148 21196
rect 15188 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15472 21196
rect 24512 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24796 21196
rect 29260 21140 29316 21420
rect 33836 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34120 21196
rect 29250 21084 29260 21140
rect 29316 21084 29326 21140
rect 2706 20972 2716 21028
rect 2772 20972 16828 21028
rect 16884 20972 16894 21028
rect 24434 20972 24444 21028
rect 24500 20972 37660 21028
rect 37716 20972 37726 21028
rect 0 20916 800 20944
rect 39200 20916 40000 20944
rect 0 20860 1708 20916
rect 1764 20860 1774 20916
rect 2482 20860 2492 20916
rect 2548 20860 17948 20916
rect 18004 20860 18014 20916
rect 23538 20860 23548 20916
rect 23604 20860 37212 20916
rect 37268 20860 37278 20916
rect 38210 20860 38220 20916
rect 38276 20860 40000 20916
rect 0 20832 800 20860
rect 39200 20832 40000 20860
rect 14690 20748 14700 20804
rect 14756 20748 15596 20804
rect 15652 20748 15662 20804
rect 20178 20748 20188 20804
rect 20244 20748 20636 20804
rect 20692 20748 20702 20804
rect 26852 20748 29260 20804
rect 29316 20748 29326 20804
rect 26852 20692 26908 20748
rect 2146 20636 2156 20692
rect 2212 20636 11116 20692
rect 11172 20636 11182 20692
rect 14130 20636 14140 20692
rect 14196 20636 15260 20692
rect 15316 20636 16268 20692
rect 16324 20636 18844 20692
rect 18900 20636 18910 20692
rect 21634 20636 21644 20692
rect 21700 20636 22540 20692
rect 22596 20636 22606 20692
rect 25330 20636 25340 20692
rect 25396 20636 25788 20692
rect 25844 20636 26908 20692
rect 28130 20636 28140 20692
rect 28196 20636 38108 20692
rect 38164 20636 38174 20692
rect 1698 20524 1708 20580
rect 1764 20524 1774 20580
rect 10770 20524 10780 20580
rect 10836 20524 11788 20580
rect 11844 20524 12012 20580
rect 12068 20524 13580 20580
rect 13636 20524 13646 20580
rect 19058 20524 19068 20580
rect 19124 20524 19628 20580
rect 19684 20524 19694 20580
rect 20738 20524 20748 20580
rect 20804 20524 21756 20580
rect 21812 20524 21822 20580
rect 26674 20524 26684 20580
rect 26740 20524 37884 20580
rect 37940 20524 37950 20580
rect 0 20244 800 20272
rect 1708 20244 1764 20524
rect 10526 20356 10536 20412
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10800 20356 10810 20412
rect 19850 20356 19860 20412
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 20124 20356 20134 20412
rect 29174 20356 29184 20412
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29448 20356 29458 20412
rect 38498 20356 38508 20412
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38772 20356 38782 20412
rect 39200 20244 40000 20272
rect 0 20188 1764 20244
rect 2034 20188 2044 20244
rect 2100 20188 11788 20244
rect 11844 20188 11854 20244
rect 15092 20188 15372 20244
rect 15428 20188 16156 20244
rect 16212 20188 16222 20244
rect 38434 20188 38444 20244
rect 38500 20188 40000 20244
rect 0 20160 800 20188
rect 15092 20132 15148 20188
rect 39200 20160 40000 20188
rect 2594 20076 2604 20132
rect 2660 20076 10780 20132
rect 10836 20076 11676 20132
rect 11732 20076 12124 20132
rect 12180 20076 12190 20132
rect 14242 20076 14252 20132
rect 14308 20076 15148 20132
rect 19954 20076 19964 20132
rect 20020 20076 22092 20132
rect 22148 20076 23996 20132
rect 24052 20076 24062 20132
rect 28914 20076 28924 20132
rect 28980 20076 37884 20132
rect 37940 20076 37950 20132
rect 2034 19964 2044 20020
rect 2100 19964 15820 20020
rect 15876 19964 15886 20020
rect 18386 19964 18396 20020
rect 18452 19964 19628 20020
rect 19684 19964 19694 20020
rect 21410 19964 21420 20020
rect 21476 19964 22652 20020
rect 22708 19964 22718 20020
rect 28242 19964 28252 20020
rect 28308 19964 37996 20020
rect 38052 19964 38062 20020
rect 13570 19852 13580 19908
rect 13636 19852 14924 19908
rect 14980 19852 14990 19908
rect 20626 19852 20636 19908
rect 20692 19852 26012 19908
rect 26068 19852 26908 19908
rect 26964 19852 26974 19908
rect 11890 19740 11900 19796
rect 11956 19740 12796 19796
rect 12852 19740 17612 19796
rect 17668 19740 18172 19796
rect 18228 19740 18238 19796
rect 21074 19740 21084 19796
rect 21140 19740 26684 19796
rect 26740 19740 26750 19796
rect 19506 19628 19516 19684
rect 19572 19628 22428 19684
rect 22484 19628 22494 19684
rect 0 19572 800 19600
rect 5864 19572 5874 19628
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 6138 19572 6148 19628
rect 15188 19572 15198 19628
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15462 19572 15472 19628
rect 0 19516 1708 19572
rect 1764 19516 1774 19572
rect 0 19488 800 19516
rect 22428 19460 22484 19628
rect 24512 19572 24522 19628
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24786 19572 24796 19628
rect 33836 19572 33846 19628
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 34110 19572 34120 19628
rect 39200 19572 40000 19600
rect 38210 19516 38220 19572
rect 38276 19516 40000 19572
rect 39200 19488 40000 19516
rect 2034 19404 2044 19460
rect 2100 19404 16996 19460
rect 22428 19404 28364 19460
rect 28420 19404 28430 19460
rect 11666 19292 11676 19348
rect 11732 19292 13580 19348
rect 13636 19292 14028 19348
rect 14084 19292 14094 19348
rect 2818 19180 2828 19236
rect 2884 19180 14924 19236
rect 14980 19180 14990 19236
rect 14578 19068 14588 19124
rect 14644 19068 15932 19124
rect 15988 19068 15998 19124
rect 16940 19012 16996 19404
rect 21522 19292 21532 19348
rect 21588 19292 22540 19348
rect 22596 19292 22606 19348
rect 22978 19292 22988 19348
rect 23044 19292 23436 19348
rect 23492 19292 26012 19348
rect 26068 19292 26078 19348
rect 21858 19180 21868 19236
rect 21924 19180 37884 19236
rect 37940 19180 37950 19236
rect 19730 19068 19740 19124
rect 19796 19068 21084 19124
rect 21140 19068 21150 19124
rect 23090 19068 23100 19124
rect 23156 19068 23996 19124
rect 24052 19068 24062 19124
rect 24322 19068 24332 19124
rect 24388 19068 25340 19124
rect 25396 19068 25406 19124
rect 27234 19068 27244 19124
rect 27300 19068 28364 19124
rect 28420 19068 28430 19124
rect 29026 19068 29036 19124
rect 29092 19068 29596 19124
rect 29652 19068 30156 19124
rect 30212 19068 30716 19124
rect 30772 19068 30782 19124
rect 1698 18956 1708 19012
rect 1764 18956 1774 19012
rect 16930 18956 16940 19012
rect 16996 18956 17006 19012
rect 25666 18956 25676 19012
rect 25732 18956 25742 19012
rect 26338 18956 26348 19012
rect 26404 18956 28700 19012
rect 28756 18956 28766 19012
rect 28924 18956 29484 19012
rect 29540 18956 30044 19012
rect 30100 18956 30604 19012
rect 30660 18956 30670 19012
rect 38210 18956 38220 19012
rect 38276 18956 38948 19012
rect 0 18900 800 18928
rect 1708 18900 1764 18956
rect 0 18844 1764 18900
rect 0 18816 800 18844
rect 10526 18788 10536 18844
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10800 18788 10810 18844
rect 19850 18788 19860 18844
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 20124 18788 20134 18844
rect 25676 18788 25732 18956
rect 28924 18788 28980 18956
rect 38892 18900 38948 18956
rect 39200 18900 40000 18928
rect 38892 18844 40000 18900
rect 29174 18788 29184 18844
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29448 18788 29458 18844
rect 38498 18788 38508 18844
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38772 18788 38782 18844
rect 39200 18816 40000 18844
rect 25676 18732 28924 18788
rect 28980 18732 28990 18788
rect 27906 18620 27916 18676
rect 27972 18620 28588 18676
rect 28644 18620 28654 18676
rect 30930 18620 30940 18676
rect 30996 18620 31006 18676
rect 30940 18564 30996 18620
rect 15810 18508 15820 18564
rect 15876 18508 18396 18564
rect 18452 18508 19068 18564
rect 19124 18508 19134 18564
rect 26562 18508 26572 18564
rect 26628 18508 27356 18564
rect 27412 18508 27422 18564
rect 28354 18508 28364 18564
rect 28420 18508 29596 18564
rect 29652 18508 30268 18564
rect 30324 18508 30996 18564
rect 2034 18396 2044 18452
rect 2100 18396 8428 18452
rect 12114 18396 12124 18452
rect 12180 18396 13804 18452
rect 13860 18396 13870 18452
rect 14018 18396 14028 18452
rect 14084 18396 15372 18452
rect 15428 18396 16044 18452
rect 16100 18396 16110 18452
rect 16370 18396 16380 18452
rect 16436 18396 17500 18452
rect 17556 18396 17566 18452
rect 17826 18396 17836 18452
rect 17892 18396 18508 18452
rect 18564 18396 19516 18452
rect 19572 18396 19582 18452
rect 20178 18396 20188 18452
rect 20244 18396 21084 18452
rect 21140 18396 21756 18452
rect 21812 18396 21822 18452
rect 26450 18396 26460 18452
rect 26516 18396 27468 18452
rect 27524 18396 27534 18452
rect 37874 18396 37884 18452
rect 37940 18396 37950 18452
rect 8372 18340 8428 18396
rect 8372 18284 14924 18340
rect 14980 18284 14990 18340
rect 15922 18284 15932 18340
rect 15988 18284 16492 18340
rect 16548 18284 17724 18340
rect 17780 18284 18844 18340
rect 18900 18284 18910 18340
rect 20850 18284 20860 18340
rect 20916 18284 21980 18340
rect 22036 18284 22764 18340
rect 22820 18284 22830 18340
rect 28354 18284 28364 18340
rect 28420 18284 29932 18340
rect 29988 18284 30492 18340
rect 30548 18284 31724 18340
rect 31780 18284 37436 18340
rect 37492 18284 37502 18340
rect 0 18228 800 18256
rect 37884 18228 37940 18396
rect 39200 18228 40000 18256
rect 0 18172 1708 18228
rect 1764 18172 1774 18228
rect 11890 18172 11900 18228
rect 11956 18172 12796 18228
rect 12852 18172 16828 18228
rect 16884 18172 16894 18228
rect 19842 18172 19852 18228
rect 19908 18172 20300 18228
rect 20356 18172 22988 18228
rect 23044 18172 23054 18228
rect 24434 18172 24444 18228
rect 24500 18172 37940 18228
rect 38210 18172 38220 18228
rect 38276 18172 40000 18228
rect 0 18144 800 18172
rect 39200 18144 40000 18172
rect 5864 18004 5874 18060
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 6138 18004 6148 18060
rect 15188 18004 15198 18060
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15462 18004 15472 18060
rect 24512 18004 24522 18060
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24786 18004 24796 18060
rect 33836 18004 33846 18060
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 34110 18004 34120 18060
rect 2034 17836 2044 17892
rect 2100 17836 12572 17892
rect 12628 17836 12638 17892
rect 14130 17836 14140 17892
rect 14196 17836 16268 17892
rect 16324 17836 18172 17892
rect 18228 17836 18238 17892
rect 2706 17612 2716 17668
rect 2772 17612 10892 17668
rect 10948 17612 10958 17668
rect 14578 17612 14588 17668
rect 14644 17612 15148 17668
rect 15204 17612 15214 17668
rect 20748 17612 37884 17668
rect 37940 17612 37950 17668
rect 0 17556 800 17584
rect 0 17500 1708 17556
rect 1764 17500 3164 17556
rect 3220 17500 3230 17556
rect 12898 17500 12908 17556
rect 12964 17500 13692 17556
rect 13748 17500 13758 17556
rect 0 17472 800 17500
rect 20748 17444 20804 17612
rect 39200 17556 40000 17584
rect 22082 17500 22092 17556
rect 22148 17500 22652 17556
rect 22708 17500 23100 17556
rect 23156 17500 23660 17556
rect 23716 17500 24332 17556
rect 24388 17500 24398 17556
rect 24770 17500 24780 17556
rect 24836 17500 37212 17556
rect 37268 17500 37278 17556
rect 38210 17500 38220 17556
rect 38276 17500 40000 17556
rect 39200 17472 40000 17500
rect 2034 17388 2044 17444
rect 2100 17388 15036 17444
rect 15092 17388 16380 17444
rect 16436 17388 16604 17444
rect 16660 17388 18284 17444
rect 18340 17388 18350 17444
rect 20738 17388 20748 17444
rect 20804 17388 20814 17444
rect 27122 17388 27132 17444
rect 27188 17388 28476 17444
rect 28532 17388 29260 17444
rect 29316 17388 30380 17444
rect 30436 17388 30716 17444
rect 30772 17388 30782 17444
rect 10526 17220 10536 17276
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10800 17220 10810 17276
rect 19850 17220 19860 17276
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 20124 17220 20134 17276
rect 29174 17220 29184 17276
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29448 17220 29458 17276
rect 38498 17220 38508 17276
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38772 17220 38782 17276
rect 1260 17052 2380 17108
rect 2436 17052 2446 17108
rect 18274 17052 18284 17108
rect 18340 17052 25452 17108
rect 25508 17052 25518 17108
rect 26562 17052 26572 17108
rect 26628 17052 26908 17108
rect 0 16884 800 16912
rect 1260 16884 1316 17052
rect 26852 16996 26908 17052
rect 2258 16940 2268 16996
rect 2324 16940 11340 16996
rect 11396 16940 12908 16996
rect 12964 16940 14364 16996
rect 14420 16940 14430 16996
rect 20290 16940 20300 16996
rect 20356 16940 21084 16996
rect 21140 16940 21532 16996
rect 21588 16940 21598 16996
rect 26852 16940 37884 16996
rect 37940 16940 37950 16996
rect 39200 16884 40000 16912
rect 0 16828 1316 16884
rect 2034 16828 2044 16884
rect 2100 16828 12572 16884
rect 12628 16828 12638 16884
rect 15922 16828 15932 16884
rect 15988 16828 16716 16884
rect 16772 16828 17612 16884
rect 17668 16828 17678 16884
rect 19394 16828 19404 16884
rect 19460 16828 20412 16884
rect 20468 16828 22876 16884
rect 22932 16828 23324 16884
rect 23380 16828 24276 16884
rect 26450 16828 26460 16884
rect 26516 16828 26908 16884
rect 26964 16828 29820 16884
rect 29876 16828 30492 16884
rect 30548 16828 30558 16884
rect 30706 16828 30716 16884
rect 30772 16828 32396 16884
rect 32452 16828 37100 16884
rect 37156 16828 37166 16884
rect 37538 16828 37548 16884
rect 37604 16828 40000 16884
rect 0 16800 800 16828
rect 24220 16660 24276 16828
rect 39200 16800 40000 16828
rect 25554 16716 25564 16772
rect 25620 16716 26236 16772
rect 26292 16716 27020 16772
rect 27076 16716 27468 16772
rect 27524 16716 27534 16772
rect 24210 16604 24220 16660
rect 24276 16604 24286 16660
rect 29138 16604 29148 16660
rect 29204 16604 30044 16660
rect 30100 16604 30940 16660
rect 30996 16604 31006 16660
rect 5864 16436 5874 16492
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 6138 16436 6148 16492
rect 15188 16436 15198 16492
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15462 16436 15472 16492
rect 24512 16436 24522 16492
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24786 16436 24796 16492
rect 33836 16436 33846 16492
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 34110 16436 34120 16492
rect 18610 16268 18620 16324
rect 18676 16268 19516 16324
rect 19572 16268 20524 16324
rect 20580 16268 21532 16324
rect 21588 16268 21598 16324
rect 0 16212 800 16240
rect 39200 16212 40000 16240
rect 0 16156 1708 16212
rect 1764 16156 1774 16212
rect 21298 16156 21308 16212
rect 21364 16156 23100 16212
rect 23156 16156 23166 16212
rect 24210 16156 24220 16212
rect 24276 16156 25900 16212
rect 25956 16156 25966 16212
rect 38210 16156 38220 16212
rect 38276 16156 40000 16212
rect 0 16128 800 16156
rect 39200 16128 40000 16156
rect 18386 16044 18396 16100
rect 18452 16044 20188 16100
rect 20244 16044 20254 16100
rect 22754 16044 22764 16100
rect 22820 16044 23548 16100
rect 23604 16044 24444 16100
rect 24500 16044 24510 16100
rect 31938 16044 31948 16100
rect 32004 16044 37884 16100
rect 37940 16044 37950 16100
rect 14242 15932 14252 15988
rect 14308 15932 16716 15988
rect 16772 15932 18508 15988
rect 18564 15932 18574 15988
rect 18722 15932 18732 15988
rect 18788 15932 20076 15988
rect 20132 15932 20142 15988
rect 24770 15932 24780 15988
rect 24836 15932 25116 15988
rect 25172 15932 25182 15988
rect 1698 15820 1708 15876
rect 1764 15820 1774 15876
rect 18946 15820 18956 15876
rect 19012 15820 20412 15876
rect 20468 15820 20478 15876
rect 21858 15820 21868 15876
rect 21924 15820 24332 15876
rect 24388 15820 24398 15876
rect 0 15540 800 15568
rect 1708 15540 1764 15820
rect 10526 15652 10536 15708
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10800 15652 10810 15708
rect 19850 15652 19860 15708
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 20124 15652 20134 15708
rect 29174 15652 29184 15708
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29448 15652 29458 15708
rect 38498 15652 38508 15708
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38772 15652 38782 15708
rect 39200 15540 40000 15568
rect 0 15484 1764 15540
rect 38434 15484 38444 15540
rect 38500 15484 40000 15540
rect 0 15456 800 15484
rect 39200 15456 40000 15484
rect 20178 15372 20188 15428
rect 20244 15372 21868 15428
rect 21924 15372 21934 15428
rect 2034 15260 2044 15316
rect 2100 15260 12124 15316
rect 12180 15260 12190 15316
rect 23762 15260 23772 15316
rect 23828 15260 25228 15316
rect 25284 15260 25294 15316
rect 27122 15260 27132 15316
rect 27188 15260 28028 15316
rect 28084 15260 28094 15316
rect 28466 15260 28476 15316
rect 28532 15260 29820 15316
rect 29876 15260 30156 15316
rect 30212 15260 31500 15316
rect 31556 15260 37996 15316
rect 38052 15260 38062 15316
rect 2146 15148 2156 15204
rect 2212 15148 14700 15204
rect 14756 15148 15596 15204
rect 15652 15148 15662 15204
rect 23202 15148 23212 15204
rect 23268 15148 24220 15204
rect 24276 15148 24286 15204
rect 27346 15148 27356 15204
rect 27412 15148 28924 15204
rect 28980 15148 37772 15204
rect 37828 15148 37838 15204
rect 19058 15036 19068 15092
rect 19124 15036 19740 15092
rect 19796 15036 19806 15092
rect 0 14868 800 14896
rect 5864 14868 5874 14924
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 6138 14868 6148 14924
rect 15188 14868 15198 14924
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15462 14868 15472 14924
rect 24512 14868 24522 14924
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24786 14868 24796 14924
rect 33836 14868 33846 14924
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 34110 14868 34120 14924
rect 39200 14868 40000 14896
rect 0 14812 1708 14868
rect 1764 14812 1774 14868
rect 38210 14812 38220 14868
rect 38276 14812 40000 14868
rect 0 14784 800 14812
rect 39200 14784 40000 14812
rect 16818 14700 16828 14756
rect 16884 14700 18284 14756
rect 18340 14700 19404 14756
rect 19460 14700 19470 14756
rect 37436 14588 37884 14644
rect 37940 14588 37950 14644
rect 15698 14476 15708 14532
rect 15764 14476 19068 14532
rect 19124 14476 19134 14532
rect 25554 14476 25564 14532
rect 25620 14476 37212 14532
rect 37268 14476 37278 14532
rect 37436 14420 37492 14588
rect 17042 14364 17052 14420
rect 17108 14364 18060 14420
rect 18116 14364 19180 14420
rect 19236 14364 19246 14420
rect 27458 14364 27468 14420
rect 27524 14364 37492 14420
rect 37874 14364 37884 14420
rect 37940 14364 37950 14420
rect 37884 14308 37940 14364
rect 2034 14252 2044 14308
rect 2100 14252 14924 14308
rect 14980 14252 15484 14308
rect 15540 14252 15550 14308
rect 16146 14252 16156 14308
rect 16212 14252 19068 14308
rect 19124 14252 19134 14308
rect 29810 14252 29820 14308
rect 29876 14252 37940 14308
rect 38210 14252 38220 14308
rect 38276 14252 38948 14308
rect 0 14196 800 14224
rect 38892 14196 38948 14252
rect 39200 14196 40000 14224
rect 0 14140 1708 14196
rect 1764 14140 2492 14196
rect 2548 14140 2558 14196
rect 38892 14140 40000 14196
rect 0 14112 800 14140
rect 10526 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10810 14140
rect 19850 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20134 14140
rect 29174 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29458 14140
rect 38498 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38782 14140
rect 39200 14112 40000 14140
rect 17602 13804 17612 13860
rect 17668 13804 18508 13860
rect 18564 13804 19964 13860
rect 20020 13804 23548 13860
rect 23604 13804 23614 13860
rect 17612 13692 18284 13748
rect 18340 13692 18350 13748
rect 23314 13692 23324 13748
rect 23380 13692 23884 13748
rect 23940 13692 23950 13748
rect 24210 13692 24220 13748
rect 24276 13692 25228 13748
rect 25284 13692 25294 13748
rect 28130 13692 28140 13748
rect 28196 13692 37884 13748
rect 37940 13692 37950 13748
rect 17612 13636 17668 13692
rect 14802 13580 14812 13636
rect 14868 13580 16828 13636
rect 16884 13580 17388 13636
rect 17444 13580 17454 13636
rect 17602 13580 17612 13636
rect 17668 13580 17678 13636
rect 18050 13580 18060 13636
rect 18116 13580 18126 13636
rect 21858 13580 21868 13636
rect 21924 13580 22316 13636
rect 22372 13580 22764 13636
rect 22820 13580 24668 13636
rect 24724 13580 25900 13636
rect 25956 13580 25966 13636
rect 0 13524 800 13552
rect 18060 13524 18116 13580
rect 39200 13524 40000 13552
rect 0 13468 1708 13524
rect 1764 13468 2492 13524
rect 2548 13468 2558 13524
rect 17612 13468 18116 13524
rect 38210 13468 38220 13524
rect 38276 13468 40000 13524
rect 0 13440 800 13468
rect 17612 13412 17668 13468
rect 39200 13440 40000 13468
rect 17602 13356 17612 13412
rect 17668 13356 17678 13412
rect 5864 13300 5874 13356
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 6138 13300 6148 13356
rect 15188 13300 15198 13356
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15462 13300 15472 13356
rect 24512 13300 24522 13356
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24786 13300 24796 13356
rect 33836 13300 33846 13356
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 34110 13300 34120 13356
rect 20626 12908 20636 12964
rect 20692 12908 21980 12964
rect 22036 12908 22046 12964
rect 0 12852 800 12880
rect 39200 12852 40000 12880
rect 0 12796 1708 12852
rect 1764 12796 2492 12852
rect 2548 12796 2558 12852
rect 31042 12796 31052 12852
rect 31108 12796 37884 12852
rect 37940 12796 37950 12852
rect 38210 12796 38220 12852
rect 38276 12796 40000 12852
rect 0 12768 800 12796
rect 39200 12768 40000 12796
rect 16594 12684 16604 12740
rect 16660 12684 17388 12740
rect 17444 12684 17454 12740
rect 20178 12684 20188 12740
rect 20244 12684 21420 12740
rect 21476 12684 23660 12740
rect 23716 12684 24444 12740
rect 24500 12684 26572 12740
rect 26628 12684 26638 12740
rect 10526 12516 10536 12572
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10800 12516 10810 12572
rect 19850 12516 19860 12572
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 20124 12516 20134 12572
rect 29174 12516 29184 12572
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29448 12516 29458 12572
rect 38498 12516 38508 12572
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38772 12516 38782 12572
rect 37538 12236 37548 12292
rect 37604 12236 38500 12292
rect 38444 12180 38500 12236
rect 39200 12180 40000 12208
rect 37650 12124 37660 12180
rect 37716 12124 38220 12180
rect 38276 12124 38286 12180
rect 38444 12124 40000 12180
rect 39200 12096 40000 12124
rect 17938 11788 17948 11844
rect 18004 11788 18844 11844
rect 18900 11788 18910 11844
rect 22754 11788 22764 11844
rect 22820 11788 24108 11844
rect 24164 11788 24174 11844
rect 5864 11732 5874 11788
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 6138 11732 6148 11788
rect 15188 11732 15198 11788
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15462 11732 15472 11788
rect 24512 11732 24522 11788
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24786 11732 24796 11788
rect 33836 11732 33846 11788
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 34110 11732 34120 11788
rect 39200 11508 40000 11536
rect 38210 11452 38220 11508
rect 38276 11452 40000 11508
rect 39200 11424 40000 11452
rect 25442 11228 25452 11284
rect 25508 11228 37884 11284
rect 37940 11228 37950 11284
rect 10526 10948 10536 11004
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10800 10948 10810 11004
rect 19850 10948 19860 11004
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 20124 10948 20134 11004
rect 29174 10948 29184 11004
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29448 10948 29458 11004
rect 38498 10948 38508 11004
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38772 10948 38782 11004
rect 30818 10892 30828 10948
rect 30884 10892 37324 10948
rect 37380 10892 37390 10948
rect 39200 10836 40000 10864
rect 38434 10780 38444 10836
rect 38500 10780 40000 10836
rect 39200 10752 40000 10780
rect 27906 10556 27916 10612
rect 27972 10556 37884 10612
rect 37940 10556 37950 10612
rect 5864 10164 5874 10220
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 6138 10164 6148 10220
rect 15188 10164 15198 10220
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15462 10164 15472 10220
rect 24512 10164 24522 10220
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24786 10164 24796 10220
rect 33836 10164 33846 10220
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 34110 10164 34120 10220
rect 39200 10164 40000 10192
rect 38210 10108 38220 10164
rect 38276 10108 40000 10164
rect 39200 10080 40000 10108
rect 37650 9548 37660 9604
rect 37716 9548 38220 9604
rect 38276 9548 38948 9604
rect 38892 9492 38948 9548
rect 39200 9492 40000 9520
rect 38892 9436 40000 9492
rect 10526 9380 10536 9436
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10800 9380 10810 9436
rect 19850 9380 19860 9436
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 20124 9380 20134 9436
rect 29174 9380 29184 9436
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29448 9380 29458 9436
rect 38498 9380 38508 9436
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38772 9380 38782 9436
rect 39200 9408 40000 9436
rect 39200 8820 40000 8848
rect 38210 8764 38220 8820
rect 38276 8764 40000 8820
rect 39200 8736 40000 8764
rect 5864 8596 5874 8652
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 6138 8596 6148 8652
rect 15188 8596 15198 8652
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15462 8596 15472 8652
rect 24512 8596 24522 8652
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24786 8596 24796 8652
rect 33836 8596 33846 8652
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 34110 8596 34120 8652
rect 39200 8148 40000 8176
rect 37650 8092 37660 8148
rect 37716 8092 38220 8148
rect 38276 8092 40000 8148
rect 39200 8064 40000 8092
rect 24882 7980 24892 8036
rect 24948 7980 36428 8036
rect 36484 7980 37212 8036
rect 37268 7980 37278 8036
rect 10526 7812 10536 7868
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10800 7812 10810 7868
rect 19850 7812 19860 7868
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 20124 7812 20134 7868
rect 29174 7812 29184 7868
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29448 7812 29458 7868
rect 38498 7812 38508 7868
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38772 7812 38782 7868
rect 39200 7476 40000 7504
rect 37538 7420 37548 7476
rect 37604 7420 40000 7476
rect 39200 7392 40000 7420
rect 28578 7308 28588 7364
rect 28644 7308 37212 7364
rect 37268 7308 37884 7364
rect 37940 7308 37950 7364
rect 5864 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6148 7084
rect 15188 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15472 7084
rect 24512 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24796 7084
rect 33836 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34120 7084
rect 39200 6804 40000 6832
rect 38210 6748 38220 6804
rect 38276 6748 40000 6804
rect 39200 6720 40000 6748
rect 26674 6524 26684 6580
rect 26740 6524 37548 6580
rect 37604 6524 37614 6580
rect 10526 6244 10536 6300
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10800 6244 10810 6300
rect 19850 6244 19860 6300
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 20124 6244 20134 6300
rect 29174 6244 29184 6300
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29448 6244 29458 6300
rect 38498 6244 38508 6300
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38772 6244 38782 6300
rect 38210 6188 38220 6244
rect 38276 6188 38286 6244
rect 38220 6132 38276 6188
rect 39200 6132 40000 6160
rect 38220 6076 40000 6132
rect 39200 6048 40000 6076
rect 29922 5740 29932 5796
rect 29988 5740 37660 5796
rect 37716 5740 37726 5796
rect 5864 5460 5874 5516
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 6138 5460 6148 5516
rect 15188 5460 15198 5516
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15462 5460 15472 5516
rect 24512 5460 24522 5516
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24786 5460 24796 5516
rect 33836 5460 33846 5516
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 34110 5460 34120 5516
rect 39200 5460 40000 5488
rect 38210 5404 38220 5460
rect 38276 5404 40000 5460
rect 39200 5376 40000 5404
rect 31266 5068 31276 5124
rect 31332 5068 37548 5124
rect 37604 5068 37996 5124
rect 38052 5068 38062 5124
rect 23538 4956 23548 5012
rect 23604 4956 27468 5012
rect 27524 4956 27534 5012
rect 38210 4844 38220 4900
rect 38276 4844 38948 4900
rect 38892 4788 38948 4844
rect 39200 4788 40000 4816
rect 38892 4732 40000 4788
rect 10526 4676 10536 4732
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10800 4676 10810 4732
rect 19850 4676 19860 4732
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 20124 4676 20134 4732
rect 29174 4676 29184 4732
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29448 4676 29458 4732
rect 38498 4676 38508 4732
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38772 4676 38782 4732
rect 39200 4704 40000 4732
rect 24994 4172 25004 4228
rect 25060 4172 37660 4228
rect 37716 4172 37726 4228
rect 39200 4116 40000 4144
rect 38210 4060 38220 4116
rect 38276 4060 40000 4116
rect 39200 4032 40000 4060
rect 5864 3892 5874 3948
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 6138 3892 6148 3948
rect 15188 3892 15198 3948
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15462 3892 15472 3948
rect 24512 3892 24522 3948
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24786 3892 24796 3948
rect 33836 3892 33846 3948
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 34110 3892 34120 3948
rect 24882 3612 24892 3668
rect 24948 3612 25676 3668
rect 25732 3612 26124 3668
rect 26180 3612 26190 3668
rect 24098 3500 24108 3556
rect 24164 3500 24780 3556
rect 24836 3500 24846 3556
rect 39200 3444 40000 3472
rect 24210 3388 24220 3444
rect 24276 3388 25228 3444
rect 25284 3388 25294 3444
rect 26114 3388 26124 3444
rect 26180 3388 27244 3444
rect 27300 3388 27310 3444
rect 31826 3388 31836 3444
rect 31892 3388 36428 3444
rect 36484 3388 37884 3444
rect 37940 3388 37950 3444
rect 38210 3388 38220 3444
rect 38276 3388 40000 3444
rect 39200 3360 40000 3388
rect 10526 3108 10536 3164
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10800 3108 10810 3164
rect 19850 3108 19860 3164
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 20124 3108 20134 3164
rect 29174 3108 29184 3164
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29448 3108 29458 3164
rect 38498 3108 38508 3164
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38772 3108 38782 3164
rect 39200 2772 40000 2800
rect 37538 2716 37548 2772
rect 37604 2716 40000 2772
rect 39200 2688 40000 2716
<< via3 >>
rect 5874 36820 5930 36876
rect 5978 36820 6034 36876
rect 6082 36820 6138 36876
rect 15198 36820 15254 36876
rect 15302 36820 15358 36876
rect 15406 36820 15462 36876
rect 24522 36820 24578 36876
rect 24626 36820 24682 36876
rect 24730 36820 24786 36876
rect 33846 36820 33902 36876
rect 33950 36820 34006 36876
rect 34054 36820 34110 36876
rect 10536 36036 10592 36092
rect 10640 36036 10696 36092
rect 10744 36036 10800 36092
rect 19860 36036 19916 36092
rect 19964 36036 20020 36092
rect 20068 36036 20124 36092
rect 29184 36036 29240 36092
rect 29288 36036 29344 36092
rect 29392 36036 29448 36092
rect 38508 36036 38564 36092
rect 38612 36036 38668 36092
rect 38716 36036 38772 36092
rect 5874 35252 5930 35308
rect 5978 35252 6034 35308
rect 6082 35252 6138 35308
rect 15198 35252 15254 35308
rect 15302 35252 15358 35308
rect 15406 35252 15462 35308
rect 24522 35252 24578 35308
rect 24626 35252 24682 35308
rect 24730 35252 24786 35308
rect 33846 35252 33902 35308
rect 33950 35252 34006 35308
rect 34054 35252 34110 35308
rect 10536 34468 10592 34524
rect 10640 34468 10696 34524
rect 10744 34468 10800 34524
rect 19860 34468 19916 34524
rect 19964 34468 20020 34524
rect 20068 34468 20124 34524
rect 29184 34468 29240 34524
rect 29288 34468 29344 34524
rect 29392 34468 29448 34524
rect 38508 34468 38564 34524
rect 38612 34468 38668 34524
rect 38716 34468 38772 34524
rect 5874 33684 5930 33740
rect 5978 33684 6034 33740
rect 6082 33684 6138 33740
rect 15198 33684 15254 33740
rect 15302 33684 15358 33740
rect 15406 33684 15462 33740
rect 24522 33684 24578 33740
rect 24626 33684 24682 33740
rect 24730 33684 24786 33740
rect 33846 33684 33902 33740
rect 33950 33684 34006 33740
rect 34054 33684 34110 33740
rect 10536 32900 10592 32956
rect 10640 32900 10696 32956
rect 10744 32900 10800 32956
rect 19860 32900 19916 32956
rect 19964 32900 20020 32956
rect 20068 32900 20124 32956
rect 29184 32900 29240 32956
rect 29288 32900 29344 32956
rect 29392 32900 29448 32956
rect 38508 32900 38564 32956
rect 38612 32900 38668 32956
rect 38716 32900 38772 32956
rect 5874 32116 5930 32172
rect 5978 32116 6034 32172
rect 6082 32116 6138 32172
rect 15198 32116 15254 32172
rect 15302 32116 15358 32172
rect 15406 32116 15462 32172
rect 24522 32116 24578 32172
rect 24626 32116 24682 32172
rect 24730 32116 24786 32172
rect 33846 32116 33902 32172
rect 33950 32116 34006 32172
rect 34054 32116 34110 32172
rect 10536 31332 10592 31388
rect 10640 31332 10696 31388
rect 10744 31332 10800 31388
rect 19860 31332 19916 31388
rect 19964 31332 20020 31388
rect 20068 31332 20124 31388
rect 29184 31332 29240 31388
rect 29288 31332 29344 31388
rect 29392 31332 29448 31388
rect 38508 31332 38564 31388
rect 38612 31332 38668 31388
rect 38716 31332 38772 31388
rect 5874 30548 5930 30604
rect 5978 30548 6034 30604
rect 6082 30548 6138 30604
rect 15198 30548 15254 30604
rect 15302 30548 15358 30604
rect 15406 30548 15462 30604
rect 24522 30548 24578 30604
rect 24626 30548 24682 30604
rect 24730 30548 24786 30604
rect 33846 30548 33902 30604
rect 33950 30548 34006 30604
rect 34054 30548 34110 30604
rect 10536 29764 10592 29820
rect 10640 29764 10696 29820
rect 10744 29764 10800 29820
rect 19860 29764 19916 29820
rect 19964 29764 20020 29820
rect 20068 29764 20124 29820
rect 29184 29764 29240 29820
rect 29288 29764 29344 29820
rect 29392 29764 29448 29820
rect 38508 29764 38564 29820
rect 38612 29764 38668 29820
rect 38716 29764 38772 29820
rect 5874 28980 5930 29036
rect 5978 28980 6034 29036
rect 6082 28980 6138 29036
rect 15198 28980 15254 29036
rect 15302 28980 15358 29036
rect 15406 28980 15462 29036
rect 24522 28980 24578 29036
rect 24626 28980 24682 29036
rect 24730 28980 24786 29036
rect 33846 28980 33902 29036
rect 33950 28980 34006 29036
rect 34054 28980 34110 29036
rect 10536 28196 10592 28252
rect 10640 28196 10696 28252
rect 10744 28196 10800 28252
rect 19860 28196 19916 28252
rect 19964 28196 20020 28252
rect 20068 28196 20124 28252
rect 29184 28196 29240 28252
rect 29288 28196 29344 28252
rect 29392 28196 29448 28252
rect 38508 28196 38564 28252
rect 38612 28196 38668 28252
rect 38716 28196 38772 28252
rect 5874 27412 5930 27468
rect 5978 27412 6034 27468
rect 6082 27412 6138 27468
rect 15198 27412 15254 27468
rect 15302 27412 15358 27468
rect 15406 27412 15462 27468
rect 24522 27412 24578 27468
rect 24626 27412 24682 27468
rect 24730 27412 24786 27468
rect 33846 27412 33902 27468
rect 33950 27412 34006 27468
rect 34054 27412 34110 27468
rect 10536 26628 10592 26684
rect 10640 26628 10696 26684
rect 10744 26628 10800 26684
rect 19860 26628 19916 26684
rect 19964 26628 20020 26684
rect 20068 26628 20124 26684
rect 29184 26628 29240 26684
rect 29288 26628 29344 26684
rect 29392 26628 29448 26684
rect 38508 26628 38564 26684
rect 38612 26628 38668 26684
rect 38716 26628 38772 26684
rect 5874 25844 5930 25900
rect 5978 25844 6034 25900
rect 6082 25844 6138 25900
rect 15198 25844 15254 25900
rect 15302 25844 15358 25900
rect 15406 25844 15462 25900
rect 24522 25844 24578 25900
rect 24626 25844 24682 25900
rect 24730 25844 24786 25900
rect 33846 25844 33902 25900
rect 33950 25844 34006 25900
rect 34054 25844 34110 25900
rect 10536 25060 10592 25116
rect 10640 25060 10696 25116
rect 10744 25060 10800 25116
rect 19860 25060 19916 25116
rect 19964 25060 20020 25116
rect 20068 25060 20124 25116
rect 29184 25060 29240 25116
rect 29288 25060 29344 25116
rect 29392 25060 29448 25116
rect 38508 25060 38564 25116
rect 38612 25060 38668 25116
rect 38716 25060 38772 25116
rect 5874 24276 5930 24332
rect 5978 24276 6034 24332
rect 6082 24276 6138 24332
rect 15198 24276 15254 24332
rect 15302 24276 15358 24332
rect 15406 24276 15462 24332
rect 24522 24276 24578 24332
rect 24626 24276 24682 24332
rect 24730 24276 24786 24332
rect 33846 24276 33902 24332
rect 33950 24276 34006 24332
rect 34054 24276 34110 24332
rect 10536 23492 10592 23548
rect 10640 23492 10696 23548
rect 10744 23492 10800 23548
rect 19860 23492 19916 23548
rect 19964 23492 20020 23548
rect 20068 23492 20124 23548
rect 29184 23492 29240 23548
rect 29288 23492 29344 23548
rect 29392 23492 29448 23548
rect 38508 23492 38564 23548
rect 38612 23492 38668 23548
rect 38716 23492 38772 23548
rect 5874 22708 5930 22764
rect 5978 22708 6034 22764
rect 6082 22708 6138 22764
rect 15198 22708 15254 22764
rect 15302 22708 15358 22764
rect 15406 22708 15462 22764
rect 24522 22708 24578 22764
rect 24626 22708 24682 22764
rect 24730 22708 24786 22764
rect 33846 22708 33902 22764
rect 33950 22708 34006 22764
rect 34054 22708 34110 22764
rect 10536 21924 10592 21980
rect 10640 21924 10696 21980
rect 10744 21924 10800 21980
rect 19860 21924 19916 21980
rect 19964 21924 20020 21980
rect 20068 21924 20124 21980
rect 29184 21924 29240 21980
rect 29288 21924 29344 21980
rect 29392 21924 29448 21980
rect 38508 21924 38564 21980
rect 38612 21924 38668 21980
rect 38716 21924 38772 21980
rect 5874 21140 5930 21196
rect 5978 21140 6034 21196
rect 6082 21140 6138 21196
rect 15198 21140 15254 21196
rect 15302 21140 15358 21196
rect 15406 21140 15462 21196
rect 24522 21140 24578 21196
rect 24626 21140 24682 21196
rect 24730 21140 24786 21196
rect 33846 21140 33902 21196
rect 33950 21140 34006 21196
rect 34054 21140 34110 21196
rect 10536 20356 10592 20412
rect 10640 20356 10696 20412
rect 10744 20356 10800 20412
rect 19860 20356 19916 20412
rect 19964 20356 20020 20412
rect 20068 20356 20124 20412
rect 29184 20356 29240 20412
rect 29288 20356 29344 20412
rect 29392 20356 29448 20412
rect 38508 20356 38564 20412
rect 38612 20356 38668 20412
rect 38716 20356 38772 20412
rect 5874 19572 5930 19628
rect 5978 19572 6034 19628
rect 6082 19572 6138 19628
rect 15198 19572 15254 19628
rect 15302 19572 15358 19628
rect 15406 19572 15462 19628
rect 24522 19572 24578 19628
rect 24626 19572 24682 19628
rect 24730 19572 24786 19628
rect 33846 19572 33902 19628
rect 33950 19572 34006 19628
rect 34054 19572 34110 19628
rect 10536 18788 10592 18844
rect 10640 18788 10696 18844
rect 10744 18788 10800 18844
rect 19860 18788 19916 18844
rect 19964 18788 20020 18844
rect 20068 18788 20124 18844
rect 29184 18788 29240 18844
rect 29288 18788 29344 18844
rect 29392 18788 29448 18844
rect 38508 18788 38564 18844
rect 38612 18788 38668 18844
rect 38716 18788 38772 18844
rect 5874 18004 5930 18060
rect 5978 18004 6034 18060
rect 6082 18004 6138 18060
rect 15198 18004 15254 18060
rect 15302 18004 15358 18060
rect 15406 18004 15462 18060
rect 24522 18004 24578 18060
rect 24626 18004 24682 18060
rect 24730 18004 24786 18060
rect 33846 18004 33902 18060
rect 33950 18004 34006 18060
rect 34054 18004 34110 18060
rect 10536 17220 10592 17276
rect 10640 17220 10696 17276
rect 10744 17220 10800 17276
rect 19860 17220 19916 17276
rect 19964 17220 20020 17276
rect 20068 17220 20124 17276
rect 29184 17220 29240 17276
rect 29288 17220 29344 17276
rect 29392 17220 29448 17276
rect 38508 17220 38564 17276
rect 38612 17220 38668 17276
rect 38716 17220 38772 17276
rect 5874 16436 5930 16492
rect 5978 16436 6034 16492
rect 6082 16436 6138 16492
rect 15198 16436 15254 16492
rect 15302 16436 15358 16492
rect 15406 16436 15462 16492
rect 24522 16436 24578 16492
rect 24626 16436 24682 16492
rect 24730 16436 24786 16492
rect 33846 16436 33902 16492
rect 33950 16436 34006 16492
rect 34054 16436 34110 16492
rect 10536 15652 10592 15708
rect 10640 15652 10696 15708
rect 10744 15652 10800 15708
rect 19860 15652 19916 15708
rect 19964 15652 20020 15708
rect 20068 15652 20124 15708
rect 29184 15652 29240 15708
rect 29288 15652 29344 15708
rect 29392 15652 29448 15708
rect 38508 15652 38564 15708
rect 38612 15652 38668 15708
rect 38716 15652 38772 15708
rect 5874 14868 5930 14924
rect 5978 14868 6034 14924
rect 6082 14868 6138 14924
rect 15198 14868 15254 14924
rect 15302 14868 15358 14924
rect 15406 14868 15462 14924
rect 24522 14868 24578 14924
rect 24626 14868 24682 14924
rect 24730 14868 24786 14924
rect 33846 14868 33902 14924
rect 33950 14868 34006 14924
rect 34054 14868 34110 14924
rect 10536 14084 10592 14140
rect 10640 14084 10696 14140
rect 10744 14084 10800 14140
rect 19860 14084 19916 14140
rect 19964 14084 20020 14140
rect 20068 14084 20124 14140
rect 29184 14084 29240 14140
rect 29288 14084 29344 14140
rect 29392 14084 29448 14140
rect 38508 14084 38564 14140
rect 38612 14084 38668 14140
rect 38716 14084 38772 14140
rect 5874 13300 5930 13356
rect 5978 13300 6034 13356
rect 6082 13300 6138 13356
rect 15198 13300 15254 13356
rect 15302 13300 15358 13356
rect 15406 13300 15462 13356
rect 24522 13300 24578 13356
rect 24626 13300 24682 13356
rect 24730 13300 24786 13356
rect 33846 13300 33902 13356
rect 33950 13300 34006 13356
rect 34054 13300 34110 13356
rect 10536 12516 10592 12572
rect 10640 12516 10696 12572
rect 10744 12516 10800 12572
rect 19860 12516 19916 12572
rect 19964 12516 20020 12572
rect 20068 12516 20124 12572
rect 29184 12516 29240 12572
rect 29288 12516 29344 12572
rect 29392 12516 29448 12572
rect 38508 12516 38564 12572
rect 38612 12516 38668 12572
rect 38716 12516 38772 12572
rect 5874 11732 5930 11788
rect 5978 11732 6034 11788
rect 6082 11732 6138 11788
rect 15198 11732 15254 11788
rect 15302 11732 15358 11788
rect 15406 11732 15462 11788
rect 24522 11732 24578 11788
rect 24626 11732 24682 11788
rect 24730 11732 24786 11788
rect 33846 11732 33902 11788
rect 33950 11732 34006 11788
rect 34054 11732 34110 11788
rect 10536 10948 10592 11004
rect 10640 10948 10696 11004
rect 10744 10948 10800 11004
rect 19860 10948 19916 11004
rect 19964 10948 20020 11004
rect 20068 10948 20124 11004
rect 29184 10948 29240 11004
rect 29288 10948 29344 11004
rect 29392 10948 29448 11004
rect 38508 10948 38564 11004
rect 38612 10948 38668 11004
rect 38716 10948 38772 11004
rect 5874 10164 5930 10220
rect 5978 10164 6034 10220
rect 6082 10164 6138 10220
rect 15198 10164 15254 10220
rect 15302 10164 15358 10220
rect 15406 10164 15462 10220
rect 24522 10164 24578 10220
rect 24626 10164 24682 10220
rect 24730 10164 24786 10220
rect 33846 10164 33902 10220
rect 33950 10164 34006 10220
rect 34054 10164 34110 10220
rect 10536 9380 10592 9436
rect 10640 9380 10696 9436
rect 10744 9380 10800 9436
rect 19860 9380 19916 9436
rect 19964 9380 20020 9436
rect 20068 9380 20124 9436
rect 29184 9380 29240 9436
rect 29288 9380 29344 9436
rect 29392 9380 29448 9436
rect 38508 9380 38564 9436
rect 38612 9380 38668 9436
rect 38716 9380 38772 9436
rect 5874 8596 5930 8652
rect 5978 8596 6034 8652
rect 6082 8596 6138 8652
rect 15198 8596 15254 8652
rect 15302 8596 15358 8652
rect 15406 8596 15462 8652
rect 24522 8596 24578 8652
rect 24626 8596 24682 8652
rect 24730 8596 24786 8652
rect 33846 8596 33902 8652
rect 33950 8596 34006 8652
rect 34054 8596 34110 8652
rect 10536 7812 10592 7868
rect 10640 7812 10696 7868
rect 10744 7812 10800 7868
rect 19860 7812 19916 7868
rect 19964 7812 20020 7868
rect 20068 7812 20124 7868
rect 29184 7812 29240 7868
rect 29288 7812 29344 7868
rect 29392 7812 29448 7868
rect 38508 7812 38564 7868
rect 38612 7812 38668 7868
rect 38716 7812 38772 7868
rect 5874 7028 5930 7084
rect 5978 7028 6034 7084
rect 6082 7028 6138 7084
rect 15198 7028 15254 7084
rect 15302 7028 15358 7084
rect 15406 7028 15462 7084
rect 24522 7028 24578 7084
rect 24626 7028 24682 7084
rect 24730 7028 24786 7084
rect 33846 7028 33902 7084
rect 33950 7028 34006 7084
rect 34054 7028 34110 7084
rect 10536 6244 10592 6300
rect 10640 6244 10696 6300
rect 10744 6244 10800 6300
rect 19860 6244 19916 6300
rect 19964 6244 20020 6300
rect 20068 6244 20124 6300
rect 29184 6244 29240 6300
rect 29288 6244 29344 6300
rect 29392 6244 29448 6300
rect 38508 6244 38564 6300
rect 38612 6244 38668 6300
rect 38716 6244 38772 6300
rect 5874 5460 5930 5516
rect 5978 5460 6034 5516
rect 6082 5460 6138 5516
rect 15198 5460 15254 5516
rect 15302 5460 15358 5516
rect 15406 5460 15462 5516
rect 24522 5460 24578 5516
rect 24626 5460 24682 5516
rect 24730 5460 24786 5516
rect 33846 5460 33902 5516
rect 33950 5460 34006 5516
rect 34054 5460 34110 5516
rect 10536 4676 10592 4732
rect 10640 4676 10696 4732
rect 10744 4676 10800 4732
rect 19860 4676 19916 4732
rect 19964 4676 20020 4732
rect 20068 4676 20124 4732
rect 29184 4676 29240 4732
rect 29288 4676 29344 4732
rect 29392 4676 29448 4732
rect 38508 4676 38564 4732
rect 38612 4676 38668 4732
rect 38716 4676 38772 4732
rect 5874 3892 5930 3948
rect 5978 3892 6034 3948
rect 6082 3892 6138 3948
rect 15198 3892 15254 3948
rect 15302 3892 15358 3948
rect 15406 3892 15462 3948
rect 24522 3892 24578 3948
rect 24626 3892 24682 3948
rect 24730 3892 24786 3948
rect 33846 3892 33902 3948
rect 33950 3892 34006 3948
rect 34054 3892 34110 3948
rect 10536 3108 10592 3164
rect 10640 3108 10696 3164
rect 10744 3108 10800 3164
rect 19860 3108 19916 3164
rect 19964 3108 20020 3164
rect 20068 3108 20124 3164
rect 29184 3108 29240 3164
rect 29288 3108 29344 3164
rect 29392 3108 29448 3164
rect 38508 3108 38564 3164
rect 38612 3108 38668 3164
rect 38716 3108 38772 3164
<< metal4 >>
rect 5846 36876 6166 36908
rect 5846 36820 5874 36876
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 6138 36820 6166 36876
rect 5846 35308 6166 36820
rect 5846 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6166 35308
rect 5846 33740 6166 35252
rect 5846 33684 5874 33740
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 6138 33684 6166 33740
rect 5846 32172 6166 33684
rect 5846 32116 5874 32172
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 6138 32116 6166 32172
rect 5846 30604 6166 32116
rect 5846 30548 5874 30604
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 6138 30548 6166 30604
rect 5846 29036 6166 30548
rect 5846 28980 5874 29036
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 6138 28980 6166 29036
rect 5846 27468 6166 28980
rect 5846 27412 5874 27468
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 6138 27412 6166 27468
rect 5846 25900 6166 27412
rect 5846 25844 5874 25900
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 6138 25844 6166 25900
rect 5846 24332 6166 25844
rect 5846 24276 5874 24332
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 6138 24276 6166 24332
rect 5846 22764 6166 24276
rect 5846 22708 5874 22764
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 6138 22708 6166 22764
rect 5846 21196 6166 22708
rect 5846 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6166 21196
rect 5846 19628 6166 21140
rect 5846 19572 5874 19628
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 6138 19572 6166 19628
rect 5846 18060 6166 19572
rect 5846 18004 5874 18060
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 6138 18004 6166 18060
rect 5846 16492 6166 18004
rect 5846 16436 5874 16492
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 6138 16436 6166 16492
rect 5846 14924 6166 16436
rect 5846 14868 5874 14924
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 6138 14868 6166 14924
rect 5846 13356 6166 14868
rect 5846 13300 5874 13356
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 6138 13300 6166 13356
rect 5846 11788 6166 13300
rect 5846 11732 5874 11788
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 6138 11732 6166 11788
rect 5846 10220 6166 11732
rect 5846 10164 5874 10220
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 6138 10164 6166 10220
rect 5846 8652 6166 10164
rect 5846 8596 5874 8652
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 6138 8596 6166 8652
rect 5846 7084 6166 8596
rect 5846 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6166 7084
rect 5846 5516 6166 7028
rect 5846 5460 5874 5516
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 6138 5460 6166 5516
rect 5846 3948 6166 5460
rect 5846 3892 5874 3948
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 6138 3892 6166 3948
rect 5846 3076 6166 3892
rect 10508 36092 10828 36908
rect 10508 36036 10536 36092
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10800 36036 10828 36092
rect 10508 34524 10828 36036
rect 10508 34468 10536 34524
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10800 34468 10828 34524
rect 10508 32956 10828 34468
rect 10508 32900 10536 32956
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10800 32900 10828 32956
rect 10508 31388 10828 32900
rect 10508 31332 10536 31388
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10800 31332 10828 31388
rect 10508 29820 10828 31332
rect 10508 29764 10536 29820
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10800 29764 10828 29820
rect 10508 28252 10828 29764
rect 10508 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10828 28252
rect 10508 26684 10828 28196
rect 10508 26628 10536 26684
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10800 26628 10828 26684
rect 10508 25116 10828 26628
rect 10508 25060 10536 25116
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10800 25060 10828 25116
rect 10508 23548 10828 25060
rect 10508 23492 10536 23548
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10800 23492 10828 23548
rect 10508 21980 10828 23492
rect 10508 21924 10536 21980
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10800 21924 10828 21980
rect 10508 20412 10828 21924
rect 10508 20356 10536 20412
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10800 20356 10828 20412
rect 10508 18844 10828 20356
rect 10508 18788 10536 18844
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10800 18788 10828 18844
rect 10508 17276 10828 18788
rect 10508 17220 10536 17276
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10800 17220 10828 17276
rect 10508 15708 10828 17220
rect 10508 15652 10536 15708
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10800 15652 10828 15708
rect 10508 14140 10828 15652
rect 10508 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10828 14140
rect 10508 12572 10828 14084
rect 10508 12516 10536 12572
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10800 12516 10828 12572
rect 10508 11004 10828 12516
rect 10508 10948 10536 11004
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10800 10948 10828 11004
rect 10508 9436 10828 10948
rect 10508 9380 10536 9436
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10800 9380 10828 9436
rect 10508 7868 10828 9380
rect 10508 7812 10536 7868
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10800 7812 10828 7868
rect 10508 6300 10828 7812
rect 10508 6244 10536 6300
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10800 6244 10828 6300
rect 10508 4732 10828 6244
rect 10508 4676 10536 4732
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10800 4676 10828 4732
rect 10508 3164 10828 4676
rect 10508 3108 10536 3164
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10800 3108 10828 3164
rect 10508 3076 10828 3108
rect 15170 36876 15490 36908
rect 15170 36820 15198 36876
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15462 36820 15490 36876
rect 15170 35308 15490 36820
rect 15170 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15490 35308
rect 15170 33740 15490 35252
rect 15170 33684 15198 33740
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15462 33684 15490 33740
rect 15170 32172 15490 33684
rect 15170 32116 15198 32172
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15462 32116 15490 32172
rect 15170 30604 15490 32116
rect 15170 30548 15198 30604
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15462 30548 15490 30604
rect 15170 29036 15490 30548
rect 15170 28980 15198 29036
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15462 28980 15490 29036
rect 15170 27468 15490 28980
rect 15170 27412 15198 27468
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15462 27412 15490 27468
rect 15170 25900 15490 27412
rect 15170 25844 15198 25900
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15462 25844 15490 25900
rect 15170 24332 15490 25844
rect 15170 24276 15198 24332
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15462 24276 15490 24332
rect 15170 22764 15490 24276
rect 15170 22708 15198 22764
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15462 22708 15490 22764
rect 15170 21196 15490 22708
rect 15170 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15490 21196
rect 15170 19628 15490 21140
rect 15170 19572 15198 19628
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15462 19572 15490 19628
rect 15170 18060 15490 19572
rect 15170 18004 15198 18060
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15462 18004 15490 18060
rect 15170 16492 15490 18004
rect 15170 16436 15198 16492
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15462 16436 15490 16492
rect 15170 14924 15490 16436
rect 15170 14868 15198 14924
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15462 14868 15490 14924
rect 15170 13356 15490 14868
rect 15170 13300 15198 13356
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15462 13300 15490 13356
rect 15170 11788 15490 13300
rect 15170 11732 15198 11788
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15462 11732 15490 11788
rect 15170 10220 15490 11732
rect 15170 10164 15198 10220
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15462 10164 15490 10220
rect 15170 8652 15490 10164
rect 15170 8596 15198 8652
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15462 8596 15490 8652
rect 15170 7084 15490 8596
rect 15170 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15490 7084
rect 15170 5516 15490 7028
rect 15170 5460 15198 5516
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15462 5460 15490 5516
rect 15170 3948 15490 5460
rect 15170 3892 15198 3948
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15462 3892 15490 3948
rect 15170 3076 15490 3892
rect 19832 36092 20152 36908
rect 19832 36036 19860 36092
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 20124 36036 20152 36092
rect 19832 34524 20152 36036
rect 19832 34468 19860 34524
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 20124 34468 20152 34524
rect 19832 32956 20152 34468
rect 19832 32900 19860 32956
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 20124 32900 20152 32956
rect 19832 31388 20152 32900
rect 19832 31332 19860 31388
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 20124 31332 20152 31388
rect 19832 29820 20152 31332
rect 19832 29764 19860 29820
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 20124 29764 20152 29820
rect 19832 28252 20152 29764
rect 19832 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20152 28252
rect 19832 26684 20152 28196
rect 19832 26628 19860 26684
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 20124 26628 20152 26684
rect 19832 25116 20152 26628
rect 19832 25060 19860 25116
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 20124 25060 20152 25116
rect 19832 23548 20152 25060
rect 19832 23492 19860 23548
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 20124 23492 20152 23548
rect 19832 21980 20152 23492
rect 19832 21924 19860 21980
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 20124 21924 20152 21980
rect 19832 20412 20152 21924
rect 19832 20356 19860 20412
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 20124 20356 20152 20412
rect 19832 18844 20152 20356
rect 19832 18788 19860 18844
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 20124 18788 20152 18844
rect 19832 17276 20152 18788
rect 19832 17220 19860 17276
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 20124 17220 20152 17276
rect 19832 15708 20152 17220
rect 19832 15652 19860 15708
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 20124 15652 20152 15708
rect 19832 14140 20152 15652
rect 19832 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20152 14140
rect 19832 12572 20152 14084
rect 19832 12516 19860 12572
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 20124 12516 20152 12572
rect 19832 11004 20152 12516
rect 19832 10948 19860 11004
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 20124 10948 20152 11004
rect 19832 9436 20152 10948
rect 19832 9380 19860 9436
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 20124 9380 20152 9436
rect 19832 7868 20152 9380
rect 19832 7812 19860 7868
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 20124 7812 20152 7868
rect 19832 6300 20152 7812
rect 19832 6244 19860 6300
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 20124 6244 20152 6300
rect 19832 4732 20152 6244
rect 19832 4676 19860 4732
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 20124 4676 20152 4732
rect 19832 3164 20152 4676
rect 19832 3108 19860 3164
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 20124 3108 20152 3164
rect 19832 3076 20152 3108
rect 24494 36876 24814 36908
rect 24494 36820 24522 36876
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24786 36820 24814 36876
rect 24494 35308 24814 36820
rect 24494 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24814 35308
rect 24494 33740 24814 35252
rect 24494 33684 24522 33740
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24786 33684 24814 33740
rect 24494 32172 24814 33684
rect 24494 32116 24522 32172
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24786 32116 24814 32172
rect 24494 30604 24814 32116
rect 24494 30548 24522 30604
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24786 30548 24814 30604
rect 24494 29036 24814 30548
rect 24494 28980 24522 29036
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24786 28980 24814 29036
rect 24494 27468 24814 28980
rect 24494 27412 24522 27468
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24786 27412 24814 27468
rect 24494 25900 24814 27412
rect 24494 25844 24522 25900
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24786 25844 24814 25900
rect 24494 24332 24814 25844
rect 24494 24276 24522 24332
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24786 24276 24814 24332
rect 24494 22764 24814 24276
rect 24494 22708 24522 22764
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24786 22708 24814 22764
rect 24494 21196 24814 22708
rect 24494 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24814 21196
rect 24494 19628 24814 21140
rect 24494 19572 24522 19628
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24786 19572 24814 19628
rect 24494 18060 24814 19572
rect 24494 18004 24522 18060
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24786 18004 24814 18060
rect 24494 16492 24814 18004
rect 24494 16436 24522 16492
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24786 16436 24814 16492
rect 24494 14924 24814 16436
rect 24494 14868 24522 14924
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24786 14868 24814 14924
rect 24494 13356 24814 14868
rect 24494 13300 24522 13356
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24786 13300 24814 13356
rect 24494 11788 24814 13300
rect 24494 11732 24522 11788
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24786 11732 24814 11788
rect 24494 10220 24814 11732
rect 24494 10164 24522 10220
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24786 10164 24814 10220
rect 24494 8652 24814 10164
rect 24494 8596 24522 8652
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24786 8596 24814 8652
rect 24494 7084 24814 8596
rect 24494 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24814 7084
rect 24494 5516 24814 7028
rect 24494 5460 24522 5516
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24786 5460 24814 5516
rect 24494 3948 24814 5460
rect 24494 3892 24522 3948
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24786 3892 24814 3948
rect 24494 3076 24814 3892
rect 29156 36092 29476 36908
rect 29156 36036 29184 36092
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29448 36036 29476 36092
rect 29156 34524 29476 36036
rect 29156 34468 29184 34524
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29448 34468 29476 34524
rect 29156 32956 29476 34468
rect 29156 32900 29184 32956
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29448 32900 29476 32956
rect 29156 31388 29476 32900
rect 29156 31332 29184 31388
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29448 31332 29476 31388
rect 29156 29820 29476 31332
rect 29156 29764 29184 29820
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29448 29764 29476 29820
rect 29156 28252 29476 29764
rect 29156 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29476 28252
rect 29156 26684 29476 28196
rect 29156 26628 29184 26684
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29448 26628 29476 26684
rect 29156 25116 29476 26628
rect 29156 25060 29184 25116
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29448 25060 29476 25116
rect 29156 23548 29476 25060
rect 29156 23492 29184 23548
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29448 23492 29476 23548
rect 29156 21980 29476 23492
rect 29156 21924 29184 21980
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29448 21924 29476 21980
rect 29156 20412 29476 21924
rect 29156 20356 29184 20412
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29448 20356 29476 20412
rect 29156 18844 29476 20356
rect 29156 18788 29184 18844
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29448 18788 29476 18844
rect 29156 17276 29476 18788
rect 29156 17220 29184 17276
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29448 17220 29476 17276
rect 29156 15708 29476 17220
rect 29156 15652 29184 15708
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29448 15652 29476 15708
rect 29156 14140 29476 15652
rect 29156 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29476 14140
rect 29156 12572 29476 14084
rect 29156 12516 29184 12572
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29448 12516 29476 12572
rect 29156 11004 29476 12516
rect 29156 10948 29184 11004
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29448 10948 29476 11004
rect 29156 9436 29476 10948
rect 29156 9380 29184 9436
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29448 9380 29476 9436
rect 29156 7868 29476 9380
rect 29156 7812 29184 7868
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29448 7812 29476 7868
rect 29156 6300 29476 7812
rect 29156 6244 29184 6300
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29448 6244 29476 6300
rect 29156 4732 29476 6244
rect 29156 4676 29184 4732
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29448 4676 29476 4732
rect 29156 3164 29476 4676
rect 29156 3108 29184 3164
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29448 3108 29476 3164
rect 29156 3076 29476 3108
rect 33818 36876 34138 36908
rect 33818 36820 33846 36876
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 34110 36820 34138 36876
rect 33818 35308 34138 36820
rect 33818 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34138 35308
rect 33818 33740 34138 35252
rect 33818 33684 33846 33740
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 34110 33684 34138 33740
rect 33818 32172 34138 33684
rect 33818 32116 33846 32172
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 34110 32116 34138 32172
rect 33818 30604 34138 32116
rect 33818 30548 33846 30604
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 34110 30548 34138 30604
rect 33818 29036 34138 30548
rect 33818 28980 33846 29036
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 34110 28980 34138 29036
rect 33818 27468 34138 28980
rect 33818 27412 33846 27468
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 34110 27412 34138 27468
rect 33818 25900 34138 27412
rect 33818 25844 33846 25900
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 34110 25844 34138 25900
rect 33818 24332 34138 25844
rect 33818 24276 33846 24332
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 34110 24276 34138 24332
rect 33818 22764 34138 24276
rect 33818 22708 33846 22764
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 34110 22708 34138 22764
rect 33818 21196 34138 22708
rect 33818 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34138 21196
rect 33818 19628 34138 21140
rect 33818 19572 33846 19628
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 34110 19572 34138 19628
rect 33818 18060 34138 19572
rect 33818 18004 33846 18060
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 34110 18004 34138 18060
rect 33818 16492 34138 18004
rect 33818 16436 33846 16492
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 34110 16436 34138 16492
rect 33818 14924 34138 16436
rect 33818 14868 33846 14924
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 34110 14868 34138 14924
rect 33818 13356 34138 14868
rect 33818 13300 33846 13356
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 34110 13300 34138 13356
rect 33818 11788 34138 13300
rect 33818 11732 33846 11788
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 34110 11732 34138 11788
rect 33818 10220 34138 11732
rect 33818 10164 33846 10220
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 34110 10164 34138 10220
rect 33818 8652 34138 10164
rect 33818 8596 33846 8652
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 34110 8596 34138 8652
rect 33818 7084 34138 8596
rect 33818 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34138 7084
rect 33818 5516 34138 7028
rect 33818 5460 33846 5516
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 34110 5460 34138 5516
rect 33818 3948 34138 5460
rect 33818 3892 33846 3948
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 34110 3892 34138 3948
rect 33818 3076 34138 3892
rect 38480 36092 38800 36908
rect 38480 36036 38508 36092
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38772 36036 38800 36092
rect 38480 34524 38800 36036
rect 38480 34468 38508 34524
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38772 34468 38800 34524
rect 38480 32956 38800 34468
rect 38480 32900 38508 32956
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38772 32900 38800 32956
rect 38480 31388 38800 32900
rect 38480 31332 38508 31388
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38772 31332 38800 31388
rect 38480 29820 38800 31332
rect 38480 29764 38508 29820
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38772 29764 38800 29820
rect 38480 28252 38800 29764
rect 38480 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38800 28252
rect 38480 26684 38800 28196
rect 38480 26628 38508 26684
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38772 26628 38800 26684
rect 38480 25116 38800 26628
rect 38480 25060 38508 25116
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38772 25060 38800 25116
rect 38480 23548 38800 25060
rect 38480 23492 38508 23548
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38772 23492 38800 23548
rect 38480 21980 38800 23492
rect 38480 21924 38508 21980
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38772 21924 38800 21980
rect 38480 20412 38800 21924
rect 38480 20356 38508 20412
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38772 20356 38800 20412
rect 38480 18844 38800 20356
rect 38480 18788 38508 18844
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38772 18788 38800 18844
rect 38480 17276 38800 18788
rect 38480 17220 38508 17276
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38772 17220 38800 17276
rect 38480 15708 38800 17220
rect 38480 15652 38508 15708
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38772 15652 38800 15708
rect 38480 14140 38800 15652
rect 38480 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38800 14140
rect 38480 12572 38800 14084
rect 38480 12516 38508 12572
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38772 12516 38800 12572
rect 38480 11004 38800 12516
rect 38480 10948 38508 11004
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38772 10948 38800 11004
rect 38480 9436 38800 10948
rect 38480 9380 38508 9436
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38772 9380 38800 9436
rect 38480 7868 38800 9380
rect 38480 7812 38508 7868
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38772 7812 38800 7868
rect 38480 6300 38800 7812
rect 38480 6244 38508 6300
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38772 6244 38800 6300
rect 38480 4732 38800 6244
rect 38480 4676 38508 4732
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38772 4676 38800 4732
rect 38480 3164 38800 4676
rect 38480 3108 38508 3164
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38772 3108 38800 3164
rect 38480 3076 38800 3108
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _126_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15344 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _127_
timestamp 1698431365
transform 1 0 15456 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _128_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18704 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18704 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _130_
timestamp 1698431365
transform -1 0 19824 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _131_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _132_
timestamp 1698431365
transform -1 0 20720 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _133_
timestamp 1698431365
transform 1 0 17248 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _134_
timestamp 1698431365
transform -1 0 18256 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _135_
timestamp 1698431365
transform 1 0 18256 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _136_
timestamp 1698431365
transform -1 0 20160 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _137_
timestamp 1698431365
transform -1 0 19040 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _138_
timestamp 1698431365
transform -1 0 18256 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _139_
timestamp 1698431365
transform -1 0 28672 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _140_
timestamp 1698431365
transform 1 0 27664 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _141_
timestamp 1698431365
transform 1 0 28112 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _142_
timestamp 1698431365
transform 1 0 27216 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _143_
timestamp 1698431365
transform 1 0 28112 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _144_
timestamp 1698431365
transform 1 0 28560 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _145_
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _146_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _147_
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _148_
timestamp 1698431365
transform 1 0 22288 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _149_
timestamp 1698431365
transform 1 0 22624 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _150_
timestamp 1698431365
transform 1 0 23072 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _151_
timestamp 1698431365
transform 1 0 23520 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _152_
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _153_
timestamp 1698431365
transform 1 0 24080 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _154_
timestamp 1698431365
transform 1 0 24976 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _155_
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _156_
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _157_
timestamp 1698431365
transform 1 0 28672 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _158_
timestamp 1698431365
transform 1 0 30576 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _159_
timestamp 1698431365
transform 1 0 31472 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _160_
timestamp 1698431365
transform 1 0 29680 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _161_
timestamp 1698431365
transform 1 0 30576 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _162_
timestamp 1698431365
transform 1 0 29680 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _163_
timestamp 1698431365
transform 1 0 30352 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _164_
timestamp 1698431365
transform 1 0 28784 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _165_
timestamp 1698431365
transform 1 0 29344 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _166_
timestamp 1698431365
transform -1 0 18704 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _167_
timestamp 1698431365
transform -1 0 13216 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _168_
timestamp 1698431365
transform -1 0 12432 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _169_
timestamp 1698431365
transform -1 0 12320 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _170_
timestamp 1698431365
transform -1 0 11648 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _171_
timestamp 1698431365
transform 1 0 11648 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _172_
timestamp 1698431365
transform -1 0 12880 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _173_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _174_
timestamp 1698431365
transform 1 0 19488 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _175_
timestamp 1698431365
transform 1 0 19936 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _176_
timestamp 1698431365
transform 1 0 18704 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _177_
timestamp 1698431365
transform 1 0 20608 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _178_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _179_
timestamp 1698431365
transform 1 0 22960 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _180_
timestamp 1698431365
transform 1 0 21616 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _181_
timestamp 1698431365
transform 1 0 22960 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _182_
timestamp 1698431365
transform 1 0 20832 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _183_
timestamp 1698431365
transform 1 0 22288 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _184_
timestamp 1698431365
transform 1 0 21616 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _185_
timestamp 1698431365
transform 1 0 23632 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _186_
timestamp 1698431365
transform 1 0 26880 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _187_
timestamp 1698431365
transform 1 0 26320 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _188_
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _189_
timestamp 1698431365
transform 1 0 29792 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _190_
timestamp 1698431365
transform 1 0 26992 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _191_
timestamp 1698431365
transform 1 0 27664 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _192_
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _193_
timestamp 1698431365
transform 1 0 30128 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _194_
timestamp 1698431365
transform 1 0 28672 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _195_
timestamp 1698431365
transform 1 0 30800 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _196_
timestamp 1698431365
transform -1 0 20944 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _197_
timestamp 1698431365
transform 1 0 19600 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _198_
timestamp 1698431365
transform 1 0 20608 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _199_
timestamp 1698431365
transform 1 0 21392 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _200_
timestamp 1698431365
transform -1 0 22288 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _201_
timestamp 1698431365
transform 1 0 20272 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _202_
timestamp 1698431365
transform -1 0 20608 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _203_
timestamp 1698431365
transform -1 0 20272 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _204_
timestamp 1698431365
transform 1 0 20720 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _205_
timestamp 1698431365
transform 1 0 21840 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _206_
timestamp 1698431365
transform 1 0 25872 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _207_
timestamp 1698431365
transform 1 0 26544 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _208_
timestamp 1698431365
transform 1 0 26992 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _209_
timestamp 1698431365
transform 1 0 28448 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _210_
timestamp 1698431365
transform 1 0 26992 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _211_
timestamp 1698431365
transform 1 0 27776 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _212_
timestamp 1698431365
transform -1 0 26992 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _213_
timestamp 1698431365
transform 1 0 26320 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _214_
timestamp 1698431365
transform 1 0 26992 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _215_
timestamp 1698431365
transform 1 0 28112 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _216_
timestamp 1698431365
transform -1 0 19376 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _217_
timestamp 1698431365
transform -1 0 16688 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _218_
timestamp 1698431365
transform 1 0 14896 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _219_
timestamp 1698431365
transform -1 0 15456 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _220_
timestamp 1698431365
transform 1 0 13776 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _221_
timestamp 1698431365
transform -1 0 15904 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _222_
timestamp 1698431365
transform 1 0 13776 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _223_
timestamp 1698431365
transform -1 0 15232 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _224_
timestamp 1698431365
transform 1 0 19488 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _225_
timestamp 1698431365
transform -1 0 23072 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _226_
timestamp 1698431365
transform 1 0 17584 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _227_
timestamp 1698431365
transform 1 0 19376 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _228_
timestamp 1698431365
transform 1 0 20272 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _229_
timestamp 1698431365
transform 1 0 21280 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _230_
timestamp 1698431365
transform 1 0 23072 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _231_
timestamp 1698431365
transform 1 0 21504 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _232_
timestamp 1698431365
transform 1 0 22736 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _233_
timestamp 1698431365
transform 1 0 21280 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _234_
timestamp 1698431365
transform 1 0 22624 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _235_
timestamp 1698431365
transform 1 0 21504 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _236_
timestamp 1698431365
transform 1 0 23408 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _237_
timestamp 1698431365
transform 1 0 23856 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _238_
timestamp 1698431365
transform 1 0 23184 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _239_
timestamp 1698431365
transform 1 0 25088 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _240_
timestamp 1698431365
transform 1 0 26208 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _241_
timestamp 1698431365
transform -1 0 24864 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _242_
timestamp 1698431365
transform 1 0 23968 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _243_
timestamp 1698431365
transform 1 0 24864 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _244_
timestamp 1698431365
transform 1 0 25648 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _245_
timestamp 1698431365
transform 1 0 25984 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _246_
timestamp 1698431365
transform 1 0 27104 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _247_
timestamp 1698431365
transform -1 0 24528 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _248_
timestamp 1698431365
transform 1 0 22960 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _249_
timestamp 1698431365
transform 1 0 22736 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _250_
timestamp 1698431365
transform 1 0 24528 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _251_
timestamp 1698431365
transform 1 0 22848 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _252_
timestamp 1698431365
transform 1 0 23968 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _253_
timestamp 1698431365
transform 1 0 23072 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _254_
timestamp 1698431365
transform 1 0 24528 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _255_
timestamp 1698431365
transform 1 0 22960 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _256_
timestamp 1698431365
transform 1 0 24192 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _257_
timestamp 1698431365
transform 1 0 25200 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _258_
timestamp 1698431365
transform 1 0 25872 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _259_
timestamp 1698431365
transform 1 0 30240 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _260_
timestamp 1698431365
transform 1 0 31360 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _261_
timestamp 1698431365
transform 1 0 29120 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _262_
timestamp 1698431365
transform 1 0 29904 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _263_
timestamp 1698431365
transform 1 0 29680 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _264_
timestamp 1698431365
transform 1 0 30800 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _265_
timestamp 1698431365
transform 1 0 28560 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _266_
timestamp 1698431365
transform 1 0 29456 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _267_
timestamp 1698431365
transform -1 0 15904 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _268_
timestamp 1698431365
transform -1 0 18704 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _269_
timestamp 1698431365
transform -1 0 14672 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _270_
timestamp 1698431365
transform -1 0 13104 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _271_
timestamp 1698431365
transform 1 0 13664 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _272_
timestamp 1698431365
transform -1 0 16128 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _273_
timestamp 1698431365
transform 1 0 13664 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _274_
timestamp 1698431365
transform -1 0 15456 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _275_
timestamp 1698431365
transform 1 0 15232 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _276_
timestamp 1698431365
transform 1 0 17472 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _277_
timestamp 1698431365
transform 1 0 18368 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _278_
timestamp 1698431365
transform -1 0 20048 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _279_
timestamp 1698431365
transform 1 0 19264 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _280_
timestamp 1698431365
transform -1 0 19040 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _281_
timestamp 1698431365
transform -1 0 18256 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _282_
timestamp 1698431365
transform 1 0 19040 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _283_
timestamp 1698431365
transform -1 0 20608 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _284_
timestamp 1698431365
transform 1 0 17248 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _285_
timestamp 1698431365
transform -1 0 18256 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _286_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _287_
timestamp 1698431365
transform 1 0 25984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _288_
timestamp 1698431365
transform 1 0 26208 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _289_
timestamp 1698431365
transform -1 0 25088 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _290_
timestamp 1698431365
transform 1 0 23520 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _291_
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _292_
timestamp 1698431365
transform 1 0 25536 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _293_
timestamp 1698431365
transform 1 0 25648 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _294_
timestamp 1698431365
transform 1 0 26544 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _295_
timestamp 1698431365
transform 1 0 18144 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _296_
timestamp 1698431365
transform -1 0 22064 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _297_
timestamp 1698431365
transform 1 0 20496 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _298_
timestamp 1698431365
transform 1 0 20048 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _299_
timestamp 1698431365
transform -1 0 22288 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _300_
timestamp 1698431365
transform -1 0 19936 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _301_
timestamp 1698431365
transform -1 0 19488 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _302_
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _303_
timestamp 1698431365
transform -1 0 24640 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _304_
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _305_
timestamp 1698431365
transform 1 0 27104 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _306_
timestamp 1698431365
transform 1 0 28000 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _307_
timestamp 1698431365
transform -1 0 28448 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _308_
timestamp 1698431365
transform 1 0 27552 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _309_
timestamp 1698431365
transform -1 0 26656 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _310_
timestamp 1698431365
transform 1 0 26096 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _311_
timestamp 1698431365
transform -1 0 27552 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _312_
timestamp 1698431365
transform 1 0 26992 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _313_
timestamp 1698431365
transform -1 0 17024 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _314_
timestamp 1698431365
transform 1 0 11536 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _315_
timestamp 1698431365
transform -1 0 12656 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _316_
timestamp 1698431365
transform -1 0 13216 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _317_
timestamp 1698431365
transform -1 0 13104 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _318_
timestamp 1698431365
transform -1 0 12320 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _319_
timestamp 1698431365
transform -1 0 11424 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _320_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17920 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _321_
timestamp 1698431365
transform -1 0 20608 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _322_
timestamp 1698431365
transform 1 0 17472 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _323_
timestamp 1698431365
transform 1 0 17920 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _324_
timestamp 1698431365
transform 1 0 19040 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _325__1
timestamp 1698431365
transform -1 0 20160 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _326_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18144 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _327_
timestamp 1698431365
transform -1 0 19824 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _328_
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _329_
timestamp 1698431365
transform -1 0 18480 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _330_
timestamp 1698431365
transform 1 0 16016 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _331_
timestamp 1698431365
transform -1 0 17808 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _332_
timestamp 1698431365
transform 1 0 15904 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _333_
timestamp 1698431365
transform -1 0 17472 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _334_
timestamp 1698431365
transform 1 0 16464 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _335_
timestamp 1698431365
transform -1 0 18032 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _336_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13776 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _337_
timestamp 1698431365
transform 1 0 14000 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__131__A1 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__A1
timestamp 1698431365
transform 1 0 16576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__A1
timestamp 1698431365
transform 1 0 19152 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__137__A1
timestamp 1698431365
transform 1 0 17024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__A1
timestamp 1698431365
transform 1 0 29680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__A1
timestamp 1698431365
transform 1 0 28896 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__A1
timestamp 1698431365
transform 1 0 30128 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__A1
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__151__A1
timestamp 1698431365
transform 1 0 24416 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__153__A1
timestamp 1698431365
transform 1 0 25872 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__A1
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__A1
timestamp 1698431365
transform 1 0 31472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__A1
timestamp 1698431365
transform 1 0 30576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__A1
timestamp 1698431365
transform 1 0 11200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__A1
timestamp 1698431365
transform 1 0 10752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__A1
timestamp 1698431365
transform 1 0 10752 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__A1
timestamp 1698431365
transform 1 0 22288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__A1
timestamp 1698431365
transform 1 0 21392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__A1
timestamp 1698431365
transform 1 0 22176 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__A1
timestamp 1698431365
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__A1
timestamp 1698431365
transform 1 0 30352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__A1
timestamp 1698431365
transform -1 0 28560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__A1
timestamp 1698431365
transform 1 0 30128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__A1
timestamp 1698431365
transform 1 0 21952 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__A1
timestamp 1698431365
transform -1 0 22736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__A1
timestamp 1698431365
transform -1 0 19488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__A1
timestamp 1698431365
transform 1 0 29232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__A1
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__A1
timestamp 1698431365
transform 1 0 28336 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__A1
timestamp 1698431365
transform 1 0 13552 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__A1
timestamp 1698431365
transform 1 0 13552 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__A1
timestamp 1698431365
transform 1 0 13552 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__A1
timestamp 1698431365
transform -1 0 22624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__A1
timestamp 1698431365
transform -1 0 21504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__A1
timestamp 1698431365
transform 1 0 22624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__A1
timestamp 1698431365
transform -1 0 21056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__A1
timestamp 1698431365
transform -1 0 25872 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__A1
timestamp 1698431365
transform -1 0 25536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__A1
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__A1
timestamp 1698431365
transform 1 0 22736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__A1
timestamp 1698431365
transform -1 0 24416 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__A1
timestamp 1698431365
transform 1 0 22848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__A1
timestamp 1698431365
transform -1 0 32480 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__A1
timestamp 1698431365
transform -1 0 31024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__A1
timestamp 1698431365
transform 1 0 31696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__A1
timestamp 1698431365
transform 1 0 12880 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__A1
timestamp 1698431365
transform 1 0 13440 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__273__A1
timestamp 1698431365
transform -1 0 13552 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__A1
timestamp 1698431365
transform 1 0 20272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__280__A1
timestamp 1698431365
transform 1 0 17024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__A1
timestamp 1698431365
transform -1 0 20608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__A1
timestamp 1698431365
transform -1 0 16800 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__A1
timestamp 1698431365
transform 1 0 27104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__A1
timestamp 1698431365
transform 1 0 25312 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__291__A1
timestamp 1698431365
transform 1 0 27104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__A1
timestamp 1698431365
transform 1 0 22288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__A1
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__A1
timestamp 1698431365
transform -1 0 19040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__A1
timestamp 1698431365
transform 1 0 28448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__A1
timestamp 1698431365
transform 1 0 28448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__A1
timestamp 1698431365
transform 1 0 26880 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__314__A1
timestamp 1698431365
transform 1 0 11312 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__A1
timestamp 1698431365
transform 1 0 11536 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__318__A1
timestamp 1698431365
transform 1 0 10528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__A1
timestamp 1698431365
transform 1 0 17696 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__A3
timestamp 1698431365
transform 1 0 15792 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__332__A3
timestamp 1698431365
transform 1 0 15008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__A1
timestamp 1698431365
transform 1 0 18256 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 25760 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 15904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 37072 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 37744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 37744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 37744 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 2464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 2464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 15232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 21616 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 16240 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 37744 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 37296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 37744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 25760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 26432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 3136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 2464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output44_I
timestamp 1698431365
transform -1 0 35616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output53_I
timestamp 1698431365
transform 1 0 37520 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output54_I
timestamp 1698431365
transform -1 0 37296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output55_I
timestamp 1698431365
transform 1 0 2464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output61_I
timestamp 1698431365
transform -1 0 37744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output62_I
timestamp 1698431365
transform -1 0 37744 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output64_I
timestamp 1698431365
transform -1 0 37744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output67_I
timestamp 1698431365
transform -1 0 37744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output69_I
timestamp 1698431365
transform 1 0 36400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output72_I
timestamp 1698431365
transform 1 0 36400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output74_I
timestamp 1698431365
transform 1 0 37520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output75_I
timestamp 1698431365
transform -1 0 37744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output82_I
timestamp 1698431365
transform 1 0 37520 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output84_I
timestamp 1698431365
transform 1 0 37072 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output85_I
timestamp 1698431365
transform -1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output86_I
timestamp 1698431365
transform -1 0 37744 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output87_I
timestamp 1698431365
transform 1 0 37520 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output103_I
timestamp 1698431365
transform 1 0 2464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698431365
transform -1 0 19040 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_104 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_120 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_199
timestamp 1698431365
transform 1 0 23632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698431365
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_312
timestamp 1698431365
transform 1 0 36288 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_315
timestamp 1698431365
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_104
timestamp 1698431365
transform 1 0 12992 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_120 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14784 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_128
timestamp 1698431365
transform 1 0 15680 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_132
timestamp 1698431365
transform 1 0 16128 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_218
timestamp 1698431365
transform 1 0 25760 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_224
timestamp 1698431365
transform 1 0 26432 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_256
timestamp 1698431365
transform 1 0 30016 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_272
timestamp 1698431365
transform 1 0 31808 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_314
timestamp 1698431365
transform 1 0 36512 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_322
timestamp 1698431365
transform 1 0 37408 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_321
timestamp 1698431365
transform 1 0 37296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_314
timestamp 1698431365
transform 1 0 36512 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_322
timestamp 1698431365
transform 1 0 37408 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_321
timestamp 1698431365
transform 1 0 37296 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_314
timestamp 1698431365
transform 1 0 36512 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_318
timestamp 1698431365
transform 1 0 36960 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_321
timestamp 1698431365
transform 1 0 37296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_314
timestamp 1698431365
transform 1 0 36512 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_322
timestamp 1698431365
transform 1 0 37408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_324
timestamp 1698431365
transform 1 0 37632 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_321
timestamp 1698431365
transform 1 0 37296 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_314
timestamp 1698431365
transform 1 0 36512 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_322
timestamp 1698431365
transform 1 0 37408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_324
timestamp 1698431365
transform 1 0 37632 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_314
timestamp 1698431365
transform 1 0 36512 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_322
timestamp 1698431365
transform 1 0 37408 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_8
timestamp 1698431365
transform 1 0 2240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_12
timestamp 1698431365
transform 1 0 2688 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_28
timestamp 1698431365
transform 1 0 4480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698431365
transform 1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_139
timestamp 1698431365
transform 1 0 16912 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_150
timestamp 1698431365
transform 1 0 18144 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_166
timestamp 1698431365
transform 1 0 19936 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_187
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_191
timestamp 1698431365
transform 1 0 22736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_193
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_200
timestamp 1698431365
transform 1 0 23744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_204
timestamp 1698431365
transform 1 0 24192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_208
timestamp 1698431365
transform 1 0 24640 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_240
timestamp 1698431365
transform 1 0 28224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_8
timestamp 1698431365
transform 1 0 2240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_12
timestamp 1698431365
transform 1 0 2688 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_44
timestamp 1698431365
transform 1 0 6272 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_60
timestamp 1698431365
transform 1 0 8064 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_68
timestamp 1698431365
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_104
timestamp 1698431365
transform 1 0 12992 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_120
timestamp 1698431365
transform 1 0 14784 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_124
timestamp 1698431365
transform 1 0 15232 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_131
timestamp 1698431365
transform 1 0 16016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_135
timestamp 1698431365
transform 1 0 16464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_137
timestamp 1698431365
transform 1 0 16688 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_168
timestamp 1698431365
transform 1 0 20160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_170
timestamp 1698431365
transform 1 0 20384 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_185
timestamp 1698431365
transform 1 0 22064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_189
timestamp 1698431365
transform 1 0 22512 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_218
timestamp 1698431365
transform 1 0 25760 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_250
timestamp 1698431365
transform 1 0 29344 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_266
timestamp 1698431365
transform 1 0 31136 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_274
timestamp 1698431365
transform 1 0 32032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_314
timestamp 1698431365
transform 1 0 36512 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_322
timestamp 1698431365
transform 1 0 37408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_324
timestamp 1698431365
transform 1 0 37632 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_8
timestamp 1698431365
transform 1 0 2240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_12
timestamp 1698431365
transform 1 0 2688 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_28
timestamp 1698431365
transform 1 0 4480 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_32
timestamp 1698431365
transform 1 0 4928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_111
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_142
timestamp 1698431365
transform 1 0 17248 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_165
timestamp 1698431365
transform 1 0 19824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_227
timestamp 1698431365
transform 1 0 26768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_235
timestamp 1698431365
transform 1 0 27664 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_239
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_241
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_249
timestamp 1698431365
transform 1 0 29232 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_256
timestamp 1698431365
transform 1 0 30016 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_288
timestamp 1698431365
transform 1 0 33600 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_304
timestamp 1698431365
transform 1 0 35392 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_312
timestamp 1698431365
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_8
timestamp 1698431365
transform 1 0 2240 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_40
timestamp 1698431365
transform 1 0 5824 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_56
timestamp 1698431365
transform 1 0 7616 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_64
timestamp 1698431365
transform 1 0 8512 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1698431365
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_104
timestamp 1698431365
transform 1 0 12992 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_108
timestamp 1698431365
transform 1 0 13440 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_110
timestamp 1698431365
transform 1 0 13664 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_192
timestamp 1698431365
transform 1 0 22848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_218
timestamp 1698431365
transform 1 0 25760 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_242
timestamp 1698431365
transform 1 0 28448 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_244
timestamp 1698431365
transform 1 0 28672 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_267
timestamp 1698431365
transform 1 0 31248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_271
timestamp 1698431365
transform 1 0 31696 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698431365
transform 1 0 36512 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_322
timestamp 1698431365
transform 1 0 37408 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_324
timestamp 1698431365
transform 1 0 37632 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_8
timestamp 1698431365
transform 1 0 2240 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_24
timestamp 1698431365
transform 1 0 4032 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698431365
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_185
timestamp 1698431365
transform 1 0 22064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_217
timestamp 1698431365
transform 1 0 25648 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_227
timestamp 1698431365
transform 1 0 26768 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_231
timestamp 1698431365
transform 1 0 27216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_233
timestamp 1698431365
transform 1 0 27440 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_240
timestamp 1698431365
transform 1 0 28224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_255
timestamp 1698431365
transform 1 0 29904 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_265
timestamp 1698431365
transform 1 0 31024 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_297
timestamp 1698431365
transform 1 0 34608 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_313
timestamp 1698431365
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_8
timestamp 1698431365
transform 1 0 2240 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_40
timestamp 1698431365
transform 1 0 5824 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_56
timestamp 1698431365
transform 1 0 7616 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_64
timestamp 1698431365
transform 1 0 8512 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698431365
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_88
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_92
timestamp 1698431365
transform 1 0 11648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_94
timestamp 1698431365
transform 1 0 11872 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_101
timestamp 1698431365
transform 1 0 12656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_105
timestamp 1698431365
transform 1 0 13104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_119
timestamp 1698431365
transform 1 0 14672 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_123
timestamp 1698431365
transform 1 0 15120 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_132
timestamp 1698431365
transform 1 0 16128 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_172
timestamp 1698431365
transform 1 0 20608 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_189
timestamp 1698431365
transform 1 0 22512 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_191
timestamp 1698431365
transform 1 0 22736 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_226
timestamp 1698431365
transform 1 0 26656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_250
timestamp 1698431365
transform 1 0 29344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_252
timestamp 1698431365
transform 1 0 29568 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_275
timestamp 1698431365
transform 1 0 32144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698431365
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_322
timestamp 1698431365
transform 1 0 37408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_324
timestamp 1698431365
transform 1 0 37632 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_14
timestamp 1698431365
transform 1 0 2912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_18
timestamp 1698431365
transform 1 0 3360 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_69
timestamp 1698431365
transform 1 0 9072 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_85
timestamp 1698431365
transform 1 0 10864 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_109
timestamp 1698431365
transform 1 0 13552 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_132
timestamp 1698431365
transform 1 0 16128 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_134
timestamp 1698431365
transform 1 0 16352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_149
timestamp 1698431365
transform 1 0 18032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_153
timestamp 1698431365
transform 1 0 18480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_155
timestamp 1698431365
transform 1 0 18704 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_158
timestamp 1698431365
transform 1 0 19040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_162
timestamp 1698431365
transform 1 0 19488 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_187
timestamp 1698431365
transform 1 0 22288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_191
timestamp 1698431365
transform 1 0 22736 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_202
timestamp 1698431365
transform 1 0 23968 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_206
timestamp 1698431365
transform 1 0 24416 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_213
timestamp 1698431365
transform 1 0 25200 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_221
timestamp 1698431365
transform 1 0 26096 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_257
timestamp 1698431365
transform 1 0 30128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_263
timestamp 1698431365
transform 1 0 30800 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_295
timestamp 1698431365
transform 1 0 34384 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_8
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_40
timestamp 1698431365
transform 1 0 5824 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_56
timestamp 1698431365
transform 1 0 7616 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_64
timestamp 1698431365
transform 1 0 8512 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_80
timestamp 1698431365
transform 1 0 10304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_106
timestamp 1698431365
transform 1 0 13216 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_120
timestamp 1698431365
transform 1 0 14784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_167
timestamp 1698431365
transform 1 0 20048 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_171
timestamp 1698431365
transform 1 0 20496 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_182
timestamp 1698431365
transform 1 0 21728 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_186
timestamp 1698431365
transform 1 0 22176 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_190
timestamp 1698431365
transform 1 0 22624 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_199
timestamp 1698431365
transform 1 0 23632 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_201
timestamp 1698431365
transform 1 0 23856 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698431365
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_216
timestamp 1698431365
transform 1 0 25536 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_218
timestamp 1698431365
transform 1 0 25760 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_239
timestamp 1698431365
transform 1 0 28112 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_269
timestamp 1698431365
transform 1 0 31472 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_273
timestamp 1698431365
transform 1 0 31920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698431365
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698431365
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_322
timestamp 1698431365
transform 1 0 37408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_324
timestamp 1698431365
transform 1 0 37632 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_8
timestamp 1698431365
transform 1 0 2240 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_24
timestamp 1698431365
transform 1 0 4032 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698431365
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_69
timestamp 1698431365
transform 1 0 9072 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_85
timestamp 1698431365
transform 1 0 10864 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_89
timestamp 1698431365
transform 1 0 11312 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_111
timestamp 1698431365
transform 1 0 13776 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_119
timestamp 1698431365
transform 1 0 14672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_132
timestamp 1698431365
transform 1 0 16128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_136
timestamp 1698431365
transform 1 0 16576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_144
timestamp 1698431365
transform 1 0 17472 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_148
timestamp 1698431365
transform 1 0 17920 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_161
timestamp 1698431365
transform 1 0 19376 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_185
timestamp 1698431365
transform 1 0 22064 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_187
timestamp 1698431365
transform 1 0 22288 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_190
timestamp 1698431365
transform 1 0 22624 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_225
timestamp 1698431365
transform 1 0 26544 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_239
timestamp 1698431365
transform 1 0 28112 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698431365
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_274
timestamp 1698431365
transform 1 0 32032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_278
timestamp 1698431365
transform 1 0 32480 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_310
timestamp 1698431365
transform 1 0 36064 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_8
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_40
timestamp 1698431365
transform 1 0 5824 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_56
timestamp 1698431365
transform 1 0 7616 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_64
timestamp 1698431365
transform 1 0 8512 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698431365
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698431365
transform 1 0 10304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_86
timestamp 1698431365
transform 1 0 10976 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_106
timestamp 1698431365
transform 1 0 13216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_108
timestamp 1698431365
transform 1 0 13440 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698431365
transform 1 0 16688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_161
timestamp 1698431365
transform 1 0 19376 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_168
timestamp 1698431365
transform 1 0 20160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_172
timestamp 1698431365
transform 1 0 20608 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_176
timestamp 1698431365
transform 1 0 21056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_188
timestamp 1698431365
transform 1 0 22400 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_192
timestamp 1698431365
transform 1 0 22848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_194
timestamp 1698431365
transform 1 0 23072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698431365
transform 1 0 24528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_216
timestamp 1698431365
transform 1 0 25536 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_231
timestamp 1698431365
transform 1 0 27216 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_235
timestamp 1698431365
transform 1 0 27664 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_248
timestamp 1698431365
transform 1 0 29120 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_252
timestamp 1698431365
transform 1 0 29568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_254
timestamp 1698431365
transform 1 0 29792 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_261
timestamp 1698431365
transform 1 0 30576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_265
timestamp 1698431365
transform 1 0 31024 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_273
timestamp 1698431365
transform 1 0 31920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698431365
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698431365
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_322
timestamp 1698431365
transform 1 0 37408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_324
timestamp 1698431365
transform 1 0 37632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_8
timestamp 1698431365
transform 1 0 2240 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_24
timestamp 1698431365
transform 1 0 4032 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698431365
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_69
timestamp 1698431365
transform 1 0 9072 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_77
timestamp 1698431365
transform 1 0 9968 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_81
timestamp 1698431365
transform 1 0 10416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_83
timestamp 1698431365
transform 1 0 10640 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_100
timestamp 1698431365
transform 1 0 12544 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_121
timestamp 1698431365
transform 1 0 14896 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_153
timestamp 1698431365
transform 1 0 18480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_161
timestamp 1698431365
transform 1 0 19376 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_168
timestamp 1698431365
transform 1 0 20160 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_200
timestamp 1698431365
transform 1 0 23744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_208
timestamp 1698431365
transform 1 0 24640 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_234
timestamp 1698431365
transform 1 0 27552 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_257
timestamp 1698431365
transform 1 0 30128 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_261
timestamp 1698431365
transform 1 0 30576 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_293
timestamp 1698431365
transform 1 0 34160 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_309
timestamp 1698431365
transform 1 0 35952 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_313
timestamp 1698431365
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_8
timestamp 1698431365
transform 1 0 2240 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_40
timestamp 1698431365
transform 1 0 5824 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_56
timestamp 1698431365
transform 1 0 7616 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_64
timestamp 1698431365
transform 1 0 8512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_88
timestamp 1698431365
transform 1 0 11200 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_96
timestamp 1698431365
transform 1 0 12096 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_103
timestamp 1698431365
transform 1 0 12880 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_111
timestamp 1698431365
transform 1 0 13776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_115
timestamp 1698431365
transform 1 0 14224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_117
timestamp 1698431365
transform 1 0 14448 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_130
timestamp 1698431365
transform 1 0 15904 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698431365
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_144
timestamp 1698431365
transform 1 0 17472 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_151
timestamp 1698431365
transform 1 0 18256 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_172
timestamp 1698431365
transform 1 0 20608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_176
timestamp 1698431365
transform 1 0 21056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_196
timestamp 1698431365
transform 1 0 23296 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_216
timestamp 1698431365
transform 1 0 25536 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_239
timestamp 1698431365
transform 1 0 28112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_243
timestamp 1698431365
transform 1 0 28560 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_260
timestamp 1698431365
transform 1 0 30464 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698431365
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_322
timestamp 1698431365
transform 1 0 37408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_324
timestamp 1698431365
transform 1 0 37632 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_14
timestamp 1698431365
transform 1 0 2912 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_30
timestamp 1698431365
transform 1 0 4704 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_123
timestamp 1698431365
transform 1 0 15120 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_131
timestamp 1698431365
transform 1 0 16016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_135
timestamp 1698431365
transform 1 0 16464 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_138
timestamp 1698431365
transform 1 0 16800 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_158
timestamp 1698431365
transform 1 0 19040 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_167
timestamp 1698431365
transform 1 0 20048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_179
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_190
timestamp 1698431365
transform 1 0 22624 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_206
timestamp 1698431365
transform 1 0 24416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_236
timestamp 1698431365
transform 1 0 27776 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_269
timestamp 1698431365
transform 1 0 31472 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_301
timestamp 1698431365
transform 1 0 35056 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_309
timestamp 1698431365
transform 1 0 35952 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_313
timestamp 1698431365
transform 1 0 36400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_8
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_40
timestamp 1698431365
transform 1 0 5824 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_56
timestamp 1698431365
transform 1 0 7616 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_64
timestamp 1698431365
transform 1 0 8512 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698431365
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_144
timestamp 1698431365
transform 1 0 17472 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_151
timestamp 1698431365
transform 1 0 18256 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_159
timestamp 1698431365
transform 1 0 19152 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_178
timestamp 1698431365
transform 1 0 21280 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_180
timestamp 1698431365
transform 1 0 21504 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_203
timestamp 1698431365
transform 1 0 24080 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698431365
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_218
timestamp 1698431365
transform 1 0 25760 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_222
timestamp 1698431365
transform 1 0 26208 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_244
timestamp 1698431365
transform 1 0 28672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_248
timestamp 1698431365
transform 1 0 29120 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_256
timestamp 1698431365
transform 1 0 30016 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_259
timestamp 1698431365
transform 1 0 30352 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_275
timestamp 1698431365
transform 1 0 32144 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698431365
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_322
timestamp 1698431365
transform 1 0 37408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_324
timestamp 1698431365
transform 1 0 37632 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_8
timestamp 1698431365
transform 1 0 2240 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_24
timestamp 1698431365
transform 1 0 4032 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_123
timestamp 1698431365
transform 1 0 15120 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_131
timestamp 1698431365
transform 1 0 16016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_135
timestamp 1698431365
transform 1 0 16464 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_138
timestamp 1698431365
transform 1 0 16800 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_158
timestamp 1698431365
transform 1 0 19040 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_165
timestamp 1698431365
transform 1 0 19824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_169
timestamp 1698431365
transform 1 0 20272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698431365
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_191
timestamp 1698431365
transform 1 0 22736 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_195
timestamp 1698431365
transform 1 0 23184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_197
timestamp 1698431365
transform 1 0 23408 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_212
timestamp 1698431365
transform 1 0 25088 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_216
timestamp 1698431365
transform 1 0 25536 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_261
timestamp 1698431365
transform 1 0 30576 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_293
timestamp 1698431365
transform 1 0 34160 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_309
timestamp 1698431365
transform 1 0 35952 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_313
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_8
timestamp 1698431365
transform 1 0 2240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_12
timestamp 1698431365
transform 1 0 2688 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_44
timestamp 1698431365
transform 1 0 6272 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698431365
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_144
timestamp 1698431365
transform 1 0 17472 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_173
timestamp 1698431365
transform 1 0 20720 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_184
timestamp 1698431365
transform 1 0 21952 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_188
timestamp 1698431365
transform 1 0 22400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_192
timestamp 1698431365
transform 1 0 22848 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_205
timestamp 1698431365
transform 1 0 24304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_228
timestamp 1698431365
transform 1 0 26880 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_232
timestamp 1698431365
transform 1 0 27328 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_234
timestamp 1698431365
transform 1 0 27552 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_251
timestamp 1698431365
transform 1 0 29456 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_255
timestamp 1698431365
transform 1 0 29904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_259
timestamp 1698431365
transform 1 0 30352 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_275
timestamp 1698431365
transform 1 0 32144 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698431365
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_322
timestamp 1698431365
transform 1 0 37408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_324
timestamp 1698431365
transform 1 0 37632 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_8
timestamp 1698431365
transform 1 0 2240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_12
timestamp 1698431365
transform 1 0 2688 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_139
timestamp 1698431365
transform 1 0 16912 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_143
timestamp 1698431365
transform 1 0 17360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_151
timestamp 1698431365
transform 1 0 18256 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_161
timestamp 1698431365
transform 1 0 19376 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_168
timestamp 1698431365
transform 1 0 20160 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698431365
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_199
timestamp 1698431365
transform 1 0 23632 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_215
timestamp 1698431365
transform 1 0 25424 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_228
timestamp 1698431365
transform 1 0 26880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_232
timestamp 1698431365
transform 1 0 27328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_236
timestamp 1698431365
transform 1 0 27776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_238
timestamp 1698431365
transform 1 0 28000 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_253
timestamp 1698431365
transform 1 0 29680 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_285
timestamp 1698431365
transform 1 0 33264 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_301
timestamp 1698431365
transform 1 0 35056 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_309
timestamp 1698431365
transform 1 0 35952 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698431365
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698431365
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_8
timestamp 1698431365
transform 1 0 2240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_12
timestamp 1698431365
transform 1 0 2688 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_44
timestamp 1698431365
transform 1 0 6272 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698431365
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_174
timestamp 1698431365
transform 1 0 20832 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_182
timestamp 1698431365
transform 1 0 21728 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_186
timestamp 1698431365
transform 1 0 22176 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_189
timestamp 1698431365
transform 1 0 22512 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_205
timestamp 1698431365
transform 1 0 24304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698431365
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698431365
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_8
timestamp 1698431365
transform 1 0 2240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_12
timestamp 1698431365
transform 1 0 2688 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698431365
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698431365
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_314
timestamp 1698431365
transform 1 0 36512 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_322
timestamp 1698431365
transform 1 0 37408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_324
timestamp 1698431365
transform 1 0 37632 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_321
timestamp 1698431365
transform 1 0 37296 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_314
timestamp 1698431365
transform 1 0 36512 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_322
timestamp 1698431365
transform 1 0 37408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_324
timestamp 1698431365
transform 1 0 37632 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_321
timestamp 1698431365
transform 1 0 37296 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_314
timestamp 1698431365
transform 1 0 36512 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_322
timestamp 1698431365
transform 1 0 37408 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_314
timestamp 1698431365
transform 1 0 36512 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_318
timestamp 1698431365
transform 1 0 36960 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_321
timestamp 1698431365
transform 1 0 37296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_314
timestamp 1698431365
transform 1 0 36512 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_322
timestamp 1698431365
transform 1 0 37408 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_104
timestamp 1698431365
transform 1 0 12992 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_120
timestamp 1698431365
transform 1 0 14784 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_126
timestamp 1698431365
transform 1 0 15456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_130
timestamp 1698431365
transform 1 0 15904 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_174
timestamp 1698431365
transform 1 0 20832 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_178
timestamp 1698431365
transform 1 0 21280 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_181
timestamp 1698431365
transform 1 0 21616 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_197
timestamp 1698431365
transform 1 0 23408 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_205
timestamp 1698431365
transform 1 0 24304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_209
timestamp 1698431365
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_218
timestamp 1698431365
transform 1 0 25760 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_250
timestamp 1698431365
transform 1 0 29344 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_266
timestamp 1698431365
transform 1 0 31136 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_274
timestamp 1698431365
transform 1 0 32032 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_278
timestamp 1698431365
transform 1 0 32480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_314
timestamp 1698431365
transform 1 0 36512 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_318
timestamp 1698431365
transform 1 0 36960 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_321
timestamp 1698431365
transform 1 0 37296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_36
timestamp 1698431365
transform 1 0 5376 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_70
timestamp 1698431365
transform 1 0 9184 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_112
timestamp 1698431365
transform 1 0 13888 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_116
timestamp 1698431365
transform 1 0 14336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_138
timestamp 1698431365
transform 1 0 16800 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_172
timestamp 1698431365
transform 1 0 20608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_199
timestamp 1698431365
transform 1 0 23632 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_203
timestamp 1698431365
transform 1 0 24080 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_224
timestamp 1698431365
transform 1 0 26432 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_232
timestamp 1698431365
transform 1 0 27328 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_236
timestamp 1698431365
transform 1 0 27776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_240
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_274
timestamp 1698431365
transform 1 0 32032 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_290
timestamp 1698431365
transform 1 0 33824 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_298
timestamp 1698431365
transform 1 0 34720 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_302
timestamp 1698431365
transform 1 0 35168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_308
timestamp 1698431365
transform 1 0 35840 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_310
timestamp 1698431365
transform 1 0 36064 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698431365
transform -1 0 26432 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input2
timestamp 1698431365
transform 1 0 15232 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 25088 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform -1 0 37744 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698431365
transform -1 0 38416 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 38416 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 38416 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input10
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input11
timestamp 1698431365
transform 1 0 14560 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 21616 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input13
timestamp 1698431365
transform 1 0 16240 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input14
timestamp 1698431365
transform -1 0 37744 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input15
timestamp 1698431365
transform -1 0 38416 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input16
timestamp 1698431365
transform -1 0 38416 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 38416 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform -1 0 26432 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 27104 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  net99_2
timestamp 1698431365
transform 1 0 17472 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output23
timestamp 1698431365
transform 1 0 18368 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output24
timestamp 1698431365
transform 1 0 19040 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output25
timestamp 1698431365
transform -1 0 16912 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output26
timestamp 1698431365
transform 1 0 15904 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output27
timestamp 1698431365
transform 1 0 19712 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output28
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output29
timestamp 1698431365
transform 1 0 37072 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output30
timestamp 1698431365
transform 1 0 37744 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output31
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output32
timestamp 1698431365
transform 1 0 37744 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output33
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output34
timestamp 1698431365
transform -1 0 2240 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output35
timestamp 1698431365
transform -1 0 2240 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output36
timestamp 1698431365
transform -1 0 2240 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output37
timestamp 1698431365
transform -1 0 23632 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output38
timestamp 1698431365
transform -1 0 15904 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output39
timestamp 1698431365
transform -1 0 25760 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output40
timestamp 1698431365
transform -1 0 22960 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output41
timestamp 1698431365
transform -1 0 25088 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output42
timestamp 1698431365
transform 1 0 37744 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output43
timestamp 1698431365
transform 1 0 37744 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output44
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output45
timestamp 1698431365
transform 1 0 37744 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output46
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output47
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output48
timestamp 1698431365
transform 1 0 19712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output49
timestamp 1698431365
transform 1 0 18368 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output50
timestamp 1698431365
transform -1 0 23632 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output51
timestamp 1698431365
transform 1 0 37744 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output52
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output53
timestamp 1698431365
transform 1 0 37744 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output54
timestamp 1698431365
transform 1 0 37744 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output55
timestamp 1698431365
transform -1 0 2240 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output56
timestamp 1698431365
transform -1 0 2240 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output57
timestamp 1698431365
transform -1 0 2240 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output58
timestamp 1698431365
transform 1 0 37072 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output59
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output60
timestamp 1698431365
transform 1 0 17024 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output61
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output62
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output63
timestamp 1698431365
transform 1 0 37744 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output64
timestamp 1698431365
transform 1 0 37744 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output65
timestamp 1698431365
transform 1 0 37744 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output66
timestamp 1698431365
transform 1 0 37072 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output67
timestamp 1698431365
transform 1 0 37744 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output68
timestamp 1698431365
transform 1 0 37744 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output69
timestamp 1698431365
transform 1 0 37072 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output70
timestamp 1698431365
transform 1 0 37072 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output71
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output72
timestamp 1698431365
transform 1 0 37744 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output73
timestamp 1698431365
transform 1 0 37744 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output74
timestamp 1698431365
transform 1 0 37744 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output75
timestamp 1698431365
transform 1 0 37744 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output76
timestamp 1698431365
transform -1 0 2240 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output77
timestamp 1698431365
transform -1 0 2240 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output78
timestamp 1698431365
transform -1 0 2240 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output79
timestamp 1698431365
transform -1 0 21616 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output80
timestamp 1698431365
transform 1 0 15904 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output81
timestamp 1698431365
transform 1 0 19040 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output82
timestamp 1698431365
transform 1 0 37744 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output83
timestamp 1698431365
transform 1 0 17696 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output84
timestamp 1698431365
transform 1 0 37744 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output85
timestamp 1698431365
transform 1 0 37072 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output86
timestamp 1698431365
transform 1 0 37744 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output87
timestamp 1698431365
transform 1 0 37744 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output88
timestamp 1698431365
transform -1 0 22288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output89
timestamp 1698431365
transform -1 0 21616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output90
timestamp 1698431365
transform 1 0 17696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output91
timestamp 1698431365
transform -1 0 22960 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output92
timestamp 1698431365
transform 1 0 37744 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output93
timestamp 1698431365
transform 1 0 37744 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output94
timestamp 1698431365
transform 1 0 37744 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output95
timestamp 1698431365
transform 1 0 37744 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output96
timestamp 1698431365
transform 1 0 37744 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output97
timestamp 1698431365
transform -1 0 2240 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output98
timestamp 1698431365
transform -1 0 2240 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output99
timestamp 1698431365
transform -1 0 2912 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output100
timestamp 1698431365
transform 1 0 37744 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output101
timestamp 1698431365
transform -1 0 27776 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output102
timestamp 1698431365
transform -1 0 25760 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output103
timestamp 1698431365
transform -1 0 2240 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output104
timestamp 1698431365
transform -1 0 2912 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output105
timestamp 1698431365
transform -1 0 2240 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output106
timestamp 1698431365
transform 1 0 17024 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_43 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_44
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 38640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_45
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 38640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_46
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_47
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_48
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 38640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_49
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 38640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_50
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 38640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_51
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_52
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 38640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_53
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 38640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 38640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 38640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 38640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 38640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 38640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 38640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 38640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 38640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 38640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 38640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 38640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 38640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 38640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 38640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 38640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 38640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 38640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 38640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 38640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_86 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_87
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_88
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_89
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_95
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_96
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_97
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_98
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_99
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_100
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_101
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_102
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_103
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_104
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_105
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_106
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_107
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_108
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_109
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_110
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_111
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_112
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_113
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_114
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_115
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_116
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_117
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_118
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_119
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_120
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_121
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_122
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_123
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_124
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_125
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_126
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_127
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_128
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_129
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_130
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_131
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_132
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_133
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_134
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_135
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_136
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_137
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_138
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_139
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_140
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_141
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_142
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_143
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_144
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_145
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_146
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_147
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_148
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_149
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_150
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_151
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_152
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_153
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_154
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_155
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_156
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_157
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_158
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_159
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_160
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_161
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_162
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_163
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_164
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_165
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_166
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_167
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_168
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_169
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_170
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_171
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_172
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_173
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_174
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_175
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_176
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_177
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_178
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_179
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_180
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_181
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_182
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_183
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_184
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_185
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_186
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_187
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_188
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_189
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_190
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_191
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_192
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_193
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_194
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_195
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_196
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_197
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_198
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_199
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_200
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_201
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_202
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_203
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_204
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_205
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_206
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_207
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_208
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_209
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_210
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_211
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_212
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_213
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_214
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_215
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_216
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_217
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_218
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_219
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_220
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_221
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_222
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_223
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_224
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_225
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_226
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_227
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_228
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_229
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_230
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_231
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_232
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_233
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_234
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_235
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_236
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_237
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_238
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_239
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_240
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_241
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_242
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_243
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_244
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_245
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_246
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_247
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_248
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_249
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_250
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_251
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_252
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_253
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_254
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_255
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_256
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_257
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_258
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_259
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_260
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_261
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_262
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_263
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_264
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_265
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_266
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_267
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_268
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_269
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_270
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_271
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_272
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_273
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_274
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_275
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_276
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_277
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_278
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_279
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_280
timestamp 1698431365
transform 1 0 8960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_281
timestamp 1698431365
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_282
timestamp 1698431365
transform 1 0 16576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_283
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698431365
transform 1 0 24192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698431365
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698431365
transform 1 0 31808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 310 870
<< labels >>
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 24864 39200 24976 40000 0 FreeSans 448 90 0 0 in[0]
port 1 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 in[10]
port 2 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 in[11]
port 3 nsew signal input
flabel metal3 s 39200 2688 40000 2800 0 FreeSans 448 0 0 0 in[12]
port 4 nsew signal input
flabel metal3 s 39200 8064 40000 8176 0 FreeSans 448 0 0 0 in[13]
port 5 nsew signal input
flabel metal3 s 39200 9408 40000 9520 0 FreeSans 448 0 0 0 in[14]
port 6 nsew signal input
flabel metal3 s 39200 11424 40000 11536 0 FreeSans 448 0 0 0 in[15]
port 7 nsew signal input
flabel metal3 s 0 12768 800 12880 0 FreeSans 448 0 0 0 in[16]
port 8 nsew signal input
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 in[17]
port 9 nsew signal input
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 in[18]
port 10 nsew signal input
flabel metal2 s 14784 39200 14896 40000 0 FreeSans 448 90 0 0 in[1]
port 11 nsew signal input
flabel metal2 s 21504 39200 21616 40000 0 FreeSans 448 90 0 0 in[2]
port 12 nsew signal input
flabel metal2 s 16128 39200 16240 40000 0 FreeSans 448 90 0 0 in[3]
port 13 nsew signal input
flabel metal3 s 39200 36960 40000 37072 0 FreeSans 448 0 0 0 in[4]
port 14 nsew signal input
flabel metal3 s 39200 32256 40000 32368 0 FreeSans 448 0 0 0 in[5]
port 15 nsew signal input
flabel metal3 s 39200 35616 40000 35728 0 FreeSans 448 0 0 0 in[6]
port 16 nsew signal input
flabel metal3 s 39200 25536 40000 25648 0 FreeSans 448 0 0 0 in[7]
port 17 nsew signal input
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 in[8]
port 18 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 in[9]
port 19 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 proj_clk[0]
port 20 nsew signal tristate
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 proj_clk[1]
port 21 nsew signal tristate
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 proj_clk[2]
port 22 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 proj_clk[3]
port 23 nsew signal tristate
flabel metal2 s 20160 39200 20272 40000 0 FreeSans 448 90 0 0 proj_in[0]
port 24 nsew signal tristate
flabel metal3 s 39200 10752 40000 10864 0 FreeSans 448 0 0 0 proj_in[10]
port 25 nsew signal tristate
flabel metal3 s 39200 12096 40000 12208 0 FreeSans 448 0 0 0 proj_in[11]
port 26 nsew signal tristate
flabel metal3 s 39200 15456 40000 15568 0 FreeSans 448 0 0 0 proj_in[12]
port 27 nsew signal tristate
flabel metal3 s 39200 12768 40000 12880 0 FreeSans 448 0 0 0 proj_in[13]
port 28 nsew signal tristate
flabel metal3 s 39200 8736 40000 8848 0 FreeSans 448 0 0 0 proj_in[14]
port 29 nsew signal tristate
flabel metal3 s 39200 14112 40000 14224 0 FreeSans 448 0 0 0 proj_in[15]
port 30 nsew signal tristate
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 proj_in[16]
port 31 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 proj_in[17]
port 32 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 proj_in[18]
port 33 nsew signal tristate
flabel metal2 s 22848 39200 22960 40000 0 FreeSans 448 90 0 0 proj_in[19]
port 34 nsew signal tristate
flabel metal2 s 15456 39200 15568 40000 0 FreeSans 448 90 0 0 proj_in[1]
port 35 nsew signal tristate
flabel metal2 s 24192 39200 24304 40000 0 FreeSans 448 90 0 0 proj_in[20]
port 36 nsew signal tristate
flabel metal2 s 22176 39200 22288 40000 0 FreeSans 448 90 0 0 proj_in[21]
port 37 nsew signal tristate
flabel metal2 s 23520 39200 23632 40000 0 FreeSans 448 90 0 0 proj_in[22]
port 38 nsew signal tristate
flabel metal3 s 39200 22176 40000 22288 0 FreeSans 448 0 0 0 proj_in[23]
port 39 nsew signal tristate
flabel metal3 s 39200 26208 40000 26320 0 FreeSans 448 0 0 0 proj_in[24]
port 40 nsew signal tristate
flabel metal3 s 39200 36288 40000 36400 0 FreeSans 448 0 0 0 proj_in[25]
port 41 nsew signal tristate
flabel metal3 s 39200 28896 40000 29008 0 FreeSans 448 0 0 0 proj_in[26]
port 42 nsew signal tristate
flabel metal3 s 39200 18816 40000 18928 0 FreeSans 448 0 0 0 proj_in[27]
port 43 nsew signal tristate
flabel metal3 s 39200 17472 40000 17584 0 FreeSans 448 0 0 0 proj_in[28]
port 44 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 proj_in[29]
port 45 nsew signal tristate
flabel metal2 s 18816 39200 18928 40000 0 FreeSans 448 90 0 0 proj_in[2]
port 46 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 proj_in[30]
port 47 nsew signal tristate
flabel metal3 s 39200 19488 40000 19600 0 FreeSans 448 0 0 0 proj_in[31]
port 48 nsew signal tristate
flabel metal3 s 39200 20160 40000 20272 0 FreeSans 448 0 0 0 proj_in[32]
port 49 nsew signal tristate
flabel metal3 s 39200 6048 40000 6160 0 FreeSans 448 0 0 0 proj_in[33]
port 50 nsew signal tristate
flabel metal3 s 39200 6720 40000 6832 0 FreeSans 448 0 0 0 proj_in[34]
port 51 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 proj_in[35]
port 52 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 proj_in[36]
port 53 nsew signal tristate
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 proj_in[37]
port 54 nsew signal tristate
flabel metal3 s 39200 21504 40000 21616 0 FreeSans 448 0 0 0 proj_in[38]
port 55 nsew signal tristate
flabel metal3 s 39200 23520 40000 23632 0 FreeSans 448 0 0 0 proj_in[39]
port 56 nsew signal tristate
flabel metal2 s 17472 39200 17584 40000 0 FreeSans 448 90 0 0 proj_in[3]
port 57 nsew signal tristate
flabel metal3 s 39200 28224 40000 28336 0 FreeSans 448 0 0 0 proj_in[40]
port 58 nsew signal tristate
flabel metal3 s 39200 29568 40000 29680 0 FreeSans 448 0 0 0 proj_in[41]
port 59 nsew signal tristate
flabel metal3 s 39200 20832 40000 20944 0 FreeSans 448 0 0 0 proj_in[42]
port 60 nsew signal tristate
flabel metal3 s 39200 24864 40000 24976 0 FreeSans 448 0 0 0 proj_in[43]
port 61 nsew signal tristate
flabel metal3 s 39200 22848 40000 22960 0 FreeSans 448 0 0 0 proj_in[44]
port 62 nsew signal tristate
flabel metal3 s 39200 26880 40000 26992 0 FreeSans 448 0 0 0 proj_in[45]
port 63 nsew signal tristate
flabel metal3 s 39200 4032 40000 4144 0 FreeSans 448 0 0 0 proj_in[46]
port 64 nsew signal tristate
flabel metal3 s 39200 18144 40000 18256 0 FreeSans 448 0 0 0 proj_in[47]
port 65 nsew signal tristate
flabel metal3 s 39200 7392 40000 7504 0 FreeSans 448 0 0 0 proj_in[48]
port 66 nsew signal tristate
flabel metal3 s 39200 16800 40000 16912 0 FreeSans 448 0 0 0 proj_in[49]
port 67 nsew signal tristate
flabel metal3 s 39200 32928 40000 33040 0 FreeSans 448 0 0 0 proj_in[4]
port 68 nsew signal tristate
flabel metal3 s 39200 3360 40000 3472 0 FreeSans 448 0 0 0 proj_in[50]
port 69 nsew signal tristate
flabel metal3 s 39200 24192 40000 24304 0 FreeSans 448 0 0 0 proj_in[51]
port 70 nsew signal tristate
flabel metal3 s 39200 4704 40000 4816 0 FreeSans 448 0 0 0 proj_in[52]
port 71 nsew signal tristate
flabel metal3 s 39200 5376 40000 5488 0 FreeSans 448 0 0 0 proj_in[53]
port 72 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 proj_in[54]
port 73 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 proj_in[55]
port 74 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 proj_in[56]
port 75 nsew signal tristate
flabel metal2 s 20832 39200 20944 40000 0 FreeSans 448 90 0 0 proj_in[57]
port 76 nsew signal tristate
flabel metal2 s 16800 39200 16912 40000 0 FreeSans 448 90 0 0 proj_in[58]
port 77 nsew signal tristate
flabel metal2 s 19488 39200 19600 40000 0 FreeSans 448 90 0 0 proj_in[59]
port 78 nsew signal tristate
flabel metal3 s 39200 33600 40000 33712 0 FreeSans 448 0 0 0 proj_in[5]
port 79 nsew signal tristate
flabel metal2 s 18144 39200 18256 40000 0 FreeSans 448 90 0 0 proj_in[60]
port 80 nsew signal tristate
flabel metal3 s 39200 34944 40000 35056 0 FreeSans 448 0 0 0 proj_in[61]
port 81 nsew signal tristate
flabel metal3 s 39200 31584 40000 31696 0 FreeSans 448 0 0 0 proj_in[62]
port 82 nsew signal tristate
flabel metal3 s 39200 30912 40000 31024 0 FreeSans 448 0 0 0 proj_in[63]
port 83 nsew signal tristate
flabel metal3 s 39200 30240 40000 30352 0 FreeSans 448 0 0 0 proj_in[64]
port 84 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 proj_in[65]
port 85 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 proj_in[66]
port 86 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 proj_in[67]
port 87 nsew signal tristate
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 proj_in[68]
port 88 nsew signal tristate
flabel metal3 s 39200 10080 40000 10192 0 FreeSans 448 0 0 0 proj_in[69]
port 89 nsew signal tristate
flabel metal3 s 39200 34272 40000 34384 0 FreeSans 448 0 0 0 proj_in[6]
port 90 nsew signal tristate
flabel metal3 s 39200 13440 40000 13552 0 FreeSans 448 0 0 0 proj_in[70]
port 91 nsew signal tristate
flabel metal3 s 39200 16128 40000 16240 0 FreeSans 448 0 0 0 proj_in[71]
port 92 nsew signal tristate
flabel metal3 s 39200 14784 40000 14896 0 FreeSans 448 0 0 0 proj_in[72]
port 93 nsew signal tristate
flabel metal3 s 0 14784 800 14896 0 FreeSans 448 0 0 0 proj_in[73]
port 94 nsew signal tristate
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 proj_in[74]
port 95 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 proj_in[75]
port 96 nsew signal tristate
flabel metal3 s 39200 27552 40000 27664 0 FreeSans 448 0 0 0 proj_in[7]
port 97 nsew signal tristate
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 proj_in[8]
port 98 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 proj_in[9]
port 99 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 proj_rst_n[0]
port 100 nsew signal tristate
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 proj_rst_n[1]
port 101 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 proj_rst_n[2]
port 102 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 proj_rst_n[3]
port 103 nsew signal tristate
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 rst_n
port 104 nsew signal input
flabel metal3 s 0 13440 800 13552 0 FreeSans 448 0 0 0 sel[0]
port 105 nsew signal input
flabel metal3 s 0 14112 800 14224 0 FreeSans 448 0 0 0 sel[1]
port 106 nsew signal input
flabel metal4 s 5846 3076 6166 36908 0 FreeSans 1280 90 0 0 vdd
port 107 nsew power bidirectional
flabel metal4 s 15170 3076 15490 36908 0 FreeSans 1280 90 0 0 vdd
port 107 nsew power bidirectional
flabel metal4 s 24494 3076 24814 36908 0 FreeSans 1280 90 0 0 vdd
port 107 nsew power bidirectional
flabel metal4 s 33818 3076 34138 36908 0 FreeSans 1280 90 0 0 vdd
port 107 nsew power bidirectional
flabel metal4 s 10508 3076 10828 36908 0 FreeSans 1280 90 0 0 vss
port 108 nsew ground bidirectional
flabel metal4 s 19832 3076 20152 36908 0 FreeSans 1280 90 0 0 vss
port 108 nsew ground bidirectional
flabel metal4 s 29156 3076 29476 36908 0 FreeSans 1280 90 0 0 vss
port 108 nsew ground bidirectional
flabel metal4 s 38480 3076 38800 36908 0 FreeSans 1280 90 0 0 vss
port 108 nsew ground bidirectional
rlabel metal1 19992 36848 19992 36848 0 vdd
rlabel via1 20072 36064 20072 36064 0 vss
rlabel metal2 15792 18424 15792 18424 0 _000_
rlabel metal3 16856 18312 16856 18312 0 _001_
rlabel metal2 18984 19656 18984 19656 0 _002_
rlabel metal2 19208 20216 19208 20216 0 _003_
rlabel metal3 19096 24472 19096 24472 0 _004_
rlabel metal3 20216 24696 20216 24696 0 _005_
rlabel metal2 17976 24416 17976 24416 0 _006_
rlabel metal2 18984 25200 18984 25200 0 _007_
rlabel metal2 18312 24752 18312 24752 0 _008_
rlabel metal2 29400 24304 29400 24304 0 _009_
rlabel metal2 28392 25200 28392 25200 0 _010_
rlabel metal2 28112 23800 28112 23800 0 _011_
rlabel metal2 29176 24920 29176 24920 0 _012_
rlabel metal2 29904 23800 29904 23800 0 _013_
rlabel metal2 22792 16016 22792 16016 0 _014_
rlabel metal2 23352 13216 23352 13216 0 _015_
rlabel metal3 24752 13720 24752 13720 0 _016_
rlabel metal3 24976 15960 24976 15960 0 _017_
rlabel metal3 24528 15288 24528 15288 0 _018_
rlabel metal3 30520 16632 30520 16632 0 _019_
rlabel metal2 31472 16856 31472 16856 0 _020_
rlabel metal2 30576 15288 30576 15288 0 _021_
rlabel metal2 30520 16352 30520 16352 0 _022_
rlabel metal2 29512 14784 29512 14784 0 _023_
rlabel metal2 11984 20776 11984 20776 0 _024_
rlabel metal2 12264 19488 12264 19488 0 _025_
rlabel metal2 11536 20216 11536 20216 0 _026_
rlabel metal2 12432 21000 12432 21000 0 _027_
rlabel metal2 19096 20496 19096 20496 0 _028_
rlabel metal2 19992 20720 19992 20720 0 _029_
rlabel via2 21224 23128 21224 23128 0 _030_
rlabel metal2 19768 18872 19768 18872 0 _031_
rlabel metal2 21336 24864 21336 24864 0 _032_
rlabel metal3 22624 25480 22624 25480 0 _033_
rlabel metal2 22568 24416 22568 24416 0 _034_
rlabel metal2 21784 25144 21784 25144 0 _035_
rlabel metal2 22624 23352 22624 23352 0 _036_
rlabel metal2 29064 22064 29064 22064 0 _037_
rlabel metal3 28336 21672 28336 21672 0 _038_
rlabel metal2 29960 21280 29960 21280 0 _039_
rlabel metal2 27944 21056 27944 21056 0 _040_
rlabel metal2 30128 22232 30128 22232 0 _041_
rlabel metal2 29624 21840 29624 21840 0 _042_
rlabel metal2 21000 18760 21000 18760 0 _043_
rlabel metal3 20664 18424 20664 18424 0 _044_
rlabel metal2 21560 18872 21560 18872 0 _045_
rlabel metal2 20552 17696 20552 17696 0 _046_
rlabel metal2 19656 17360 19656 17360 0 _047_
rlabel metal2 21840 16856 21840 16856 0 _048_
rlabel metal2 26600 19320 26600 19320 0 _049_
rlabel metal2 27496 19656 27496 19656 0 _050_
rlabel metal2 27944 18536 27944 18536 0 _051_
rlabel metal2 27944 19712 27944 19712 0 _052_
rlabel metal2 26488 17920 26488 17920 0 _053_
rlabel metal2 28112 17528 28112 17528 0 _054_
rlabel metal2 14168 20384 14168 20384 0 _055_
rlabel metal2 14280 20384 14280 20384 0 _056_
rlabel metal2 15456 19208 15456 19208 0 _057_
rlabel metal2 14728 20440 14728 20440 0 _058_
rlabel metal2 14784 21000 14784 21000 0 _059_
rlabel metal2 22792 20608 22792 20608 0 _060_
rlabel metal2 21896 21952 21896 21952 0 _061_
rlabel metal3 19040 18424 19040 18424 0 _062_
rlabel metal2 23464 19656 23464 19656 0 _063_
rlabel metal2 22008 21952 22008 21952 0 _064_
rlabel metal2 22232 20272 22232 20272 0 _065_
rlabel metal2 22456 22848 22456 22848 0 _066_
rlabel metal2 22232 21280 22232 21280 0 _067_
rlabel metal2 22456 22008 22456 22008 0 _068_
rlabel metal2 25256 21952 25256 21952 0 _069_
rlabel metal3 24024 21560 24024 21560 0 _070_
rlabel metal2 26208 20664 26208 20664 0 _071_
rlabel metal2 24136 21056 24136 21056 0 _072_
rlabel metal2 25816 21896 25816 21896 0 _073_
rlabel metal2 27104 22232 27104 22232 0 _074_
rlabel metal3 23576 19096 23576 19096 0 _075_
rlabel metal2 23464 18872 23464 18872 0 _076_
rlabel metal2 24696 18984 24696 18984 0 _077_
rlabel metal2 23800 18144 23800 18144 0 _078_
rlabel metal2 24024 17136 24024 17136 0 _079_
rlabel metal2 23912 16576 23912 16576 0 _080_
rlabel metal3 25704 18872 25704 18872 0 _081_
rlabel metal2 29064 18760 29064 18760 0 _082_
rlabel metal2 31360 19096 31360 19096 0 _083_
rlabel metal2 30072 19712 30072 19712 0 _084_
rlabel metal2 30800 18424 30800 18424 0 _085_
rlabel metal2 29568 17640 29568 17640 0 _086_
rlabel metal2 14056 18032 14056 18032 0 _087_
rlabel metal2 14168 18144 14168 18144 0 _088_
rlabel metal2 13720 17304 13720 17304 0 _089_
rlabel metal2 14616 18760 14616 18760 0 _090_
rlabel metal3 14896 17640 14896 17640 0 _091_
rlabel metal3 16352 16856 16352 16856 0 _092_
rlabel metal2 25424 16856 25424 16856 0 _093_
rlabel metal3 18144 22344 18144 22344 0 _094_
rlabel metal2 19320 22848 19320 22848 0 _095_
rlabel metal2 18312 22848 18312 22848 0 _096_
rlabel metal2 20328 21504 20328 21504 0 _097_
rlabel metal2 17976 21840 17976 21840 0 _098_
rlabel metal2 26040 24304 26040 24304 0 _099_
rlabel metal2 26656 24920 26656 24920 0 _100_
rlabel metal2 23800 23744 23800 23744 0 _101_
rlabel metal2 25816 25200 25816 25200 0 _102_
rlabel metal2 26544 23800 26544 23800 0 _103_
rlabel metal3 19096 16296 19096 16296 0 _104_
rlabel metal2 20776 13664 20776 13664 0 _105_
rlabel metal3 21336 12936 21336 12936 0 _106_
rlabel metal2 19208 16576 19208 16576 0 _107_
rlabel metal2 24360 15568 24360 15568 0 _108_
rlabel metal2 25592 16856 25592 16856 0 _109_
rlabel metal2 28000 16856 28000 16856 0 _110_
rlabel metal2 27720 15736 27720 15736 0 _111_
rlabel metal2 26208 16072 26208 16072 0 _112_
rlabel metal2 27104 14504 27104 14504 0 _113_
rlabel metal3 12376 18200 12376 18200 0 _114_
rlabel metal2 12320 16856 12320 16856 0 _115_
rlabel metal2 12488 18928 12488 18928 0 _116_
rlabel metal2 11424 18424 11424 18424 0 _117_
rlabel metal3 19712 15848 19712 15848 0 _118_
rlabel metal2 17752 13216 17752 13216 0 _119_
rlabel metal2 19096 13720 19096 13720 0 _120_
rlabel metal2 18032 20216 18032 20216 0 _122_
rlabel metal2 17248 20776 17248 20776 0 _123_
rlabel metal2 16856 18928 16856 18928 0 _124_
rlabel metal2 17472 17640 17472 17640 0 _125_
rlabel metal2 14840 7182 14840 7182 0 clk
rlabel metal2 20216 15736 20216 15736 0 clknet_0_clk
rlabel metal2 14280 15232 14280 15232 0 clknet_1_0__leaf_clk
rlabel metal3 21784 13832 21784 13832 0 clknet_1_1__leaf_clk
rlabel metal3 25536 36456 25536 36456 0 in[0]
rlabel metal2 15736 3192 15736 3192 0 in[10]
rlabel metal2 23856 2184 23856 2184 0 in[11]
rlabel metal2 37576 3080 37576 3080 0 in[12]
rlabel metal3 38738 8120 38738 8120 0 in[13]
rlabel metal2 38248 9632 38248 9632 0 in[14]
rlabel metal2 38248 11816 38248 11816 0 in[15]
rlabel metal3 1246 12824 1246 12824 0 in[16]
rlabel metal3 1302 26264 1302 26264 0 in[17]
rlabel metal2 1848 25200 1848 25200 0 in[18]
rlabel metal2 14840 37842 14840 37842 0 in[1]
rlabel metal2 21672 36456 21672 36456 0 in[2]
rlabel metal2 16184 37562 16184 37562 0 in[3]
rlabel metal2 37576 36680 37576 36680 0 in[4]
rlabel metal2 38248 32424 38248 32424 0 in[5]
rlabel metal2 38304 36232 38304 36232 0 in[6]
rlabel metal2 38248 25928 38248 25928 0 in[7]
rlabel metal2 26264 3584 26264 3584 0 in[8]
rlabel metal1 26208 2520 26208 2520 0 in[9]
rlabel metal3 24136 26488 24136 26488 0 net1
rlabel metal2 10584 20552 10584 20552 0 net10
rlabel metal3 34160 27832 34160 27832 0 net100
rlabel metal2 27496 4256 27496 4256 0 net101
rlabel metal2 25592 8680 25592 8680 0 net102
rlabel metal2 2520 22736 2520 22736 0 net103
rlabel metal2 2744 21616 2744 21616 0 net104
rlabel metal2 2072 19320 2072 19320 0 net105
rlabel metal2 17304 8232 17304 8232 0 net106
rlabel metal2 19824 13944 19824 13944 0 net107
rlabel metal2 17976 13104 17976 13104 0 net108
rlabel metal2 15064 30128 15064 30128 0 net11
rlabel metal2 22176 31920 22176 31920 0 net12
rlabel metal2 16912 24024 16912 24024 0 net13
rlabel metal2 39200 35224 39200 35224 0 net14
rlabel metal2 38472 31920 38472 31920 0 net15
rlabel metal2 37408 34888 37408 34888 0 net16
rlabel metal2 26264 23128 26264 23128 0 net17
rlabel metal2 22008 17808 22008 17808 0 net18
rlabel metal3 23408 17528 23408 17528 0 net19
rlabel metal3 25088 16184 25088 16184 0 net2
rlabel metal2 15064 17864 15064 17864 0 net20
rlabel metal2 2128 13944 2128 13944 0 net21
rlabel metal2 14952 14336 14952 14336 0 net22
rlabel metal3 19432 15960 19432 15960 0 net23
rlabel metal2 19320 8680 19320 8680 0 net24
rlabel metal2 16632 8512 16632 8512 0 net25
rlabel metal2 16072 8904 16072 8904 0 net26
rlabel metal3 19656 30072 19656 30072 0 net27
rlabel metal2 25480 13552 25480 13552 0 net28
rlabel metal2 37240 13720 37240 13720 0 net29
rlabel metal2 21336 16240 21336 16240 0 net3
rlabel metal3 34944 16072 34944 16072 0 net30
rlabel metal3 34496 12824 34496 12824 0 net31
rlabel metal2 37352 10024 37352 10024 0 net32
rlabel metal3 37912 14336 37912 14336 0 net33
rlabel metal2 11872 19096 11872 19096 0 net34
rlabel metal2 2184 22232 2184 22232 0 net35
rlabel metal3 8400 21616 8400 21616 0 net36
rlabel metal2 23464 30856 23464 30856 0 net37
rlabel metal3 16688 28616 16688 28616 0 net38
rlabel metal3 24472 36344 24472 36344 0 net39
rlabel metal2 37184 3416 37184 3416 0 net4
rlabel metal2 22792 30856 22792 30856 0 net40
rlabel metal2 24416 35448 24416 35448 0 net41
rlabel metal2 30296 21896 30296 21896 0 net42
rlabel metal3 33152 20664 33152 20664 0 net43
rlabel metal2 36568 34132 36568 34132 0 net44
rlabel metal2 37968 27272 37968 27272 0 net45
rlabel metal2 21896 19152 21896 19152 0 net46
rlabel metal3 20776 17528 20776 17528 0 net47
rlabel metal2 19712 16296 19712 16296 0 net48
rlabel metal2 19488 33992 19488 33992 0 net49
rlabel metal2 37912 8260 37912 8260 0 net5
rlabel metal2 22344 16044 22344 16044 0 net50
rlabel metal3 33432 20104 33432 20104 0 net51
rlabel metal2 28280 20048 28280 20048 0 net52
rlabel metal2 37744 6552 37744 6552 0 net53
rlabel metal2 37912 7392 37912 7392 0 net54
rlabel metal2 14952 19152 14952 19152 0 net55
rlabel metal2 15512 21784 15512 21784 0 net56
rlabel metal2 14728 22008 14728 22008 0 net57
rlabel metal2 23576 20776 23576 20776 0 net58
rlabel metal2 23240 22904 23240 22904 0 net59
rlabel metal2 37912 10024 37912 10024 0 net6
rlabel metal2 17584 34104 17584 34104 0 net60
rlabel metal2 37912 28504 37912 28504 0 net61
rlabel metal2 37688 29288 37688 29288 0 net62
rlabel metal2 37912 21056 37912 21056 0 net63
rlabel metal2 24472 20832 24472 20832 0 net64
rlabel metal2 26152 22456 26152 22456 0 net65
rlabel metal2 27776 27160 27776 27160 0 net66
rlabel metal2 37912 4256 37912 4256 0 net67
rlabel metal2 24472 18368 24472 18368 0 net68
rlabel metal2 37240 8064 37240 8064 0 net69
rlabel metal2 37856 12376 37856 12376 0 net7
rlabel metal2 24752 17080 24752 17080 0 net70
rlabel metal3 33264 33208 33264 33208 0 net71
rlabel metal3 37184 3416 37184 3416 0 net72
rlabel metal2 30464 20104 30464 20104 0 net73
rlabel metal2 31304 6748 31304 6748 0 net74
rlabel metal2 37912 5824 37912 5824 0 net75
rlabel metal2 12600 17136 12600 17136 0 net76
rlabel metal2 15680 18984 15680 18984 0 net77
rlabel metal2 14952 17920 14952 17920 0 net78
rlabel metal2 21056 31920 21056 31920 0 net79
rlabel metal2 2184 12824 2184 12824 0 net8
rlabel metal2 17416 31920 17416 31920 0 net80
rlabel metal2 19208 31612 19208 31612 0 net81
rlabel metal2 38024 33712 38024 33712 0 net82
rlabel metal2 17808 21784 17808 21784 0 net83
rlabel metal2 38080 35672 38080 35672 0 net84
rlabel metal2 37240 31584 37240 31584 0 net85
rlabel metal2 37912 31836 37912 31836 0 net86
rlabel metal2 37912 30912 37912 30912 0 net87
rlabel metal2 21952 3528 21952 3528 0 net88
rlabel metal2 21504 3528 21504 3528 0 net89
rlabel metal2 12152 20048 12152 20048 0 net9
rlabel metal2 18928 16184 18928 16184 0 net90
rlabel metal2 22792 7672 22792 7672 0 net91
rlabel metal3 32928 10584 32928 10584 0 net92
rlabel metal2 37520 34776 37520 34776 0 net93
rlabel metal3 33040 13720 33040 13720 0 net94
rlabel metal2 26600 16520 26600 16520 0 net95
rlabel metal3 37464 14504 37464 14504 0 net96
rlabel metal2 12152 16128 12152 16128 0 net97
rlabel metal2 12600 18424 12600 18424 0 net98
rlabel metal2 10920 18088 10920 18088 0 net99
rlabel metal2 18872 2030 18872 2030 0 proj_clk[0]
rlabel metal2 19544 2030 19544 2030 0 proj_clk[1]
rlabel metal2 16296 4424 16296 4424 0 proj_clk[2]
rlabel metal2 16856 2058 16856 2058 0 proj_clk[3]
rlabel metal2 20216 37786 20216 37786 0 proj_in[0]
rlabel metal2 38304 11144 38304 11144 0 proj_in[10]
rlabel metal2 37576 12488 37576 12488 0 proj_in[11]
rlabel metal2 38304 15848 38304 15848 0 proj_in[12]
rlabel metal3 38738 12824 38738 12824 0 proj_in[13]
rlabel metal2 38248 8960 38248 8960 0 proj_in[14]
rlabel metal3 38584 14280 38584 14280 0 proj_in[15]
rlabel metal3 1246 20216 1246 20216 0 proj_in[16]
rlabel metal3 1246 23576 1246 23576 0 proj_in[17]
rlabel metal3 1246 20888 1246 20888 0 proj_in[18]
rlabel metal2 23016 36344 23016 36344 0 proj_in[19]
rlabel metal2 15512 36344 15512 36344 0 proj_in[1]
rlabel metal2 25256 36512 25256 36512 0 proj_in[20]
rlabel metal2 22344 36344 22344 36344 0 proj_in[21]
rlabel metal2 24584 36400 24584 36400 0 proj_in[22]
rlabel metal3 38738 22232 38738 22232 0 proj_in[23]
rlabel metal2 38192 26936 38192 26936 0 proj_in[24]
rlabel metal3 38066 36344 38066 36344 0 proj_in[25]
rlabel metal2 38248 29232 38248 29232 0 proj_in[26]
rlabel metal3 38584 18984 38584 18984 0 proj_in[27]
rlabel metal3 38738 17528 38738 17528 0 proj_in[28]
rlabel metal2 20216 2030 20216 2030 0 proj_in[29]
rlabel metal2 18872 37786 18872 37786 0 proj_in[2]
rlabel metal2 22904 2030 22904 2030 0 proj_in[30]
rlabel metal2 38248 19824 38248 19824 0 proj_in[31]
rlabel metal2 38304 20552 38304 20552 0 proj_in[32]
rlabel metal2 38248 6328 38248 6328 0 proj_in[33]
rlabel metal2 38248 7168 38248 7168 0 proj_in[34]
rlabel metal3 1246 25592 1246 25592 0 proj_in[35]
rlabel metal3 1246 22904 1246 22904 0 proj_in[36]
rlabel metal3 1246 22232 1246 22232 0 proj_in[37]
rlabel metal2 37576 21840 37576 21840 0 proj_in[38]
rlabel metal3 38584 23688 38584 23688 0 proj_in[39]
rlabel metal2 17528 37786 17528 37786 0 proj_in[3]
rlabel metal3 38584 28392 38584 28392 0 proj_in[40]
rlabel metal2 38248 29848 38248 29848 0 proj_in[41]
rlabel metal2 38248 21280 38248 21280 0 proj_in[42]
rlabel metal2 38248 25144 38248 25144 0 proj_in[43]
rlabel metal2 38248 23072 38248 23072 0 proj_in[44]
rlabel metal2 37576 26992 37576 26992 0 proj_in[45]
rlabel metal2 38248 4256 38248 4256 0 proj_in[46]
rlabel metal2 38248 18368 38248 18368 0 proj_in[47]
rlabel metal2 37576 7728 37576 7728 0 proj_in[48]
rlabel metal2 37576 17136 37576 17136 0 proj_in[49]
rlabel metal3 38584 33096 38584 33096 0 proj_in[4]
rlabel metal3 38738 3416 38738 3416 0 proj_in[50]
rlabel metal2 38248 24528 38248 24528 0 proj_in[51]
rlabel metal3 38584 4872 38584 4872 0 proj_in[52]
rlabel metal2 38248 5712 38248 5712 0 proj_in[53]
rlabel metal3 1246 16184 1246 16184 0 proj_in[54]
rlabel metal3 1246 19544 1246 19544 0 proj_in[55]
rlabel metal3 1246 18200 1246 18200 0 proj_in[56]
rlabel metal2 21000 36344 21000 36344 0 proj_in[57]
rlabel metal2 16408 36624 16408 36624 0 proj_in[58]
rlabel metal2 19544 37786 19544 37786 0 proj_in[59]
rlabel metal2 38248 33936 38248 33936 0 proj_in[5]
rlabel metal2 18200 37786 18200 37786 0 proj_in[60]
rlabel metal2 38248 35392 38248 35392 0 proj_in[61]
rlabel metal3 38402 31640 38402 31640 0 proj_in[62]
rlabel metal2 38304 31528 38304 31528 0 proj_in[63]
rlabel metal2 38248 30688 38248 30688 0 proj_in[64]
rlabel metal2 21560 2030 21560 2030 0 proj_in[65]
rlabel metal2 20888 2030 20888 2030 0 proj_in[66]
rlabel metal2 18200 2030 18200 2030 0 proj_in[67]
rlabel metal2 22232 2030 22232 2030 0 proj_in[68]
rlabel metal2 38248 10416 38248 10416 0 proj_in[69]
rlabel metal2 38304 34664 38304 34664 0 proj_in[6]
rlabel metal2 38248 13664 38248 13664 0 proj_in[70]
rlabel metal2 38248 16576 38248 16576 0 proj_in[71]
rlabel metal3 38738 14840 38738 14840 0 proj_in[72]
rlabel metal3 1246 14840 1246 14840 0 proj_in[73]
rlabel metal3 1246 15512 1246 15512 0 proj_in[74]
rlabel metal3 1022 16856 1022 16856 0 proj_in[75]
rlabel metal2 38248 27776 38248 27776 0 proj_in[7]
rlabel metal2 26264 2058 26264 2058 0 proj_in[8]
rlabel metal3 24752 3416 24752 3416 0 proj_in[9]
rlabel metal3 1246 24248 1246 24248 0 proj_rst_n[0]
rlabel metal3 854 21560 854 21560 0 proj_rst_n[1]
rlabel metal3 1246 18872 1246 18872 0 proj_rst_n[2]
rlabel metal2 17528 2030 17528 2030 0 proj_rst_n[3]
rlabel metal3 1246 17528 1246 17528 0 rst_n
rlabel metal2 1736 13608 1736 13608 0 sel[0]
rlabel metal2 1736 14280 1736 14280 0 sel[1]
rlabel metal3 17584 14728 17584 14728 0 sel_latched\[0\]
rlabel metal2 18088 14448 18088 14448 0 sel_latched\[1\]
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
