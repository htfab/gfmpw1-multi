VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rotfpga2a
  CLASS BLOCK ;
  FOREIGN rotfpga2a ;
  ORIGIN 0.000 0.000 ;
  SIZE 320.000 BY 320.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.560 4.000 ;
    END
  END clk
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 272.160 4.000 272.720 ;
    END
  END in[0]
  PIN in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 147.840 320.000 148.400 ;
    END
  END in[10]
  PIN in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 151.200 320.000 151.760 ;
    END
  END in[11]
  PIN in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END in[12]
  PIN in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END in[13]
  PIN in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 144.480 320.000 145.040 ;
    END
  END in[14]
  PIN in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 137.760 320.000 138.320 ;
    END
  END in[15]
  PIN in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 141.120 320.000 141.680 ;
    END
  END in[16]
  PIN in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 4.000 ;
    END
  END in[17]
  PIN in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 0.000 7.280 4.000 ;
    END
  END in[18]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 4.000 ;
    END
  END in[1]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 164.640 320.000 165.200 ;
    END
  END in[2]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 0.000 148.400 4.000 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 4.000 57.680 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END in[7]
  PIN in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.760 4.000 222.320 ;
    END
  END in[8]
  PIN in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 316.000 148.400 320.000 ;
    END
  END in[9]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 215.040 320.000 215.600 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 292.320 320.000 292.880 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 316.000 192.080 320.000 ;
    END
  END out[11]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 316.000 154.560 320.000 155.120 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 4.000 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 316.000 81.200 320.000 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 316.000 131.600 320.000 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 316.000 242.480 320.000 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 316.000 239.120 320.000 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 4.000 ;
    END
  END out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 4.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 302.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 302.140 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 302.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 302.140 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 313.040 302.140 ;
      LAYER Metal2 ;
        RECT 4.620 315.700 80.340 316.000 ;
        RECT 81.500 315.700 130.740 316.000 ;
        RECT 131.900 315.700 147.540 316.000 ;
        RECT 148.700 315.700 191.220 316.000 ;
        RECT 192.380 315.700 238.260 316.000 ;
        RECT 239.420 315.700 241.620 316.000 ;
        RECT 242.780 315.700 315.140 316.000 ;
        RECT 4.620 4.300 315.140 315.700 ;
        RECT 4.620 3.500 6.420 4.300 ;
        RECT 7.580 3.500 9.780 4.300 ;
        RECT 10.940 3.500 36.660 4.300 ;
        RECT 37.820 3.500 147.540 4.300 ;
        RECT 148.700 3.500 157.620 4.300 ;
        RECT 158.780 3.500 160.980 4.300 ;
        RECT 162.140 3.500 164.340 4.300 ;
        RECT 165.500 3.500 171.060 4.300 ;
        RECT 172.220 3.500 191.220 4.300 ;
        RECT 192.380 3.500 315.140 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 293.180 316.000 302.820 ;
        RECT 4.000 292.020 315.700 293.180 ;
        RECT 4.000 273.020 316.000 292.020 ;
        RECT 4.300 271.860 316.000 273.020 ;
        RECT 4.000 222.620 316.000 271.860 ;
        RECT 4.300 221.460 316.000 222.620 ;
        RECT 4.000 215.900 316.000 221.460 ;
        RECT 4.000 214.740 315.700 215.900 ;
        RECT 4.000 168.860 316.000 214.740 ;
        RECT 4.300 167.700 316.000 168.860 ;
        RECT 4.000 165.500 316.000 167.700 ;
        RECT 4.000 164.340 315.700 165.500 ;
        RECT 4.000 155.420 316.000 164.340 ;
        RECT 4.300 154.260 315.700 155.420 ;
        RECT 4.000 152.060 316.000 154.260 ;
        RECT 4.000 150.900 315.700 152.060 ;
        RECT 4.000 148.700 316.000 150.900 ;
        RECT 4.000 147.540 315.700 148.700 ;
        RECT 4.000 145.340 316.000 147.540 ;
        RECT 4.000 144.180 315.700 145.340 ;
        RECT 4.000 141.980 316.000 144.180 ;
        RECT 4.000 140.820 315.700 141.980 ;
        RECT 4.000 138.620 316.000 140.820 ;
        RECT 4.000 137.460 315.700 138.620 ;
        RECT 4.000 125.180 316.000 137.460 ;
        RECT 4.300 124.020 316.000 125.180 ;
        RECT 4.000 121.820 316.000 124.020 ;
        RECT 4.300 120.660 316.000 121.820 ;
        RECT 4.000 57.980 316.000 120.660 ;
        RECT 4.300 56.820 316.000 57.980 ;
        RECT 4.000 14.700 316.000 56.820 ;
      LAYER Metal4 ;
        RECT 8.540 15.080 21.940 292.790 ;
        RECT 24.140 15.080 98.740 292.790 ;
        RECT 100.940 15.080 175.540 292.790 ;
        RECT 177.740 15.080 252.340 292.790 ;
        RECT 254.540 15.080 311.220 292.790 ;
        RECT 8.540 14.650 311.220 15.080 ;
  END
END rotfpga2a
END LIBRARY

