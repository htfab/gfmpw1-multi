magic
tech gf180mcuD
magscale 1 5
timestamp 1702353081
<< metal1 >>
rect 672 18437 19320 18454
rect 672 18411 2938 18437
rect 2964 18411 2990 18437
rect 3016 18411 3042 18437
rect 3068 18411 7600 18437
rect 7626 18411 7652 18437
rect 7678 18411 7704 18437
rect 7730 18411 12262 18437
rect 12288 18411 12314 18437
rect 12340 18411 12366 18437
rect 12392 18411 16924 18437
rect 16950 18411 16976 18437
rect 17002 18411 17028 18437
rect 17054 18411 19320 18437
rect 672 18394 19320 18411
rect 9031 18353 9057 18359
rect 9031 18321 9057 18327
rect 10151 18297 10177 18303
rect 7401 18271 7407 18297
rect 7433 18271 7439 18297
rect 10151 18265 10177 18271
rect 10879 18241 10905 18247
rect 8185 18215 8191 18241
rect 8217 18215 8223 18241
rect 8633 18215 8639 18241
rect 8665 18215 8671 18241
rect 10649 18215 10655 18241
rect 10681 18215 10687 18241
rect 11321 18215 11327 18241
rect 11353 18215 11359 18241
rect 10879 18209 10905 18215
rect 10543 18129 10569 18135
rect 10543 18097 10569 18103
rect 11047 18129 11073 18135
rect 11047 18097 11073 18103
rect 11215 18129 11241 18135
rect 11215 18097 11241 18103
rect 672 18045 19400 18062
rect 672 18019 5269 18045
rect 5295 18019 5321 18045
rect 5347 18019 5373 18045
rect 5399 18019 9931 18045
rect 9957 18019 9983 18045
rect 10009 18019 10035 18045
rect 10061 18019 14593 18045
rect 14619 18019 14645 18045
rect 14671 18019 14697 18045
rect 14723 18019 19255 18045
rect 19281 18019 19307 18045
rect 19333 18019 19359 18045
rect 19385 18019 19400 18045
rect 672 18002 19400 18019
rect 7519 17961 7545 17967
rect 7519 17929 7545 17935
rect 9871 17961 9897 17967
rect 9871 17929 9897 17935
rect 10767 17961 10793 17967
rect 10767 17929 10793 17935
rect 11103 17961 11129 17967
rect 11103 17929 11129 17935
rect 7855 17905 7881 17911
rect 7855 17873 7881 17879
rect 8023 17905 8049 17911
rect 8023 17873 8049 17879
rect 8191 17905 8217 17911
rect 8191 17873 8217 17879
rect 8359 17905 8385 17911
rect 8359 17873 8385 17879
rect 8863 17905 8889 17911
rect 8863 17873 8889 17879
rect 9031 17905 9057 17911
rect 9031 17873 9057 17879
rect 9199 17905 9225 17911
rect 9199 17873 9225 17879
rect 9535 17905 9561 17911
rect 9535 17873 9561 17879
rect 10207 17905 10233 17911
rect 10207 17873 10233 17879
rect 10375 17905 10401 17911
rect 10375 17873 10401 17879
rect 9305 17823 9311 17849
rect 9337 17823 9343 17849
rect 9641 17823 9647 17849
rect 9673 17823 9679 17849
rect 9977 17823 9983 17849
rect 10009 17823 10015 17849
rect 7743 17793 7769 17799
rect 7743 17761 7769 17767
rect 672 17653 19320 17670
rect 672 17627 2938 17653
rect 2964 17627 2990 17653
rect 3016 17627 3042 17653
rect 3068 17627 7600 17653
rect 7626 17627 7652 17653
rect 7678 17627 7704 17653
rect 7730 17627 12262 17653
rect 12288 17627 12314 17653
rect 12340 17627 12366 17653
rect 12392 17627 16924 17653
rect 16950 17627 16976 17653
rect 17002 17627 17028 17653
rect 17054 17627 19320 17653
rect 672 17610 19320 17627
rect 8751 17513 8777 17519
rect 8751 17481 8777 17487
rect 9087 17513 9113 17519
rect 9087 17481 9113 17487
rect 9423 17513 9449 17519
rect 9423 17481 9449 17487
rect 9759 17513 9785 17519
rect 9759 17481 9785 17487
rect 10095 17513 10121 17519
rect 10095 17481 10121 17487
rect 672 17261 19400 17278
rect 672 17235 5269 17261
rect 5295 17235 5321 17261
rect 5347 17235 5373 17261
rect 5399 17235 9931 17261
rect 9957 17235 9983 17261
rect 10009 17235 10035 17261
rect 10061 17235 14593 17261
rect 14619 17235 14645 17261
rect 14671 17235 14697 17261
rect 14723 17235 19255 17261
rect 19281 17235 19307 17261
rect 19333 17235 19359 17261
rect 19385 17235 19400 17261
rect 672 17218 19400 17235
rect 672 16869 19320 16886
rect 672 16843 2938 16869
rect 2964 16843 2990 16869
rect 3016 16843 3042 16869
rect 3068 16843 7600 16869
rect 7626 16843 7652 16869
rect 7678 16843 7704 16869
rect 7730 16843 12262 16869
rect 12288 16843 12314 16869
rect 12340 16843 12366 16869
rect 12392 16843 16924 16869
rect 16950 16843 16976 16869
rect 17002 16843 17028 16869
rect 17054 16843 19320 16869
rect 672 16826 19320 16843
rect 672 16477 19400 16494
rect 672 16451 5269 16477
rect 5295 16451 5321 16477
rect 5347 16451 5373 16477
rect 5399 16451 9931 16477
rect 9957 16451 9983 16477
rect 10009 16451 10035 16477
rect 10061 16451 14593 16477
rect 14619 16451 14645 16477
rect 14671 16451 14697 16477
rect 14723 16451 19255 16477
rect 19281 16451 19307 16477
rect 19333 16451 19359 16477
rect 19385 16451 19400 16477
rect 672 16434 19400 16451
rect 672 16085 19320 16102
rect 672 16059 2938 16085
rect 2964 16059 2990 16085
rect 3016 16059 3042 16085
rect 3068 16059 7600 16085
rect 7626 16059 7652 16085
rect 7678 16059 7704 16085
rect 7730 16059 12262 16085
rect 12288 16059 12314 16085
rect 12340 16059 12366 16085
rect 12392 16059 16924 16085
rect 16950 16059 16976 16085
rect 17002 16059 17028 16085
rect 17054 16059 19320 16085
rect 672 16042 19320 16059
rect 672 15693 19400 15710
rect 672 15667 5269 15693
rect 5295 15667 5321 15693
rect 5347 15667 5373 15693
rect 5399 15667 9931 15693
rect 9957 15667 9983 15693
rect 10009 15667 10035 15693
rect 10061 15667 14593 15693
rect 14619 15667 14645 15693
rect 14671 15667 14697 15693
rect 14723 15667 19255 15693
rect 19281 15667 19307 15693
rect 19333 15667 19359 15693
rect 19385 15667 19400 15693
rect 672 15650 19400 15667
rect 672 15301 19320 15318
rect 672 15275 2938 15301
rect 2964 15275 2990 15301
rect 3016 15275 3042 15301
rect 3068 15275 7600 15301
rect 7626 15275 7652 15301
rect 7678 15275 7704 15301
rect 7730 15275 12262 15301
rect 12288 15275 12314 15301
rect 12340 15275 12366 15301
rect 12392 15275 16924 15301
rect 16950 15275 16976 15301
rect 17002 15275 17028 15301
rect 17054 15275 19320 15301
rect 672 15258 19320 15275
rect 672 14909 19400 14926
rect 672 14883 5269 14909
rect 5295 14883 5321 14909
rect 5347 14883 5373 14909
rect 5399 14883 9931 14909
rect 9957 14883 9983 14909
rect 10009 14883 10035 14909
rect 10061 14883 14593 14909
rect 14619 14883 14645 14909
rect 14671 14883 14697 14909
rect 14723 14883 19255 14909
rect 19281 14883 19307 14909
rect 19333 14883 19359 14909
rect 19385 14883 19400 14909
rect 672 14866 19400 14883
rect 672 14517 19320 14534
rect 672 14491 2938 14517
rect 2964 14491 2990 14517
rect 3016 14491 3042 14517
rect 3068 14491 7600 14517
rect 7626 14491 7652 14517
rect 7678 14491 7704 14517
rect 7730 14491 12262 14517
rect 12288 14491 12314 14517
rect 12340 14491 12366 14517
rect 12392 14491 16924 14517
rect 16950 14491 16976 14517
rect 17002 14491 17028 14517
rect 17054 14491 19320 14517
rect 672 14474 19320 14491
rect 672 14125 19400 14142
rect 672 14099 5269 14125
rect 5295 14099 5321 14125
rect 5347 14099 5373 14125
rect 5399 14099 9931 14125
rect 9957 14099 9983 14125
rect 10009 14099 10035 14125
rect 10061 14099 14593 14125
rect 14619 14099 14645 14125
rect 14671 14099 14697 14125
rect 14723 14099 19255 14125
rect 19281 14099 19307 14125
rect 19333 14099 19359 14125
rect 19385 14099 19400 14125
rect 672 14082 19400 14099
rect 672 13733 19320 13750
rect 672 13707 2938 13733
rect 2964 13707 2990 13733
rect 3016 13707 3042 13733
rect 3068 13707 7600 13733
rect 7626 13707 7652 13733
rect 7678 13707 7704 13733
rect 7730 13707 12262 13733
rect 12288 13707 12314 13733
rect 12340 13707 12366 13733
rect 12392 13707 16924 13733
rect 16950 13707 16976 13733
rect 17002 13707 17028 13733
rect 17054 13707 19320 13733
rect 672 13690 19320 13707
rect 672 13341 19400 13358
rect 672 13315 5269 13341
rect 5295 13315 5321 13341
rect 5347 13315 5373 13341
rect 5399 13315 9931 13341
rect 9957 13315 9983 13341
rect 10009 13315 10035 13341
rect 10061 13315 14593 13341
rect 14619 13315 14645 13341
rect 14671 13315 14697 13341
rect 14723 13315 19255 13341
rect 19281 13315 19307 13341
rect 19333 13315 19359 13341
rect 19385 13315 19400 13341
rect 672 13298 19400 13315
rect 2137 13119 2143 13145
rect 2169 13119 2175 13145
rect 2423 13089 2449 13095
rect 2423 13057 2449 13063
rect 967 13033 993 13039
rect 967 13001 993 13007
rect 672 12949 19320 12966
rect 672 12923 2938 12949
rect 2964 12923 2990 12949
rect 3016 12923 3042 12949
rect 3068 12923 7600 12949
rect 7626 12923 7652 12949
rect 7678 12923 7704 12949
rect 7730 12923 12262 12949
rect 12288 12923 12314 12949
rect 12340 12923 12366 12949
rect 12392 12923 16924 12949
rect 16950 12923 16976 12949
rect 17002 12923 17028 12949
rect 17054 12923 19320 12949
rect 672 12906 19320 12923
rect 855 12697 881 12703
rect 855 12665 881 12671
rect 1023 12641 1049 12647
rect 1023 12609 1049 12615
rect 1247 12641 1273 12647
rect 1247 12609 1273 12615
rect 672 12557 19400 12574
rect 672 12531 5269 12557
rect 5295 12531 5321 12557
rect 5347 12531 5373 12557
rect 5399 12531 9931 12557
rect 9957 12531 9983 12557
rect 10009 12531 10035 12557
rect 10061 12531 14593 12557
rect 14619 12531 14645 12557
rect 14671 12531 14697 12557
rect 14723 12531 19255 12557
rect 19281 12531 19307 12557
rect 19333 12531 19359 12557
rect 19385 12531 19400 12557
rect 672 12514 19400 12531
rect 8689 12447 8695 12473
rect 8721 12447 8727 12473
rect 1023 12417 1049 12423
rect 1023 12385 1049 12391
rect 855 12361 881 12367
rect 8801 12335 8807 12361
rect 8833 12335 8839 12361
rect 17817 12335 17823 12361
rect 17849 12335 17855 12361
rect 855 12329 881 12335
rect 1247 12305 1273 12311
rect 1247 12273 1273 12279
rect 18999 12249 19025 12255
rect 18999 12217 19025 12223
rect 672 12165 19320 12182
rect 672 12139 2938 12165
rect 2964 12139 2990 12165
rect 3016 12139 3042 12165
rect 3068 12139 7600 12165
rect 7626 12139 7652 12165
rect 7678 12139 7704 12165
rect 7730 12139 12262 12165
rect 12288 12139 12314 12165
rect 12340 12139 12366 12165
rect 12392 12139 16924 12165
rect 16950 12139 16976 12165
rect 17002 12139 17028 12165
rect 17054 12139 19320 12165
rect 672 12122 19320 12139
rect 8023 12025 8049 12031
rect 8023 11993 8049 11999
rect 8863 11969 8889 11975
rect 8185 11943 8191 11969
rect 8217 11943 8223 11969
rect 8409 11943 8415 11969
rect 8441 11943 8447 11969
rect 9081 11943 9087 11969
rect 9113 11943 9119 11969
rect 9529 11943 9535 11969
rect 9561 11943 9567 11969
rect 8863 11937 8889 11943
rect 855 11913 881 11919
rect 855 11881 881 11887
rect 19111 11913 19137 11919
rect 19111 11881 19137 11887
rect 1023 11857 1049 11863
rect 1023 11825 1049 11831
rect 1247 11857 1273 11863
rect 18831 11857 18857 11863
rect 8521 11831 8527 11857
rect 8553 11831 8559 11857
rect 1247 11825 1273 11831
rect 18831 11825 18857 11831
rect 18943 11857 18969 11863
rect 18943 11825 18969 11831
rect 672 11773 19400 11790
rect 672 11747 5269 11773
rect 5295 11747 5321 11773
rect 5347 11747 5373 11773
rect 5399 11747 9931 11773
rect 9957 11747 9983 11773
rect 10009 11747 10035 11773
rect 10061 11747 14593 11773
rect 14619 11747 14645 11773
rect 14671 11747 14697 11773
rect 14723 11747 19255 11773
rect 19281 11747 19307 11773
rect 19333 11747 19359 11773
rect 19385 11747 19400 11773
rect 672 11730 19400 11747
rect 1023 11633 1049 11639
rect 18943 11633 18969 11639
rect 8689 11607 8695 11633
rect 8721 11607 8727 11633
rect 1023 11601 1049 11607
rect 18943 11601 18969 11607
rect 855 11577 881 11583
rect 19111 11577 19137 11583
rect 8801 11551 8807 11577
rect 8833 11551 8839 11577
rect 855 11545 881 11551
rect 19111 11545 19137 11551
rect 1247 11521 1273 11527
rect 1247 11489 1273 11495
rect 18831 11521 18857 11527
rect 18831 11489 18857 11495
rect 672 11381 19320 11398
rect 672 11355 2938 11381
rect 2964 11355 2990 11381
rect 3016 11355 3042 11381
rect 3068 11355 7600 11381
rect 7626 11355 7652 11381
rect 7678 11355 7704 11381
rect 7730 11355 12262 11381
rect 12288 11355 12314 11381
rect 12340 11355 12366 11381
rect 12392 11355 16924 11381
rect 16950 11355 16976 11381
rect 17002 11355 17028 11381
rect 17054 11355 19320 11381
rect 672 11338 19320 11355
rect 8023 11241 8049 11247
rect 8023 11209 8049 11215
rect 8863 11185 8889 11191
rect 8185 11159 8191 11185
rect 8217 11159 8223 11185
rect 8409 11159 8415 11185
rect 8441 11159 8447 11185
rect 9137 11159 9143 11185
rect 9169 11159 9175 11185
rect 9585 11159 9591 11185
rect 9617 11159 9623 11185
rect 8863 11153 8889 11159
rect 855 11129 881 11135
rect 855 11097 881 11103
rect 1023 11129 1049 11135
rect 1023 11097 1049 11103
rect 1191 11129 1217 11135
rect 18831 11129 18857 11135
rect 8521 11103 8527 11129
rect 8553 11103 8559 11129
rect 11209 11103 11215 11129
rect 11241 11103 11247 11129
rect 1191 11097 1217 11103
rect 18831 11097 18857 11103
rect 19111 11129 19137 11135
rect 19111 11097 19137 11103
rect 1359 11073 1385 11079
rect 1359 11041 1385 11047
rect 1583 11073 1609 11079
rect 1583 11041 1609 11047
rect 10711 11073 10737 11079
rect 11047 11073 11073 11079
rect 10873 11047 10879 11073
rect 10905 11047 10911 11073
rect 10711 11041 10737 11047
rect 11047 11041 11073 11047
rect 18943 11073 18969 11079
rect 18943 11041 18969 11047
rect 672 10989 19400 11006
rect 672 10963 5269 10989
rect 5295 10963 5321 10989
rect 5347 10963 5373 10989
rect 5399 10963 9931 10989
rect 9957 10963 9983 10989
rect 10009 10963 10035 10989
rect 10061 10963 14593 10989
rect 14619 10963 14645 10989
rect 14671 10963 14697 10989
rect 14723 10963 19255 10989
rect 19281 10963 19307 10989
rect 19333 10963 19359 10989
rect 19385 10963 19400 10989
rect 672 10946 19400 10963
rect 1247 10905 1273 10911
rect 10985 10879 10991 10905
rect 11017 10879 11023 10905
rect 1247 10873 1273 10879
rect 1023 10849 1049 10855
rect 1023 10817 1049 10823
rect 10487 10849 10513 10855
rect 10487 10817 10513 10823
rect 855 10793 881 10799
rect 11327 10793 11353 10799
rect 10705 10767 10711 10793
rect 10737 10767 10743 10793
rect 10929 10767 10935 10793
rect 10961 10767 10967 10793
rect 11601 10767 11607 10793
rect 11633 10767 11639 10793
rect 12049 10767 12055 10793
rect 12081 10767 12087 10793
rect 17817 10767 17823 10793
rect 17849 10767 17855 10793
rect 855 10761 881 10767
rect 11327 10761 11353 10767
rect 1471 10737 1497 10743
rect 1471 10705 1497 10711
rect 18999 10737 19025 10743
rect 18999 10705 19025 10711
rect 672 10597 19320 10614
rect 672 10571 2938 10597
rect 2964 10571 2990 10597
rect 3016 10571 3042 10597
rect 3068 10571 7600 10597
rect 7626 10571 7652 10597
rect 7678 10571 7704 10597
rect 7730 10571 12262 10597
rect 12288 10571 12314 10597
rect 12340 10571 12366 10597
rect 12392 10571 16924 10597
rect 16950 10571 16976 10597
rect 17002 10571 17028 10597
rect 17054 10571 19320 10597
rect 672 10554 19320 10571
rect 7855 10457 7881 10463
rect 7855 10425 7881 10431
rect 10655 10457 10681 10463
rect 10655 10425 10681 10431
rect 18271 10457 18297 10463
rect 18271 10425 18297 10431
rect 8695 10401 8721 10407
rect 11383 10401 11409 10407
rect 19111 10401 19137 10407
rect 8073 10375 8079 10401
rect 8105 10375 8111 10401
rect 8241 10375 8247 10401
rect 8273 10375 8279 10401
rect 8857 10375 8863 10401
rect 8889 10375 8895 10401
rect 9417 10375 9423 10401
rect 9449 10375 9455 10401
rect 10817 10375 10823 10401
rect 10849 10375 10855 10401
rect 11041 10375 11047 10401
rect 11073 10375 11079 10401
rect 11713 10375 11719 10401
rect 11745 10375 11751 10401
rect 12217 10375 12223 10401
rect 12249 10375 12255 10401
rect 8695 10369 8721 10375
rect 11383 10369 11409 10375
rect 19111 10369 19137 10375
rect 855 10345 881 10351
rect 855 10313 881 10319
rect 7743 10345 7769 10351
rect 18775 10345 18801 10351
rect 11153 10319 11159 10345
rect 11185 10319 11191 10345
rect 7743 10313 7769 10319
rect 18775 10313 18801 10319
rect 18943 10345 18969 10351
rect 18943 10313 18969 10319
rect 1023 10289 1049 10295
rect 1023 10257 1049 10263
rect 1247 10289 1273 10295
rect 18607 10289 18633 10295
rect 8353 10263 8359 10289
rect 8385 10263 8391 10289
rect 1247 10257 1273 10263
rect 18607 10257 18633 10263
rect 672 10205 19400 10222
rect 672 10179 5269 10205
rect 5295 10179 5321 10205
rect 5347 10179 5373 10205
rect 5399 10179 9931 10205
rect 9957 10179 9983 10205
rect 10009 10179 10035 10205
rect 10061 10179 14593 10205
rect 14619 10179 14645 10205
rect 14671 10179 14697 10205
rect 14723 10179 19255 10205
rect 19281 10179 19307 10205
rect 19333 10179 19359 10205
rect 19385 10179 19400 10205
rect 672 10162 19400 10179
rect 18831 10121 18857 10127
rect 18831 10089 18857 10095
rect 18943 10065 18969 10071
rect 8241 10039 8247 10065
rect 8273 10039 8279 10065
rect 8689 10039 8695 10065
rect 8721 10039 8727 10065
rect 18943 10033 18969 10039
rect 19111 10009 19137 10015
rect 2137 9983 2143 10009
rect 2169 9983 2175 10009
rect 8353 9983 8359 10009
rect 8385 9983 8391 10009
rect 8801 9983 8807 10009
rect 8833 9983 8839 10009
rect 19111 9977 19137 9983
rect 9535 9953 9561 9959
rect 9535 9921 9561 9927
rect 18607 9953 18633 9959
rect 18607 9921 18633 9927
rect 967 9897 993 9903
rect 967 9865 993 9871
rect 672 9813 19320 9830
rect 672 9787 2938 9813
rect 2964 9787 2990 9813
rect 3016 9787 3042 9813
rect 3068 9787 7600 9813
rect 7626 9787 7652 9813
rect 7678 9787 7704 9813
rect 7730 9787 12262 9813
rect 12288 9787 12314 9813
rect 12340 9787 12366 9813
rect 12392 9787 16924 9813
rect 16950 9787 16976 9813
rect 17002 9787 17028 9813
rect 17054 9787 19320 9813
rect 672 9770 19320 9787
rect 9927 9673 9953 9679
rect 9927 9641 9953 9647
rect 8695 9617 8721 9623
rect 8017 9591 8023 9617
rect 8049 9591 8055 9617
rect 8241 9591 8247 9617
rect 8273 9591 8279 9617
rect 8969 9591 8975 9617
rect 9001 9591 9007 9617
rect 9361 9591 9367 9617
rect 9393 9591 9399 9617
rect 8695 9585 8721 9591
rect 855 9561 881 9567
rect 855 9529 881 9535
rect 7743 9561 7769 9567
rect 7743 9529 7769 9535
rect 7855 9561 7881 9567
rect 18831 9561 18857 9567
rect 8353 9535 8359 9561
rect 8385 9535 8391 9561
rect 7855 9529 7881 9535
rect 18831 9529 18857 9535
rect 19111 9561 19137 9567
rect 19111 9529 19137 9535
rect 1023 9505 1049 9511
rect 1023 9473 1049 9479
rect 1247 9505 1273 9511
rect 1247 9473 1273 9479
rect 9647 9505 9673 9511
rect 9647 9473 9673 9479
rect 10095 9505 10121 9511
rect 11159 9505 11185 9511
rect 11495 9505 11521 9511
rect 18943 9505 18969 9511
rect 10257 9479 10263 9505
rect 10289 9479 10295 9505
rect 11321 9479 11327 9505
rect 11353 9479 11359 9505
rect 11657 9479 11663 9505
rect 11689 9479 11695 9505
rect 10095 9473 10121 9479
rect 11159 9473 11185 9479
rect 11495 9473 11521 9479
rect 18943 9473 18969 9479
rect 672 9421 19400 9438
rect 672 9395 5269 9421
rect 5295 9395 5321 9421
rect 5347 9395 5373 9421
rect 5399 9395 9931 9421
rect 9957 9395 9983 9421
rect 10009 9395 10035 9421
rect 10061 9395 14593 9421
rect 14619 9395 14645 9421
rect 14671 9395 14697 9421
rect 14723 9395 19255 9421
rect 19281 9395 19307 9421
rect 19333 9395 19359 9421
rect 19385 9395 19400 9421
rect 672 9378 19400 9395
rect 9137 9311 9143 9337
rect 9169 9311 9175 9337
rect 11097 9311 11103 9337
rect 11129 9311 11135 9337
rect 1023 9281 1049 9287
rect 1023 9249 1049 9255
rect 18943 9281 18969 9287
rect 18943 9249 18969 9255
rect 855 9225 881 9231
rect 855 9193 881 9199
rect 8695 9225 8721 9231
rect 9311 9225 9337 9231
rect 11327 9225 11353 9231
rect 19111 9225 19137 9231
rect 8913 9199 8919 9225
rect 8945 9199 8951 9225
rect 10817 9199 10823 9225
rect 10849 9199 10855 9225
rect 11041 9199 11047 9225
rect 11073 9199 11079 9225
rect 11713 9199 11719 9225
rect 11745 9199 11751 9225
rect 12161 9199 12167 9225
rect 12193 9199 12199 9225
rect 8695 9193 8721 9199
rect 9311 9193 9337 9199
rect 11327 9193 11353 9199
rect 19111 9193 19137 9199
rect 1247 9169 1273 9175
rect 1247 9137 1273 9143
rect 8415 9169 8441 9175
rect 8415 9137 8441 9143
rect 10599 9169 10625 9175
rect 10599 9137 10625 9143
rect 12671 9169 12697 9175
rect 12671 9137 12697 9143
rect 12951 9169 12977 9175
rect 12951 9137 12977 9143
rect 18831 9169 18857 9175
rect 18831 9137 18857 9143
rect 672 9029 19320 9046
rect 672 9003 2938 9029
rect 2964 9003 2990 9029
rect 3016 9003 3042 9029
rect 3068 9003 7600 9029
rect 7626 9003 7652 9029
rect 7678 9003 7704 9029
rect 7730 9003 12262 9029
rect 12288 9003 12314 9029
rect 12340 9003 12366 9029
rect 12392 9003 16924 9029
rect 16950 9003 16976 9029
rect 17002 9003 17028 9029
rect 17054 9003 19320 9029
rect 672 8986 19320 9003
rect 967 8889 993 8895
rect 8857 8863 8863 8889
rect 8889 8863 8895 8889
rect 967 8857 993 8863
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 9025 8807 9031 8833
rect 9057 8807 9063 8833
rect 9585 8807 9591 8833
rect 9617 8807 9623 8833
rect 10817 8807 10823 8833
rect 10849 8807 10855 8833
rect 11097 8807 11103 8833
rect 11129 8807 11135 8833
rect 11433 8807 11439 8833
rect 11465 8807 11471 8833
rect 11713 8807 11719 8833
rect 11745 8807 11751 8833
rect 12217 8807 12223 8833
rect 12249 8807 12255 8833
rect 10655 8777 10681 8783
rect 10655 8745 10681 8751
rect 18271 8777 18297 8783
rect 18271 8745 18297 8751
rect 18607 8777 18633 8783
rect 18607 8745 18633 8751
rect 18775 8777 18801 8783
rect 18775 8745 18801 8751
rect 18943 8777 18969 8783
rect 18943 8745 18969 8751
rect 19111 8777 19137 8783
rect 19111 8745 19137 8751
rect 8639 8721 8665 8727
rect 9473 8695 9479 8721
rect 9505 8695 9511 8721
rect 11153 8695 11159 8721
rect 11185 8695 11191 8721
rect 8639 8689 8665 8695
rect 672 8637 19400 8654
rect 672 8611 5269 8637
rect 5295 8611 5321 8637
rect 5347 8611 5373 8637
rect 5399 8611 9931 8637
rect 9957 8611 9983 8637
rect 10009 8611 10035 8637
rect 10061 8611 14593 8637
rect 14619 8611 14645 8637
rect 14671 8611 14697 8637
rect 14723 8611 19255 8637
rect 19281 8611 19307 8637
rect 19333 8611 19359 8637
rect 19385 8611 19400 8637
rect 672 8594 19400 8611
rect 855 8553 881 8559
rect 855 8521 881 8527
rect 1359 8497 1385 8503
rect 18943 8497 18969 8503
rect 1017 8471 1023 8497
rect 1049 8471 1055 8497
rect 7961 8471 7967 8497
rect 7993 8471 7999 8497
rect 1359 8465 1385 8471
rect 18943 8465 18969 8471
rect 1191 8441 1217 8447
rect 1191 8409 1217 8415
rect 1583 8441 1609 8447
rect 18775 8441 18801 8447
rect 8073 8415 8079 8441
rect 8105 8415 8111 8441
rect 1583 8409 1609 8415
rect 18775 8409 18801 8415
rect 19111 8441 19137 8447
rect 19111 8409 19137 8415
rect 672 8245 19320 8262
rect 672 8219 2938 8245
rect 2964 8219 2990 8245
rect 3016 8219 3042 8245
rect 3068 8219 7600 8245
rect 7626 8219 7652 8245
rect 7678 8219 7704 8245
rect 7730 8219 12262 8245
rect 12288 8219 12314 8245
rect 12340 8219 12366 8245
rect 12392 8219 16924 8245
rect 16950 8219 16976 8245
rect 17002 8219 17028 8245
rect 17054 8219 19320 8245
rect 672 8202 19320 8219
rect 1247 8105 1273 8111
rect 1247 8073 1273 8079
rect 19167 8105 19193 8111
rect 19167 8073 19193 8079
rect 905 8023 911 8049
rect 937 8023 943 8049
rect 7737 8023 7743 8049
rect 7769 8023 7775 8049
rect 7961 8023 7967 8049
rect 7993 8023 7999 8049
rect 8577 8023 8583 8049
rect 8609 8023 8615 8049
rect 9081 8023 9087 8049
rect 9113 8023 9119 8049
rect 7575 7993 7601 7999
rect 8303 7993 8329 7999
rect 8073 7967 8079 7993
rect 8105 7967 8111 7993
rect 7575 7961 7601 7967
rect 8303 7961 8329 7967
rect 1023 7937 1049 7943
rect 1023 7905 1049 7911
rect 9703 7937 9729 7943
rect 10039 7937 10065 7943
rect 9865 7911 9871 7937
rect 9897 7911 9903 7937
rect 10201 7911 10207 7937
rect 10233 7911 10239 7937
rect 9703 7905 9729 7911
rect 10039 7905 10065 7911
rect 672 7853 19400 7870
rect 672 7827 5269 7853
rect 5295 7827 5321 7853
rect 5347 7827 5373 7853
rect 5399 7827 9931 7853
rect 9957 7827 9983 7853
rect 10009 7827 10035 7853
rect 10061 7827 14593 7853
rect 14619 7827 14645 7853
rect 14671 7827 14697 7853
rect 14723 7827 19255 7853
rect 19281 7827 19307 7853
rect 19333 7827 19359 7853
rect 19385 7827 19400 7853
rect 672 7810 19400 7827
rect 911 7769 937 7775
rect 7905 7743 7911 7769
rect 7937 7743 7943 7769
rect 9641 7743 9647 7769
rect 9673 7743 9679 7769
rect 911 7737 937 7743
rect 7687 7713 7713 7719
rect 7687 7681 7713 7687
rect 9871 7657 9897 7663
rect 6897 7631 6903 7657
rect 6929 7631 6935 7657
rect 7289 7631 7295 7657
rect 7321 7631 7327 7657
rect 8017 7631 8023 7657
rect 8049 7631 8055 7657
rect 8241 7631 8247 7657
rect 8273 7631 8279 7657
rect 9305 7631 9311 7657
rect 9337 7631 9343 7657
rect 9585 7631 9591 7657
rect 9617 7631 9623 7657
rect 10257 7631 10263 7657
rect 10289 7631 10295 7657
rect 10705 7631 10711 7657
rect 10737 7631 10743 7657
rect 17817 7631 17823 7657
rect 17849 7631 17855 7657
rect 9871 7625 9897 7631
rect 8415 7601 8441 7607
rect 8415 7569 8441 7575
rect 9143 7601 9169 7607
rect 9143 7569 9169 7575
rect 18999 7601 19025 7607
rect 18999 7569 19025 7575
rect 672 7461 19320 7478
rect 672 7435 2938 7461
rect 2964 7435 2990 7461
rect 3016 7435 3042 7461
rect 3068 7435 7600 7461
rect 7626 7435 7652 7461
rect 7678 7435 7704 7461
rect 7730 7435 12262 7461
rect 12288 7435 12314 7461
rect 12340 7435 12366 7461
rect 12392 7435 16924 7461
rect 16950 7435 16976 7461
rect 17002 7435 17028 7461
rect 17054 7435 19320 7461
rect 672 7418 19320 7435
rect 18831 7321 18857 7327
rect 18831 7289 18857 7295
rect 9479 7265 9505 7271
rect 19111 7265 19137 7271
rect 8185 7239 8191 7265
rect 8217 7239 8223 7265
rect 8913 7239 8919 7265
rect 8945 7239 8951 7265
rect 9193 7239 9199 7265
rect 9225 7239 9231 7265
rect 9865 7239 9871 7265
rect 9897 7239 9903 7265
rect 10313 7239 10319 7265
rect 10345 7239 10351 7265
rect 9479 7233 9505 7239
rect 19111 7233 19137 7239
rect 8751 7209 8777 7215
rect 18943 7209 18969 7215
rect 9249 7183 9255 7209
rect 9281 7183 9287 7209
rect 8751 7177 8777 7183
rect 18943 7177 18969 7183
rect 8073 7127 8079 7153
rect 8105 7127 8111 7153
rect 672 7069 19400 7086
rect 672 7043 5269 7069
rect 5295 7043 5321 7069
rect 5347 7043 5373 7069
rect 5399 7043 9931 7069
rect 9957 7043 9983 7069
rect 10009 7043 10035 7069
rect 10061 7043 14593 7069
rect 14619 7043 14645 7069
rect 14671 7043 14697 7069
rect 14723 7043 19255 7069
rect 19281 7043 19307 7069
rect 19333 7043 19359 7069
rect 19385 7043 19400 7069
rect 672 7026 19400 7043
rect 17873 6847 17879 6873
rect 17905 6847 17911 6873
rect 17655 6817 17681 6823
rect 17655 6785 17681 6791
rect 18999 6817 19025 6823
rect 18999 6785 19025 6791
rect 672 6677 19320 6694
rect 672 6651 2938 6677
rect 2964 6651 2990 6677
rect 3016 6651 3042 6677
rect 3068 6651 7600 6677
rect 7626 6651 7652 6677
rect 7678 6651 7704 6677
rect 7730 6651 12262 6677
rect 12288 6651 12314 6677
rect 12340 6651 12366 6677
rect 12392 6651 16924 6677
rect 16950 6651 16976 6677
rect 17002 6651 17028 6677
rect 17054 6651 19320 6677
rect 672 6634 19320 6651
rect 672 6285 19400 6302
rect 672 6259 5269 6285
rect 5295 6259 5321 6285
rect 5347 6259 5373 6285
rect 5399 6259 9931 6285
rect 9957 6259 9983 6285
rect 10009 6259 10035 6285
rect 10061 6259 14593 6285
rect 14619 6259 14645 6285
rect 14671 6259 14697 6285
rect 14723 6259 19255 6285
rect 19281 6259 19307 6285
rect 19333 6259 19359 6285
rect 19385 6259 19400 6285
rect 672 6242 19400 6259
rect 672 5893 19320 5910
rect 672 5867 2938 5893
rect 2964 5867 2990 5893
rect 3016 5867 3042 5893
rect 3068 5867 7600 5893
rect 7626 5867 7652 5893
rect 7678 5867 7704 5893
rect 7730 5867 12262 5893
rect 12288 5867 12314 5893
rect 12340 5867 12366 5893
rect 12392 5867 16924 5893
rect 16950 5867 16976 5893
rect 17002 5867 17028 5893
rect 17054 5867 19320 5893
rect 672 5850 19320 5867
rect 672 5501 19400 5518
rect 672 5475 5269 5501
rect 5295 5475 5321 5501
rect 5347 5475 5373 5501
rect 5399 5475 9931 5501
rect 9957 5475 9983 5501
rect 10009 5475 10035 5501
rect 10061 5475 14593 5501
rect 14619 5475 14645 5501
rect 14671 5475 14697 5501
rect 14723 5475 19255 5501
rect 19281 5475 19307 5501
rect 19333 5475 19359 5501
rect 19385 5475 19400 5501
rect 672 5458 19400 5475
rect 672 5109 19320 5126
rect 672 5083 2938 5109
rect 2964 5083 2990 5109
rect 3016 5083 3042 5109
rect 3068 5083 7600 5109
rect 7626 5083 7652 5109
rect 7678 5083 7704 5109
rect 7730 5083 12262 5109
rect 12288 5083 12314 5109
rect 12340 5083 12366 5109
rect 12392 5083 16924 5109
rect 16950 5083 16976 5109
rect 17002 5083 17028 5109
rect 17054 5083 19320 5109
rect 672 5066 19320 5083
rect 672 4717 19400 4734
rect 672 4691 5269 4717
rect 5295 4691 5321 4717
rect 5347 4691 5373 4717
rect 5399 4691 9931 4717
rect 9957 4691 9983 4717
rect 10009 4691 10035 4717
rect 10061 4691 14593 4717
rect 14619 4691 14645 4717
rect 14671 4691 14697 4717
rect 14723 4691 19255 4717
rect 19281 4691 19307 4717
rect 19333 4691 19359 4717
rect 19385 4691 19400 4717
rect 672 4674 19400 4691
rect 672 4325 19320 4342
rect 672 4299 2938 4325
rect 2964 4299 2990 4325
rect 3016 4299 3042 4325
rect 3068 4299 7600 4325
rect 7626 4299 7652 4325
rect 7678 4299 7704 4325
rect 7730 4299 12262 4325
rect 12288 4299 12314 4325
rect 12340 4299 12366 4325
rect 12392 4299 16924 4325
rect 16950 4299 16976 4325
rect 17002 4299 17028 4325
rect 17054 4299 19320 4325
rect 672 4282 19320 4299
rect 672 3933 19400 3950
rect 672 3907 5269 3933
rect 5295 3907 5321 3933
rect 5347 3907 5373 3933
rect 5399 3907 9931 3933
rect 9957 3907 9983 3933
rect 10009 3907 10035 3933
rect 10061 3907 14593 3933
rect 14619 3907 14645 3933
rect 14671 3907 14697 3933
rect 14723 3907 19255 3933
rect 19281 3907 19307 3933
rect 19333 3907 19359 3933
rect 19385 3907 19400 3933
rect 672 3890 19400 3907
rect 672 3541 19320 3558
rect 672 3515 2938 3541
rect 2964 3515 2990 3541
rect 3016 3515 3042 3541
rect 3068 3515 7600 3541
rect 7626 3515 7652 3541
rect 7678 3515 7704 3541
rect 7730 3515 12262 3541
rect 12288 3515 12314 3541
rect 12340 3515 12366 3541
rect 12392 3515 16924 3541
rect 16950 3515 16976 3541
rect 17002 3515 17028 3541
rect 17054 3515 19320 3541
rect 672 3498 19320 3515
rect 672 3149 19400 3166
rect 672 3123 5269 3149
rect 5295 3123 5321 3149
rect 5347 3123 5373 3149
rect 5399 3123 9931 3149
rect 9957 3123 9983 3149
rect 10009 3123 10035 3149
rect 10061 3123 14593 3149
rect 14619 3123 14645 3149
rect 14671 3123 14697 3149
rect 14723 3123 19255 3149
rect 19281 3123 19307 3149
rect 19333 3123 19359 3149
rect 19385 3123 19400 3149
rect 672 3106 19400 3123
rect 672 2757 19320 2774
rect 672 2731 2938 2757
rect 2964 2731 2990 2757
rect 3016 2731 3042 2757
rect 3068 2731 7600 2757
rect 7626 2731 7652 2757
rect 7678 2731 7704 2757
rect 7730 2731 12262 2757
rect 12288 2731 12314 2757
rect 12340 2731 12366 2757
rect 12392 2731 16924 2757
rect 16950 2731 16976 2757
rect 17002 2731 17028 2757
rect 17054 2731 19320 2757
rect 672 2714 19320 2731
rect 7407 2561 7433 2567
rect 7407 2529 7433 2535
rect 7743 2449 7769 2455
rect 7743 2417 7769 2423
rect 8079 2449 8105 2455
rect 8079 2417 8105 2423
rect 8359 2449 8385 2455
rect 8359 2417 8385 2423
rect 672 2365 19400 2382
rect 672 2339 5269 2365
rect 5295 2339 5321 2365
rect 5347 2339 5373 2365
rect 5399 2339 9931 2365
rect 9957 2339 9983 2365
rect 10009 2339 10035 2365
rect 10061 2339 14593 2365
rect 14619 2339 14645 2365
rect 14671 2339 14697 2365
rect 14723 2339 19255 2365
rect 19281 2339 19307 2365
rect 19333 2339 19359 2365
rect 19385 2339 19400 2365
rect 672 2322 19400 2339
rect 6735 2281 6761 2287
rect 6735 2249 6761 2255
rect 7015 2281 7041 2287
rect 7015 2249 7041 2255
rect 7351 2281 7377 2287
rect 7351 2249 7377 2255
rect 7687 2281 7713 2287
rect 7687 2249 7713 2255
rect 8023 2281 8049 2287
rect 8023 2249 8049 2255
rect 8191 2281 8217 2287
rect 8191 2249 8217 2255
rect 7855 2225 7881 2231
rect 7855 2193 7881 2199
rect 6847 2169 6873 2175
rect 6847 2137 6873 2143
rect 7183 2169 7209 2175
rect 7569 2143 7575 2169
rect 7601 2143 7607 2169
rect 8297 2143 8303 2169
rect 8329 2143 8335 2169
rect 12609 2143 12615 2169
rect 12641 2143 12647 2169
rect 7183 2137 7209 2143
rect 6511 2113 6537 2119
rect 6511 2081 6537 2087
rect 8863 2113 8889 2119
rect 8863 2081 8889 2087
rect 9199 2113 9225 2119
rect 9199 2081 9225 2087
rect 9535 2113 9561 2119
rect 9535 2081 9561 2087
rect 9871 2113 9897 2119
rect 9871 2081 9897 2087
rect 10151 2113 10177 2119
rect 10151 2081 10177 2087
rect 10431 2113 10457 2119
rect 10431 2081 10457 2087
rect 10767 2113 10793 2119
rect 10767 2081 10793 2087
rect 11103 2113 11129 2119
rect 11103 2081 11129 2087
rect 11439 2113 11465 2119
rect 11439 2081 11465 2087
rect 13119 2057 13145 2063
rect 13119 2025 13145 2031
rect 672 1973 19320 1990
rect 672 1947 2938 1973
rect 2964 1947 2990 1973
rect 3016 1947 3042 1973
rect 3068 1947 7600 1973
rect 7626 1947 7652 1973
rect 7678 1947 7704 1973
rect 7730 1947 12262 1973
rect 12288 1947 12314 1973
rect 12340 1947 12366 1973
rect 12392 1947 16924 1973
rect 16950 1947 16976 1973
rect 17002 1947 17028 1973
rect 17054 1947 19320 1973
rect 672 1930 19320 1947
rect 6679 1833 6705 1839
rect 6679 1801 6705 1807
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 9423 1777 9449 1783
rect 7793 1751 7799 1777
rect 7825 1751 7831 1777
rect 8633 1751 8639 1777
rect 8665 1751 8671 1777
rect 8969 1751 8975 1777
rect 9001 1751 9007 1777
rect 9423 1745 9449 1751
rect 9759 1777 9785 1783
rect 9759 1745 9785 1751
rect 10095 1777 10121 1783
rect 10649 1751 10655 1777
rect 10681 1751 10687 1777
rect 10985 1751 10991 1777
rect 11017 1751 11023 1777
rect 11321 1751 11327 1777
rect 11353 1751 11359 1777
rect 11657 1751 11663 1777
rect 11689 1751 11695 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 10095 1745 10121 1751
rect 8023 1721 8049 1727
rect 8023 1689 8049 1695
rect 8191 1721 8217 1727
rect 8191 1689 8217 1695
rect 8751 1721 8777 1727
rect 8751 1689 8777 1695
rect 9087 1721 9113 1727
rect 9087 1689 9113 1695
rect 9255 1721 9281 1727
rect 9255 1689 9281 1695
rect 9591 1721 9617 1727
rect 9591 1689 9617 1695
rect 9927 1721 9953 1727
rect 9927 1689 9953 1695
rect 10543 1721 10569 1727
rect 10543 1689 10569 1695
rect 10879 1721 10905 1727
rect 10879 1689 10905 1695
rect 11215 1721 11241 1727
rect 11215 1689 11241 1695
rect 11551 1665 11577 1671
rect 11551 1633 11577 1639
rect 672 1581 19400 1598
rect 672 1555 5269 1581
rect 5295 1555 5321 1581
rect 5347 1555 5373 1581
rect 5399 1555 9931 1581
rect 9957 1555 9983 1581
rect 10009 1555 10035 1581
rect 10061 1555 14593 1581
rect 14619 1555 14645 1581
rect 14671 1555 14697 1581
rect 14723 1555 19255 1581
rect 19281 1555 19307 1581
rect 19333 1555 19359 1581
rect 19385 1555 19400 1581
rect 672 1538 19400 1555
<< via1 >>
rect 2938 18411 2964 18437
rect 2990 18411 3016 18437
rect 3042 18411 3068 18437
rect 7600 18411 7626 18437
rect 7652 18411 7678 18437
rect 7704 18411 7730 18437
rect 12262 18411 12288 18437
rect 12314 18411 12340 18437
rect 12366 18411 12392 18437
rect 16924 18411 16950 18437
rect 16976 18411 17002 18437
rect 17028 18411 17054 18437
rect 9031 18327 9057 18353
rect 7407 18271 7433 18297
rect 10151 18271 10177 18297
rect 8191 18215 8217 18241
rect 8639 18215 8665 18241
rect 10655 18215 10681 18241
rect 10879 18215 10905 18241
rect 11327 18215 11353 18241
rect 10543 18103 10569 18129
rect 11047 18103 11073 18129
rect 11215 18103 11241 18129
rect 5269 18019 5295 18045
rect 5321 18019 5347 18045
rect 5373 18019 5399 18045
rect 9931 18019 9957 18045
rect 9983 18019 10009 18045
rect 10035 18019 10061 18045
rect 14593 18019 14619 18045
rect 14645 18019 14671 18045
rect 14697 18019 14723 18045
rect 19255 18019 19281 18045
rect 19307 18019 19333 18045
rect 19359 18019 19385 18045
rect 7519 17935 7545 17961
rect 9871 17935 9897 17961
rect 10767 17935 10793 17961
rect 11103 17935 11129 17961
rect 7855 17879 7881 17905
rect 8023 17879 8049 17905
rect 8191 17879 8217 17905
rect 8359 17879 8385 17905
rect 8863 17879 8889 17905
rect 9031 17879 9057 17905
rect 9199 17879 9225 17905
rect 9535 17879 9561 17905
rect 10207 17879 10233 17905
rect 10375 17879 10401 17905
rect 9311 17823 9337 17849
rect 9647 17823 9673 17849
rect 9983 17823 10009 17849
rect 7743 17767 7769 17793
rect 2938 17627 2964 17653
rect 2990 17627 3016 17653
rect 3042 17627 3068 17653
rect 7600 17627 7626 17653
rect 7652 17627 7678 17653
rect 7704 17627 7730 17653
rect 12262 17627 12288 17653
rect 12314 17627 12340 17653
rect 12366 17627 12392 17653
rect 16924 17627 16950 17653
rect 16976 17627 17002 17653
rect 17028 17627 17054 17653
rect 8751 17487 8777 17513
rect 9087 17487 9113 17513
rect 9423 17487 9449 17513
rect 9759 17487 9785 17513
rect 10095 17487 10121 17513
rect 5269 17235 5295 17261
rect 5321 17235 5347 17261
rect 5373 17235 5399 17261
rect 9931 17235 9957 17261
rect 9983 17235 10009 17261
rect 10035 17235 10061 17261
rect 14593 17235 14619 17261
rect 14645 17235 14671 17261
rect 14697 17235 14723 17261
rect 19255 17235 19281 17261
rect 19307 17235 19333 17261
rect 19359 17235 19385 17261
rect 2938 16843 2964 16869
rect 2990 16843 3016 16869
rect 3042 16843 3068 16869
rect 7600 16843 7626 16869
rect 7652 16843 7678 16869
rect 7704 16843 7730 16869
rect 12262 16843 12288 16869
rect 12314 16843 12340 16869
rect 12366 16843 12392 16869
rect 16924 16843 16950 16869
rect 16976 16843 17002 16869
rect 17028 16843 17054 16869
rect 5269 16451 5295 16477
rect 5321 16451 5347 16477
rect 5373 16451 5399 16477
rect 9931 16451 9957 16477
rect 9983 16451 10009 16477
rect 10035 16451 10061 16477
rect 14593 16451 14619 16477
rect 14645 16451 14671 16477
rect 14697 16451 14723 16477
rect 19255 16451 19281 16477
rect 19307 16451 19333 16477
rect 19359 16451 19385 16477
rect 2938 16059 2964 16085
rect 2990 16059 3016 16085
rect 3042 16059 3068 16085
rect 7600 16059 7626 16085
rect 7652 16059 7678 16085
rect 7704 16059 7730 16085
rect 12262 16059 12288 16085
rect 12314 16059 12340 16085
rect 12366 16059 12392 16085
rect 16924 16059 16950 16085
rect 16976 16059 17002 16085
rect 17028 16059 17054 16085
rect 5269 15667 5295 15693
rect 5321 15667 5347 15693
rect 5373 15667 5399 15693
rect 9931 15667 9957 15693
rect 9983 15667 10009 15693
rect 10035 15667 10061 15693
rect 14593 15667 14619 15693
rect 14645 15667 14671 15693
rect 14697 15667 14723 15693
rect 19255 15667 19281 15693
rect 19307 15667 19333 15693
rect 19359 15667 19385 15693
rect 2938 15275 2964 15301
rect 2990 15275 3016 15301
rect 3042 15275 3068 15301
rect 7600 15275 7626 15301
rect 7652 15275 7678 15301
rect 7704 15275 7730 15301
rect 12262 15275 12288 15301
rect 12314 15275 12340 15301
rect 12366 15275 12392 15301
rect 16924 15275 16950 15301
rect 16976 15275 17002 15301
rect 17028 15275 17054 15301
rect 5269 14883 5295 14909
rect 5321 14883 5347 14909
rect 5373 14883 5399 14909
rect 9931 14883 9957 14909
rect 9983 14883 10009 14909
rect 10035 14883 10061 14909
rect 14593 14883 14619 14909
rect 14645 14883 14671 14909
rect 14697 14883 14723 14909
rect 19255 14883 19281 14909
rect 19307 14883 19333 14909
rect 19359 14883 19385 14909
rect 2938 14491 2964 14517
rect 2990 14491 3016 14517
rect 3042 14491 3068 14517
rect 7600 14491 7626 14517
rect 7652 14491 7678 14517
rect 7704 14491 7730 14517
rect 12262 14491 12288 14517
rect 12314 14491 12340 14517
rect 12366 14491 12392 14517
rect 16924 14491 16950 14517
rect 16976 14491 17002 14517
rect 17028 14491 17054 14517
rect 5269 14099 5295 14125
rect 5321 14099 5347 14125
rect 5373 14099 5399 14125
rect 9931 14099 9957 14125
rect 9983 14099 10009 14125
rect 10035 14099 10061 14125
rect 14593 14099 14619 14125
rect 14645 14099 14671 14125
rect 14697 14099 14723 14125
rect 19255 14099 19281 14125
rect 19307 14099 19333 14125
rect 19359 14099 19385 14125
rect 2938 13707 2964 13733
rect 2990 13707 3016 13733
rect 3042 13707 3068 13733
rect 7600 13707 7626 13733
rect 7652 13707 7678 13733
rect 7704 13707 7730 13733
rect 12262 13707 12288 13733
rect 12314 13707 12340 13733
rect 12366 13707 12392 13733
rect 16924 13707 16950 13733
rect 16976 13707 17002 13733
rect 17028 13707 17054 13733
rect 5269 13315 5295 13341
rect 5321 13315 5347 13341
rect 5373 13315 5399 13341
rect 9931 13315 9957 13341
rect 9983 13315 10009 13341
rect 10035 13315 10061 13341
rect 14593 13315 14619 13341
rect 14645 13315 14671 13341
rect 14697 13315 14723 13341
rect 19255 13315 19281 13341
rect 19307 13315 19333 13341
rect 19359 13315 19385 13341
rect 2143 13119 2169 13145
rect 2423 13063 2449 13089
rect 967 13007 993 13033
rect 2938 12923 2964 12949
rect 2990 12923 3016 12949
rect 3042 12923 3068 12949
rect 7600 12923 7626 12949
rect 7652 12923 7678 12949
rect 7704 12923 7730 12949
rect 12262 12923 12288 12949
rect 12314 12923 12340 12949
rect 12366 12923 12392 12949
rect 16924 12923 16950 12949
rect 16976 12923 17002 12949
rect 17028 12923 17054 12949
rect 855 12671 881 12697
rect 1023 12615 1049 12641
rect 1247 12615 1273 12641
rect 5269 12531 5295 12557
rect 5321 12531 5347 12557
rect 5373 12531 5399 12557
rect 9931 12531 9957 12557
rect 9983 12531 10009 12557
rect 10035 12531 10061 12557
rect 14593 12531 14619 12557
rect 14645 12531 14671 12557
rect 14697 12531 14723 12557
rect 19255 12531 19281 12557
rect 19307 12531 19333 12557
rect 19359 12531 19385 12557
rect 8695 12447 8721 12473
rect 1023 12391 1049 12417
rect 855 12335 881 12361
rect 8807 12335 8833 12361
rect 17823 12335 17849 12361
rect 1247 12279 1273 12305
rect 18999 12223 19025 12249
rect 2938 12139 2964 12165
rect 2990 12139 3016 12165
rect 3042 12139 3068 12165
rect 7600 12139 7626 12165
rect 7652 12139 7678 12165
rect 7704 12139 7730 12165
rect 12262 12139 12288 12165
rect 12314 12139 12340 12165
rect 12366 12139 12392 12165
rect 16924 12139 16950 12165
rect 16976 12139 17002 12165
rect 17028 12139 17054 12165
rect 8023 11999 8049 12025
rect 8191 11943 8217 11969
rect 8415 11943 8441 11969
rect 8863 11943 8889 11969
rect 9087 11943 9113 11969
rect 9535 11943 9561 11969
rect 855 11887 881 11913
rect 19111 11887 19137 11913
rect 1023 11831 1049 11857
rect 1247 11831 1273 11857
rect 8527 11831 8553 11857
rect 18831 11831 18857 11857
rect 18943 11831 18969 11857
rect 5269 11747 5295 11773
rect 5321 11747 5347 11773
rect 5373 11747 5399 11773
rect 9931 11747 9957 11773
rect 9983 11747 10009 11773
rect 10035 11747 10061 11773
rect 14593 11747 14619 11773
rect 14645 11747 14671 11773
rect 14697 11747 14723 11773
rect 19255 11747 19281 11773
rect 19307 11747 19333 11773
rect 19359 11747 19385 11773
rect 1023 11607 1049 11633
rect 8695 11607 8721 11633
rect 18943 11607 18969 11633
rect 855 11551 881 11577
rect 8807 11551 8833 11577
rect 19111 11551 19137 11577
rect 1247 11495 1273 11521
rect 18831 11495 18857 11521
rect 2938 11355 2964 11381
rect 2990 11355 3016 11381
rect 3042 11355 3068 11381
rect 7600 11355 7626 11381
rect 7652 11355 7678 11381
rect 7704 11355 7730 11381
rect 12262 11355 12288 11381
rect 12314 11355 12340 11381
rect 12366 11355 12392 11381
rect 16924 11355 16950 11381
rect 16976 11355 17002 11381
rect 17028 11355 17054 11381
rect 8023 11215 8049 11241
rect 8191 11159 8217 11185
rect 8415 11159 8441 11185
rect 8863 11159 8889 11185
rect 9143 11159 9169 11185
rect 9591 11159 9617 11185
rect 855 11103 881 11129
rect 1023 11103 1049 11129
rect 1191 11103 1217 11129
rect 8527 11103 8553 11129
rect 11215 11103 11241 11129
rect 18831 11103 18857 11129
rect 19111 11103 19137 11129
rect 1359 11047 1385 11073
rect 1583 11047 1609 11073
rect 10711 11047 10737 11073
rect 10879 11047 10905 11073
rect 11047 11047 11073 11073
rect 18943 11047 18969 11073
rect 5269 10963 5295 10989
rect 5321 10963 5347 10989
rect 5373 10963 5399 10989
rect 9931 10963 9957 10989
rect 9983 10963 10009 10989
rect 10035 10963 10061 10989
rect 14593 10963 14619 10989
rect 14645 10963 14671 10989
rect 14697 10963 14723 10989
rect 19255 10963 19281 10989
rect 19307 10963 19333 10989
rect 19359 10963 19385 10989
rect 1247 10879 1273 10905
rect 10991 10879 11017 10905
rect 1023 10823 1049 10849
rect 10487 10823 10513 10849
rect 855 10767 881 10793
rect 10711 10767 10737 10793
rect 10935 10767 10961 10793
rect 11327 10767 11353 10793
rect 11607 10767 11633 10793
rect 12055 10767 12081 10793
rect 17823 10767 17849 10793
rect 1471 10711 1497 10737
rect 18999 10711 19025 10737
rect 2938 10571 2964 10597
rect 2990 10571 3016 10597
rect 3042 10571 3068 10597
rect 7600 10571 7626 10597
rect 7652 10571 7678 10597
rect 7704 10571 7730 10597
rect 12262 10571 12288 10597
rect 12314 10571 12340 10597
rect 12366 10571 12392 10597
rect 16924 10571 16950 10597
rect 16976 10571 17002 10597
rect 17028 10571 17054 10597
rect 7855 10431 7881 10457
rect 10655 10431 10681 10457
rect 18271 10431 18297 10457
rect 8079 10375 8105 10401
rect 8247 10375 8273 10401
rect 8695 10375 8721 10401
rect 8863 10375 8889 10401
rect 9423 10375 9449 10401
rect 10823 10375 10849 10401
rect 11047 10375 11073 10401
rect 11383 10375 11409 10401
rect 11719 10375 11745 10401
rect 12223 10375 12249 10401
rect 19111 10375 19137 10401
rect 855 10319 881 10345
rect 7743 10319 7769 10345
rect 11159 10319 11185 10345
rect 18775 10319 18801 10345
rect 18943 10319 18969 10345
rect 1023 10263 1049 10289
rect 1247 10263 1273 10289
rect 8359 10263 8385 10289
rect 18607 10263 18633 10289
rect 5269 10179 5295 10205
rect 5321 10179 5347 10205
rect 5373 10179 5399 10205
rect 9931 10179 9957 10205
rect 9983 10179 10009 10205
rect 10035 10179 10061 10205
rect 14593 10179 14619 10205
rect 14645 10179 14671 10205
rect 14697 10179 14723 10205
rect 19255 10179 19281 10205
rect 19307 10179 19333 10205
rect 19359 10179 19385 10205
rect 18831 10095 18857 10121
rect 8247 10039 8273 10065
rect 8695 10039 8721 10065
rect 18943 10039 18969 10065
rect 2143 9983 2169 10009
rect 8359 9983 8385 10009
rect 8807 9983 8833 10009
rect 19111 9983 19137 10009
rect 9535 9927 9561 9953
rect 18607 9927 18633 9953
rect 967 9871 993 9897
rect 2938 9787 2964 9813
rect 2990 9787 3016 9813
rect 3042 9787 3068 9813
rect 7600 9787 7626 9813
rect 7652 9787 7678 9813
rect 7704 9787 7730 9813
rect 12262 9787 12288 9813
rect 12314 9787 12340 9813
rect 12366 9787 12392 9813
rect 16924 9787 16950 9813
rect 16976 9787 17002 9813
rect 17028 9787 17054 9813
rect 9927 9647 9953 9673
rect 8023 9591 8049 9617
rect 8247 9591 8273 9617
rect 8695 9591 8721 9617
rect 8975 9591 9001 9617
rect 9367 9591 9393 9617
rect 855 9535 881 9561
rect 7743 9535 7769 9561
rect 7855 9535 7881 9561
rect 8359 9535 8385 9561
rect 18831 9535 18857 9561
rect 19111 9535 19137 9561
rect 1023 9479 1049 9505
rect 1247 9479 1273 9505
rect 9647 9479 9673 9505
rect 10095 9479 10121 9505
rect 10263 9479 10289 9505
rect 11159 9479 11185 9505
rect 11327 9479 11353 9505
rect 11495 9479 11521 9505
rect 11663 9479 11689 9505
rect 18943 9479 18969 9505
rect 5269 9395 5295 9421
rect 5321 9395 5347 9421
rect 5373 9395 5399 9421
rect 9931 9395 9957 9421
rect 9983 9395 10009 9421
rect 10035 9395 10061 9421
rect 14593 9395 14619 9421
rect 14645 9395 14671 9421
rect 14697 9395 14723 9421
rect 19255 9395 19281 9421
rect 19307 9395 19333 9421
rect 19359 9395 19385 9421
rect 9143 9311 9169 9337
rect 11103 9311 11129 9337
rect 1023 9255 1049 9281
rect 18943 9255 18969 9281
rect 855 9199 881 9225
rect 8695 9199 8721 9225
rect 8919 9199 8945 9225
rect 9311 9199 9337 9225
rect 10823 9199 10849 9225
rect 11047 9199 11073 9225
rect 11327 9199 11353 9225
rect 11719 9199 11745 9225
rect 12167 9199 12193 9225
rect 19111 9199 19137 9225
rect 1247 9143 1273 9169
rect 8415 9143 8441 9169
rect 10599 9143 10625 9169
rect 12671 9143 12697 9169
rect 12951 9143 12977 9169
rect 18831 9143 18857 9169
rect 2938 9003 2964 9029
rect 2990 9003 3016 9029
rect 3042 9003 3068 9029
rect 7600 9003 7626 9029
rect 7652 9003 7678 9029
rect 7704 9003 7730 9029
rect 12262 9003 12288 9029
rect 12314 9003 12340 9029
rect 12366 9003 12392 9029
rect 16924 9003 16950 9029
rect 16976 9003 17002 9029
rect 17028 9003 17054 9029
rect 967 8863 993 8889
rect 8863 8863 8889 8889
rect 2143 8807 2169 8833
rect 9031 8807 9057 8833
rect 9591 8807 9617 8833
rect 10823 8807 10849 8833
rect 11103 8807 11129 8833
rect 11439 8807 11465 8833
rect 11719 8807 11745 8833
rect 12223 8807 12249 8833
rect 10655 8751 10681 8777
rect 18271 8751 18297 8777
rect 18607 8751 18633 8777
rect 18775 8751 18801 8777
rect 18943 8751 18969 8777
rect 19111 8751 19137 8777
rect 8639 8695 8665 8721
rect 9479 8695 9505 8721
rect 11159 8695 11185 8721
rect 5269 8611 5295 8637
rect 5321 8611 5347 8637
rect 5373 8611 5399 8637
rect 9931 8611 9957 8637
rect 9983 8611 10009 8637
rect 10035 8611 10061 8637
rect 14593 8611 14619 8637
rect 14645 8611 14671 8637
rect 14697 8611 14723 8637
rect 19255 8611 19281 8637
rect 19307 8611 19333 8637
rect 19359 8611 19385 8637
rect 855 8527 881 8553
rect 1023 8471 1049 8497
rect 1359 8471 1385 8497
rect 7967 8471 7993 8497
rect 18943 8471 18969 8497
rect 1191 8415 1217 8441
rect 1583 8415 1609 8441
rect 8079 8415 8105 8441
rect 18775 8415 18801 8441
rect 19111 8415 19137 8441
rect 2938 8219 2964 8245
rect 2990 8219 3016 8245
rect 3042 8219 3068 8245
rect 7600 8219 7626 8245
rect 7652 8219 7678 8245
rect 7704 8219 7730 8245
rect 12262 8219 12288 8245
rect 12314 8219 12340 8245
rect 12366 8219 12392 8245
rect 16924 8219 16950 8245
rect 16976 8219 17002 8245
rect 17028 8219 17054 8245
rect 1247 8079 1273 8105
rect 19167 8079 19193 8105
rect 911 8023 937 8049
rect 7743 8023 7769 8049
rect 7967 8023 7993 8049
rect 8583 8023 8609 8049
rect 9087 8023 9113 8049
rect 7575 7967 7601 7993
rect 8079 7967 8105 7993
rect 8303 7967 8329 7993
rect 1023 7911 1049 7937
rect 9703 7911 9729 7937
rect 9871 7911 9897 7937
rect 10039 7911 10065 7937
rect 10207 7911 10233 7937
rect 5269 7827 5295 7853
rect 5321 7827 5347 7853
rect 5373 7827 5399 7853
rect 9931 7827 9957 7853
rect 9983 7827 10009 7853
rect 10035 7827 10061 7853
rect 14593 7827 14619 7853
rect 14645 7827 14671 7853
rect 14697 7827 14723 7853
rect 19255 7827 19281 7853
rect 19307 7827 19333 7853
rect 19359 7827 19385 7853
rect 911 7743 937 7769
rect 7911 7743 7937 7769
rect 9647 7743 9673 7769
rect 7687 7687 7713 7713
rect 6903 7631 6929 7657
rect 7295 7631 7321 7657
rect 8023 7631 8049 7657
rect 8247 7631 8273 7657
rect 9311 7631 9337 7657
rect 9591 7631 9617 7657
rect 9871 7631 9897 7657
rect 10263 7631 10289 7657
rect 10711 7631 10737 7657
rect 17823 7631 17849 7657
rect 8415 7575 8441 7601
rect 9143 7575 9169 7601
rect 18999 7575 19025 7601
rect 2938 7435 2964 7461
rect 2990 7435 3016 7461
rect 3042 7435 3068 7461
rect 7600 7435 7626 7461
rect 7652 7435 7678 7461
rect 7704 7435 7730 7461
rect 12262 7435 12288 7461
rect 12314 7435 12340 7461
rect 12366 7435 12392 7461
rect 16924 7435 16950 7461
rect 16976 7435 17002 7461
rect 17028 7435 17054 7461
rect 18831 7295 18857 7321
rect 8191 7239 8217 7265
rect 8919 7239 8945 7265
rect 9199 7239 9225 7265
rect 9479 7239 9505 7265
rect 9871 7239 9897 7265
rect 10319 7239 10345 7265
rect 19111 7239 19137 7265
rect 8751 7183 8777 7209
rect 9255 7183 9281 7209
rect 18943 7183 18969 7209
rect 8079 7127 8105 7153
rect 5269 7043 5295 7069
rect 5321 7043 5347 7069
rect 5373 7043 5399 7069
rect 9931 7043 9957 7069
rect 9983 7043 10009 7069
rect 10035 7043 10061 7069
rect 14593 7043 14619 7069
rect 14645 7043 14671 7069
rect 14697 7043 14723 7069
rect 19255 7043 19281 7069
rect 19307 7043 19333 7069
rect 19359 7043 19385 7069
rect 17879 6847 17905 6873
rect 17655 6791 17681 6817
rect 18999 6791 19025 6817
rect 2938 6651 2964 6677
rect 2990 6651 3016 6677
rect 3042 6651 3068 6677
rect 7600 6651 7626 6677
rect 7652 6651 7678 6677
rect 7704 6651 7730 6677
rect 12262 6651 12288 6677
rect 12314 6651 12340 6677
rect 12366 6651 12392 6677
rect 16924 6651 16950 6677
rect 16976 6651 17002 6677
rect 17028 6651 17054 6677
rect 5269 6259 5295 6285
rect 5321 6259 5347 6285
rect 5373 6259 5399 6285
rect 9931 6259 9957 6285
rect 9983 6259 10009 6285
rect 10035 6259 10061 6285
rect 14593 6259 14619 6285
rect 14645 6259 14671 6285
rect 14697 6259 14723 6285
rect 19255 6259 19281 6285
rect 19307 6259 19333 6285
rect 19359 6259 19385 6285
rect 2938 5867 2964 5893
rect 2990 5867 3016 5893
rect 3042 5867 3068 5893
rect 7600 5867 7626 5893
rect 7652 5867 7678 5893
rect 7704 5867 7730 5893
rect 12262 5867 12288 5893
rect 12314 5867 12340 5893
rect 12366 5867 12392 5893
rect 16924 5867 16950 5893
rect 16976 5867 17002 5893
rect 17028 5867 17054 5893
rect 5269 5475 5295 5501
rect 5321 5475 5347 5501
rect 5373 5475 5399 5501
rect 9931 5475 9957 5501
rect 9983 5475 10009 5501
rect 10035 5475 10061 5501
rect 14593 5475 14619 5501
rect 14645 5475 14671 5501
rect 14697 5475 14723 5501
rect 19255 5475 19281 5501
rect 19307 5475 19333 5501
rect 19359 5475 19385 5501
rect 2938 5083 2964 5109
rect 2990 5083 3016 5109
rect 3042 5083 3068 5109
rect 7600 5083 7626 5109
rect 7652 5083 7678 5109
rect 7704 5083 7730 5109
rect 12262 5083 12288 5109
rect 12314 5083 12340 5109
rect 12366 5083 12392 5109
rect 16924 5083 16950 5109
rect 16976 5083 17002 5109
rect 17028 5083 17054 5109
rect 5269 4691 5295 4717
rect 5321 4691 5347 4717
rect 5373 4691 5399 4717
rect 9931 4691 9957 4717
rect 9983 4691 10009 4717
rect 10035 4691 10061 4717
rect 14593 4691 14619 4717
rect 14645 4691 14671 4717
rect 14697 4691 14723 4717
rect 19255 4691 19281 4717
rect 19307 4691 19333 4717
rect 19359 4691 19385 4717
rect 2938 4299 2964 4325
rect 2990 4299 3016 4325
rect 3042 4299 3068 4325
rect 7600 4299 7626 4325
rect 7652 4299 7678 4325
rect 7704 4299 7730 4325
rect 12262 4299 12288 4325
rect 12314 4299 12340 4325
rect 12366 4299 12392 4325
rect 16924 4299 16950 4325
rect 16976 4299 17002 4325
rect 17028 4299 17054 4325
rect 5269 3907 5295 3933
rect 5321 3907 5347 3933
rect 5373 3907 5399 3933
rect 9931 3907 9957 3933
rect 9983 3907 10009 3933
rect 10035 3907 10061 3933
rect 14593 3907 14619 3933
rect 14645 3907 14671 3933
rect 14697 3907 14723 3933
rect 19255 3907 19281 3933
rect 19307 3907 19333 3933
rect 19359 3907 19385 3933
rect 2938 3515 2964 3541
rect 2990 3515 3016 3541
rect 3042 3515 3068 3541
rect 7600 3515 7626 3541
rect 7652 3515 7678 3541
rect 7704 3515 7730 3541
rect 12262 3515 12288 3541
rect 12314 3515 12340 3541
rect 12366 3515 12392 3541
rect 16924 3515 16950 3541
rect 16976 3515 17002 3541
rect 17028 3515 17054 3541
rect 5269 3123 5295 3149
rect 5321 3123 5347 3149
rect 5373 3123 5399 3149
rect 9931 3123 9957 3149
rect 9983 3123 10009 3149
rect 10035 3123 10061 3149
rect 14593 3123 14619 3149
rect 14645 3123 14671 3149
rect 14697 3123 14723 3149
rect 19255 3123 19281 3149
rect 19307 3123 19333 3149
rect 19359 3123 19385 3149
rect 2938 2731 2964 2757
rect 2990 2731 3016 2757
rect 3042 2731 3068 2757
rect 7600 2731 7626 2757
rect 7652 2731 7678 2757
rect 7704 2731 7730 2757
rect 12262 2731 12288 2757
rect 12314 2731 12340 2757
rect 12366 2731 12392 2757
rect 16924 2731 16950 2757
rect 16976 2731 17002 2757
rect 17028 2731 17054 2757
rect 7407 2535 7433 2561
rect 7743 2423 7769 2449
rect 8079 2423 8105 2449
rect 8359 2423 8385 2449
rect 5269 2339 5295 2365
rect 5321 2339 5347 2365
rect 5373 2339 5399 2365
rect 9931 2339 9957 2365
rect 9983 2339 10009 2365
rect 10035 2339 10061 2365
rect 14593 2339 14619 2365
rect 14645 2339 14671 2365
rect 14697 2339 14723 2365
rect 19255 2339 19281 2365
rect 19307 2339 19333 2365
rect 19359 2339 19385 2365
rect 6735 2255 6761 2281
rect 7015 2255 7041 2281
rect 7351 2255 7377 2281
rect 7687 2255 7713 2281
rect 8023 2255 8049 2281
rect 8191 2255 8217 2281
rect 7855 2199 7881 2225
rect 6847 2143 6873 2169
rect 7183 2143 7209 2169
rect 7575 2143 7601 2169
rect 8303 2143 8329 2169
rect 12615 2143 12641 2169
rect 6511 2087 6537 2113
rect 8863 2087 8889 2113
rect 9199 2087 9225 2113
rect 9535 2087 9561 2113
rect 9871 2087 9897 2113
rect 10151 2087 10177 2113
rect 10431 2087 10457 2113
rect 10767 2087 10793 2113
rect 11103 2087 11129 2113
rect 11439 2087 11465 2113
rect 13119 2031 13145 2057
rect 2938 1947 2964 1973
rect 2990 1947 3016 1973
rect 3042 1947 3068 1973
rect 7600 1947 7626 1973
rect 7652 1947 7678 1973
rect 7704 1947 7730 1973
rect 12262 1947 12288 1973
rect 12314 1947 12340 1973
rect 12366 1947 12392 1973
rect 16924 1947 16950 1973
rect 16976 1947 17002 1973
rect 17028 1947 17054 1973
rect 6679 1807 6705 1833
rect 12783 1807 12809 1833
rect 7799 1751 7825 1777
rect 8639 1751 8665 1777
rect 8975 1751 9001 1777
rect 9423 1751 9449 1777
rect 9759 1751 9785 1777
rect 10095 1751 10121 1777
rect 10655 1751 10681 1777
rect 10991 1751 11017 1777
rect 11327 1751 11353 1777
rect 11663 1751 11689 1777
rect 12279 1751 12305 1777
rect 8023 1695 8049 1721
rect 8191 1695 8217 1721
rect 8751 1695 8777 1721
rect 9087 1695 9113 1721
rect 9255 1695 9281 1721
rect 9591 1695 9617 1721
rect 9927 1695 9953 1721
rect 10543 1695 10569 1721
rect 10879 1695 10905 1721
rect 11215 1695 11241 1721
rect 11551 1639 11577 1665
rect 5269 1555 5295 1581
rect 5321 1555 5347 1581
rect 5373 1555 5399 1581
rect 9931 1555 9957 1581
rect 9983 1555 10009 1581
rect 10035 1555 10061 1581
rect 14593 1555 14619 1581
rect 14645 1555 14671 1581
rect 14697 1555 14723 1581
rect 19255 1555 19281 1581
rect 19307 1555 19333 1581
rect 19359 1555 19385 1581
<< metal2 >>
rect 7392 19600 7448 20000
rect 7728 19600 7784 20000
rect 8064 19600 8120 20000
rect 8400 19600 8456 20000
rect 8736 19600 8792 20000
rect 9072 19600 9128 20000
rect 9408 19600 9464 20000
rect 9744 19600 9800 20000
rect 10080 19600 10136 20000
rect 10416 19600 10472 20000
rect 10752 19600 10808 20000
rect 11088 19600 11144 20000
rect 2937 18438 3069 18443
rect 2965 18410 2989 18438
rect 3017 18410 3041 18438
rect 2937 18405 3069 18410
rect 7406 18297 7434 19600
rect 7742 18522 7770 19600
rect 7742 18494 7882 18522
rect 7599 18438 7731 18443
rect 7627 18410 7651 18438
rect 7679 18410 7703 18438
rect 7599 18405 7731 18410
rect 7406 18271 7407 18297
rect 7433 18271 7434 18297
rect 7406 18265 7434 18271
rect 5268 18046 5400 18051
rect 5296 18018 5320 18046
rect 5348 18018 5372 18046
rect 5268 18013 5400 18018
rect 7518 17962 7546 17967
rect 7518 17915 7546 17934
rect 7854 17962 7882 18494
rect 8078 18018 8106 19600
rect 8414 18354 8442 19600
rect 8414 18321 8442 18326
rect 8190 18242 8218 18247
rect 8190 18241 8330 18242
rect 8190 18215 8191 18241
rect 8217 18215 8330 18241
rect 8190 18214 8330 18215
rect 8190 18209 8218 18214
rect 7854 17905 7882 17934
rect 7854 17879 7855 17905
rect 7881 17879 7882 17905
rect 7854 17873 7882 17879
rect 7910 17990 8106 18018
rect 7742 17794 7770 17799
rect 7910 17794 7938 17990
rect 7742 17793 7938 17794
rect 7742 17767 7743 17793
rect 7769 17767 7938 17793
rect 7742 17766 7938 17767
rect 8022 17905 8050 17911
rect 8022 17879 8023 17905
rect 8049 17879 8050 17905
rect 7742 17761 7770 17766
rect 2937 17654 3069 17659
rect 2965 17626 2989 17654
rect 3017 17626 3041 17654
rect 2937 17621 3069 17626
rect 7599 17654 7731 17659
rect 7627 17626 7651 17654
rect 7679 17626 7703 17654
rect 7599 17621 7731 17626
rect 5268 17262 5400 17267
rect 5296 17234 5320 17262
rect 5348 17234 5372 17262
rect 5268 17229 5400 17234
rect 2937 16870 3069 16875
rect 2965 16842 2989 16870
rect 3017 16842 3041 16870
rect 2937 16837 3069 16842
rect 7599 16870 7731 16875
rect 7627 16842 7651 16870
rect 7679 16842 7703 16870
rect 7599 16837 7731 16842
rect 5268 16478 5400 16483
rect 5296 16450 5320 16478
rect 5348 16450 5372 16478
rect 5268 16445 5400 16450
rect 2937 16086 3069 16091
rect 2965 16058 2989 16086
rect 3017 16058 3041 16086
rect 2937 16053 3069 16058
rect 7599 16086 7731 16091
rect 7627 16058 7651 16086
rect 7679 16058 7703 16086
rect 7599 16053 7731 16058
rect 5268 15694 5400 15699
rect 5296 15666 5320 15694
rect 5348 15666 5372 15694
rect 5268 15661 5400 15666
rect 2937 15302 3069 15307
rect 2965 15274 2989 15302
rect 3017 15274 3041 15302
rect 2937 15269 3069 15274
rect 7599 15302 7731 15307
rect 7627 15274 7651 15302
rect 7679 15274 7703 15302
rect 7599 15269 7731 15274
rect 8022 14994 8050 17879
rect 8078 17906 8106 17990
rect 8190 17906 8218 17911
rect 8078 17905 8218 17906
rect 8078 17879 8191 17905
rect 8217 17879 8218 17905
rect 8078 17878 8218 17879
rect 8190 17873 8218 17878
rect 8302 15106 8330 18214
rect 8638 18241 8666 18247
rect 8638 18215 8639 18241
rect 8665 18215 8666 18241
rect 8358 17905 8386 17911
rect 8358 17879 8359 17905
rect 8385 17879 8386 17905
rect 8358 15106 8386 17879
rect 8358 15078 8498 15106
rect 8302 15073 8330 15078
rect 8022 14961 8050 14966
rect 8414 14994 8442 14999
rect 5268 14910 5400 14915
rect 5296 14882 5320 14910
rect 5348 14882 5372 14910
rect 5268 14877 5400 14882
rect 2937 14518 3069 14523
rect 2965 14490 2989 14518
rect 3017 14490 3041 14518
rect 2937 14485 3069 14490
rect 7599 14518 7731 14523
rect 7627 14490 7651 14518
rect 7679 14490 7703 14518
rect 7599 14485 7731 14490
rect 5268 14126 5400 14131
rect 5296 14098 5320 14126
rect 5348 14098 5372 14126
rect 5268 14093 5400 14098
rect 2937 13734 3069 13739
rect 2965 13706 2989 13734
rect 3017 13706 3041 13734
rect 2937 13701 3069 13706
rect 7599 13734 7731 13739
rect 7627 13706 7651 13734
rect 7679 13706 7703 13734
rect 7599 13701 7731 13706
rect 5268 13342 5400 13347
rect 5296 13314 5320 13342
rect 5348 13314 5372 13342
rect 5268 13309 5400 13314
rect 2142 13145 2170 13151
rect 2142 13119 2143 13145
rect 2169 13119 2170 13145
rect 2142 13090 2170 13119
rect 2422 13090 2450 13095
rect 2142 13089 2450 13090
rect 2142 13063 2423 13089
rect 2449 13063 2450 13089
rect 2142 13062 2450 13063
rect 966 13033 994 13039
rect 966 13007 967 13033
rect 993 13007 994 13033
rect 966 12810 994 13007
rect 966 12777 994 12782
rect 854 12697 882 12703
rect 854 12671 855 12697
rect 881 12671 882 12697
rect 854 12474 882 12671
rect 1022 12642 1050 12647
rect 1022 12641 1162 12642
rect 1022 12615 1023 12641
rect 1049 12615 1162 12641
rect 1022 12614 1162 12615
rect 1022 12609 1050 12614
rect 854 12441 882 12446
rect 1022 12418 1050 12423
rect 1022 12371 1050 12390
rect 854 12361 882 12367
rect 854 12335 855 12361
rect 881 12335 882 12361
rect 854 12138 882 12335
rect 854 12105 882 12110
rect 854 11913 882 11919
rect 854 11887 855 11913
rect 881 11887 882 11913
rect 854 11802 882 11887
rect 1022 11858 1050 11863
rect 1022 11811 1050 11830
rect 854 11769 882 11774
rect 1022 11634 1050 11639
rect 1022 11633 1106 11634
rect 1022 11607 1023 11633
rect 1049 11607 1106 11633
rect 1022 11606 1106 11607
rect 1022 11601 1050 11606
rect 854 11577 882 11583
rect 854 11551 855 11577
rect 881 11551 882 11577
rect 854 11466 882 11551
rect 854 11433 882 11438
rect 1022 11186 1050 11191
rect 854 11130 882 11135
rect 854 11083 882 11102
rect 1022 11129 1050 11158
rect 1022 11103 1023 11129
rect 1049 11103 1050 11129
rect 1022 11097 1050 11103
rect 1022 10850 1050 10855
rect 1022 10803 1050 10822
rect 854 10793 882 10799
rect 854 10767 855 10793
rect 881 10767 882 10793
rect 854 10738 882 10767
rect 854 10458 882 10710
rect 854 10425 882 10430
rect 854 10345 882 10351
rect 854 10319 855 10345
rect 881 10319 882 10345
rect 854 10122 882 10319
rect 1078 10346 1106 11606
rect 1078 10313 1106 10318
rect 1022 10290 1050 10295
rect 1022 10243 1050 10262
rect 854 10089 882 10094
rect 966 9898 994 9903
rect 966 9851 994 9870
rect 854 9561 882 9567
rect 854 9535 855 9561
rect 881 9535 882 9561
rect 854 9450 882 9535
rect 1134 9562 1162 12614
rect 1246 12641 1274 12647
rect 1246 12615 1247 12641
rect 1273 12615 1274 12641
rect 1246 12474 1274 12615
rect 1246 12441 1274 12446
rect 1246 12305 1274 12311
rect 1246 12279 1247 12305
rect 1273 12279 1274 12305
rect 1246 12138 1274 12279
rect 1246 12105 1274 12110
rect 1246 11857 1274 11863
rect 1246 11831 1247 11857
rect 1273 11831 1274 11857
rect 1246 11802 1274 11831
rect 1246 11769 1274 11774
rect 1246 11521 1274 11527
rect 1246 11495 1247 11521
rect 1273 11495 1274 11521
rect 1246 11466 1274 11495
rect 1246 11433 1274 11438
rect 1190 11129 1218 11135
rect 1190 11103 1191 11129
rect 1217 11103 1218 11129
rect 1190 10794 1218 11103
rect 1246 11130 1274 11135
rect 1246 10905 1274 11102
rect 1358 11074 1386 11079
rect 1358 11027 1386 11046
rect 1582 11073 1610 11079
rect 1582 11047 1583 11073
rect 1609 11047 1610 11073
rect 1246 10879 1247 10905
rect 1273 10879 1274 10905
rect 1246 10873 1274 10879
rect 1190 10761 1218 10766
rect 1582 10794 1610 11047
rect 1582 10761 1610 10766
rect 1470 10738 1498 10743
rect 1470 10691 1498 10710
rect 1246 10289 1274 10295
rect 1246 10263 1247 10289
rect 1273 10263 1274 10289
rect 1246 10122 1274 10263
rect 1246 10089 1274 10094
rect 2422 10066 2450 13062
rect 2937 12950 3069 12955
rect 2965 12922 2989 12950
rect 3017 12922 3041 12950
rect 2937 12917 3069 12922
rect 7599 12950 7731 12955
rect 7627 12922 7651 12950
rect 7679 12922 7703 12950
rect 7599 12917 7731 12922
rect 5268 12558 5400 12563
rect 5296 12530 5320 12558
rect 5348 12530 5372 12558
rect 5268 12525 5400 12530
rect 8022 12418 8050 12423
rect 2937 12166 3069 12171
rect 2965 12138 2989 12166
rect 3017 12138 3041 12166
rect 2937 12133 3069 12138
rect 7599 12166 7731 12171
rect 7627 12138 7651 12166
rect 7679 12138 7703 12166
rect 7599 12133 7731 12138
rect 8022 12025 8050 12390
rect 8022 11999 8023 12025
rect 8049 11999 8050 12025
rect 8022 11993 8050 11999
rect 8190 11969 8218 11975
rect 8190 11943 8191 11969
rect 8217 11943 8218 11969
rect 8022 11858 8050 11863
rect 5268 11774 5400 11779
rect 5296 11746 5320 11774
rect 5348 11746 5372 11774
rect 5268 11741 5400 11746
rect 2937 11382 3069 11387
rect 2965 11354 2989 11382
rect 3017 11354 3041 11382
rect 2937 11349 3069 11354
rect 7599 11382 7731 11387
rect 7627 11354 7651 11382
rect 7679 11354 7703 11382
rect 7599 11349 7731 11354
rect 8022 11241 8050 11830
rect 8022 11215 8023 11241
rect 8049 11215 8050 11241
rect 8022 11209 8050 11215
rect 7854 11186 7882 11191
rect 8190 11186 8218 11943
rect 8414 11969 8442 14966
rect 8414 11943 8415 11969
rect 8441 11943 8442 11969
rect 8414 11937 8442 11943
rect 5268 10990 5400 10995
rect 5296 10962 5320 10990
rect 5348 10962 5372 10990
rect 5268 10957 5400 10962
rect 2937 10598 3069 10603
rect 2965 10570 2989 10598
rect 3017 10570 3041 10598
rect 2937 10565 3069 10570
rect 7599 10598 7731 10603
rect 7627 10570 7651 10598
rect 7679 10570 7703 10598
rect 7599 10565 7731 10570
rect 7854 10457 7882 11158
rect 7854 10431 7855 10457
rect 7881 10431 7882 10457
rect 7854 10425 7882 10431
rect 8078 11185 8218 11186
rect 8078 11159 8191 11185
rect 8217 11159 8218 11185
rect 8078 11158 8218 11159
rect 8078 10401 8106 11158
rect 8190 11153 8218 11158
rect 8414 11186 8442 11191
rect 8470 11186 8498 15078
rect 8638 12306 8666 18215
rect 8750 17906 8778 19600
rect 9030 18354 9058 18359
rect 9030 18307 9058 18326
rect 9086 18298 9114 19600
rect 9422 18298 9450 19600
rect 9086 18270 9338 18298
rect 8862 17906 8890 17911
rect 8750 17905 8890 17906
rect 8750 17879 8863 17905
rect 8889 17879 8890 17905
rect 8750 17878 8890 17879
rect 8750 17513 8778 17878
rect 8862 17873 8890 17878
rect 9030 17905 9058 17911
rect 9030 17879 9031 17905
rect 9057 17879 9058 17905
rect 9030 17654 9058 17879
rect 8750 17487 8751 17513
rect 8777 17487 8778 17513
rect 8750 17481 8778 17487
rect 8918 17626 9058 17654
rect 8694 15106 8722 15111
rect 8694 12473 8722 15078
rect 8694 12447 8695 12473
rect 8721 12447 8722 12473
rect 8694 12441 8722 12447
rect 8806 12362 8834 12367
rect 8750 12361 8834 12362
rect 8750 12335 8807 12361
rect 8833 12335 8834 12361
rect 8750 12334 8834 12335
rect 8638 12278 8722 12306
rect 8526 11858 8554 11863
rect 8526 11811 8554 11830
rect 8694 11633 8722 12278
rect 8694 11607 8695 11633
rect 8721 11607 8722 11633
rect 8694 11601 8722 11607
rect 8750 11522 8778 12334
rect 8806 12329 8834 12334
rect 8862 11969 8890 11975
rect 8862 11943 8863 11969
rect 8889 11943 8890 11969
rect 8806 11858 8834 11863
rect 8806 11577 8834 11830
rect 8806 11551 8807 11577
rect 8833 11551 8834 11577
rect 8806 11545 8834 11551
rect 8414 11185 8498 11186
rect 8414 11159 8415 11185
rect 8441 11159 8498 11185
rect 8414 11158 8498 11159
rect 8526 11494 8778 11522
rect 8414 11153 8442 11158
rect 8526 11129 8554 11494
rect 8862 11186 8890 11943
rect 8918 11774 8946 17626
rect 9086 17513 9114 18270
rect 9198 17905 9226 17911
rect 9198 17879 9199 17905
rect 9225 17879 9226 17905
rect 9198 17654 9226 17879
rect 9310 17849 9338 18270
rect 9310 17823 9311 17849
rect 9337 17823 9338 17849
rect 9310 17817 9338 17823
rect 9422 18270 9674 18298
rect 9086 17487 9087 17513
rect 9113 17487 9114 17513
rect 9086 17481 9114 17487
rect 9142 17626 9226 17654
rect 9142 14826 9170 17626
rect 9422 17513 9450 18270
rect 9422 17487 9423 17513
rect 9449 17487 9450 17513
rect 9422 17481 9450 17487
rect 9478 17962 9506 17967
rect 9086 14798 9170 14826
rect 9086 11969 9114 14798
rect 9478 13482 9506 17934
rect 9534 17905 9562 17911
rect 9534 17879 9535 17905
rect 9561 17879 9562 17905
rect 9534 13538 9562 17879
rect 9646 17849 9674 18270
rect 9646 17823 9647 17849
rect 9673 17823 9674 17849
rect 9646 17817 9674 17823
rect 9758 17794 9786 19600
rect 9930 18046 10062 18051
rect 9958 18018 9982 18046
rect 10010 18018 10034 18046
rect 9930 18013 10062 18018
rect 9870 17962 9898 17967
rect 9870 17915 9898 17934
rect 10094 17906 10122 19600
rect 10430 18690 10458 19600
rect 10150 18662 10682 18690
rect 10150 18297 10178 18662
rect 10150 18271 10151 18297
rect 10177 18271 10178 18297
rect 10150 18265 10178 18271
rect 10654 18241 10682 18662
rect 10654 18215 10655 18241
rect 10681 18215 10682 18241
rect 10654 18209 10682 18215
rect 10766 18242 10794 19600
rect 10878 18242 10906 18247
rect 10766 18241 10906 18242
rect 10766 18215 10879 18241
rect 10905 18215 10906 18241
rect 10766 18214 10906 18215
rect 10542 18129 10570 18135
rect 10542 18103 10543 18129
rect 10569 18103 10570 18129
rect 10206 17906 10234 17911
rect 10094 17905 10234 17906
rect 10094 17879 10207 17905
rect 10233 17879 10234 17905
rect 10094 17878 10234 17879
rect 9982 17849 10010 17855
rect 9982 17823 9983 17849
rect 10009 17823 10010 17849
rect 9982 17794 10010 17823
rect 9758 17766 10010 17794
rect 9758 17513 9786 17766
rect 9758 17487 9759 17513
rect 9785 17487 9786 17513
rect 9758 17481 9786 17487
rect 10094 17513 10122 17878
rect 10206 17873 10234 17878
rect 10374 17905 10402 17911
rect 10374 17879 10375 17905
rect 10401 17879 10402 17905
rect 10094 17487 10095 17513
rect 10121 17487 10122 17513
rect 10094 17481 10122 17487
rect 9930 17262 10062 17267
rect 9958 17234 9982 17262
rect 10010 17234 10034 17262
rect 9930 17229 10062 17234
rect 9930 16478 10062 16483
rect 9958 16450 9982 16478
rect 10010 16450 10034 16478
rect 9930 16445 10062 16450
rect 9930 15694 10062 15699
rect 9958 15666 9982 15694
rect 10010 15666 10034 15694
rect 9930 15661 10062 15666
rect 9930 14910 10062 14915
rect 9958 14882 9982 14910
rect 10010 14882 10034 14910
rect 9930 14877 10062 14882
rect 10374 14714 10402 17879
rect 10542 17654 10570 18103
rect 10766 17961 10794 18214
rect 10878 18209 10906 18214
rect 11102 18242 11130 19600
rect 12261 18438 12393 18443
rect 12289 18410 12313 18438
rect 12341 18410 12365 18438
rect 12261 18405 12393 18410
rect 16923 18438 17055 18443
rect 16951 18410 16975 18438
rect 17003 18410 17027 18438
rect 16923 18405 17055 18410
rect 11326 18242 11354 18247
rect 11102 18241 11354 18242
rect 11102 18215 11327 18241
rect 11353 18215 11354 18241
rect 11102 18214 11354 18215
rect 10766 17935 10767 17961
rect 10793 17935 10794 17961
rect 10766 17929 10794 17935
rect 11046 18129 11074 18135
rect 11046 18103 11047 18129
rect 11073 18103 11074 18129
rect 10374 14681 10402 14686
rect 10430 17626 10570 17654
rect 9930 14126 10062 14131
rect 9958 14098 9982 14126
rect 10010 14098 10034 14126
rect 9930 14093 10062 14098
rect 9534 13510 9618 13538
rect 9478 13454 9562 13482
rect 9086 11943 9087 11969
rect 9113 11943 9114 11969
rect 9086 11937 9114 11943
rect 9534 11969 9562 13454
rect 9534 11943 9535 11969
rect 9561 11943 9562 11969
rect 9534 11937 9562 11943
rect 8918 11746 9170 11774
rect 8526 11103 8527 11129
rect 8553 11103 8554 11129
rect 8526 11097 8554 11103
rect 8694 11185 8890 11186
rect 8694 11159 8863 11185
rect 8889 11159 8890 11185
rect 8694 11158 8890 11159
rect 8078 10375 8079 10401
rect 8105 10375 8106 10401
rect 7742 10346 7770 10351
rect 7742 10299 7770 10318
rect 5268 10206 5400 10211
rect 5296 10178 5320 10206
rect 5348 10178 5372 10206
rect 5268 10173 5400 10178
rect 8078 10094 8106 10375
rect 8246 10850 8274 10855
rect 8246 10401 8274 10822
rect 8694 10402 8722 11158
rect 8862 11153 8890 11158
rect 9142 11185 9170 11746
rect 9142 11159 9143 11185
rect 9169 11159 9170 11185
rect 9142 11153 9170 11159
rect 9590 11185 9618 13510
rect 9930 13342 10062 13347
rect 9958 13314 9982 13342
rect 10010 13314 10034 13342
rect 9930 13309 10062 13314
rect 9930 12558 10062 12563
rect 9958 12530 9982 12558
rect 10010 12530 10034 12558
rect 9930 12525 10062 12530
rect 9930 11774 10062 11779
rect 9958 11746 9982 11774
rect 10010 11746 10034 11774
rect 10430 11774 10458 17626
rect 10598 14714 10626 14719
rect 10430 11746 10514 11774
rect 9930 11741 10062 11746
rect 9590 11159 9591 11185
rect 9617 11159 9618 11185
rect 9590 11153 9618 11159
rect 8246 10375 8247 10401
rect 8273 10375 8274 10401
rect 8246 10369 8274 10375
rect 8638 10401 8722 10402
rect 8638 10375 8695 10401
rect 8721 10375 8722 10401
rect 8638 10374 8722 10375
rect 2422 10033 2450 10038
rect 8022 10066 8106 10094
rect 8358 10289 8386 10295
rect 8358 10263 8359 10289
rect 8385 10263 8386 10289
rect 8246 10066 8274 10071
rect 2142 10010 2170 10015
rect 2142 9963 2170 9982
rect 2937 9814 3069 9819
rect 2965 9786 2989 9814
rect 3017 9786 3041 9814
rect 2937 9781 3069 9786
rect 7599 9814 7731 9819
rect 7627 9786 7651 9814
rect 7679 9786 7703 9814
rect 7599 9781 7731 9786
rect 8022 9617 8050 10066
rect 8246 10019 8274 10038
rect 8358 10009 8386 10263
rect 8358 9983 8359 10009
rect 8385 9983 8386 10009
rect 8358 9977 8386 9983
rect 8638 9730 8666 10374
rect 8694 10369 8722 10374
rect 8862 11074 8890 11079
rect 8862 10401 8890 11046
rect 9930 10990 10062 10995
rect 9958 10962 9982 10990
rect 10010 10962 10034 10990
rect 9930 10957 10062 10962
rect 10486 10849 10514 11746
rect 10486 10823 10487 10849
rect 10513 10823 10514 10849
rect 10486 10817 10514 10823
rect 10598 10458 10626 14686
rect 11046 13454 11074 18103
rect 11102 17961 11130 18214
rect 11326 18209 11354 18214
rect 11102 17935 11103 17961
rect 11129 17935 11130 17961
rect 11102 17929 11130 17935
rect 11214 18129 11242 18135
rect 11214 18103 11215 18129
rect 11241 18103 11242 18129
rect 11214 13454 11242 18103
rect 14592 18046 14724 18051
rect 14620 18018 14644 18046
rect 14672 18018 14696 18046
rect 14592 18013 14724 18018
rect 19254 18046 19386 18051
rect 19282 18018 19306 18046
rect 19334 18018 19358 18046
rect 19254 18013 19386 18018
rect 12261 17654 12393 17659
rect 12289 17626 12313 17654
rect 12341 17626 12365 17654
rect 12261 17621 12393 17626
rect 16923 17654 17055 17659
rect 16951 17626 16975 17654
rect 17003 17626 17027 17654
rect 16923 17621 17055 17626
rect 14592 17262 14724 17267
rect 14620 17234 14644 17262
rect 14672 17234 14696 17262
rect 14592 17229 14724 17234
rect 19254 17262 19386 17267
rect 19282 17234 19306 17262
rect 19334 17234 19358 17262
rect 19254 17229 19386 17234
rect 12261 16870 12393 16875
rect 12289 16842 12313 16870
rect 12341 16842 12365 16870
rect 12261 16837 12393 16842
rect 16923 16870 17055 16875
rect 16951 16842 16975 16870
rect 17003 16842 17027 16870
rect 16923 16837 17055 16842
rect 14592 16478 14724 16483
rect 14620 16450 14644 16478
rect 14672 16450 14696 16478
rect 14592 16445 14724 16450
rect 19254 16478 19386 16483
rect 19282 16450 19306 16478
rect 19334 16450 19358 16478
rect 19254 16445 19386 16450
rect 12261 16086 12393 16091
rect 12289 16058 12313 16086
rect 12341 16058 12365 16086
rect 12261 16053 12393 16058
rect 16923 16086 17055 16091
rect 16951 16058 16975 16086
rect 17003 16058 17027 16086
rect 16923 16053 17055 16058
rect 14592 15694 14724 15699
rect 14620 15666 14644 15694
rect 14672 15666 14696 15694
rect 14592 15661 14724 15666
rect 19254 15694 19386 15699
rect 19282 15666 19306 15694
rect 19334 15666 19358 15694
rect 19254 15661 19386 15666
rect 12261 15302 12393 15307
rect 12289 15274 12313 15302
rect 12341 15274 12365 15302
rect 12261 15269 12393 15274
rect 16923 15302 17055 15307
rect 16951 15274 16975 15302
rect 17003 15274 17027 15302
rect 16923 15269 17055 15274
rect 14592 14910 14724 14915
rect 14620 14882 14644 14910
rect 14672 14882 14696 14910
rect 14592 14877 14724 14882
rect 19254 14910 19386 14915
rect 19282 14882 19306 14910
rect 19334 14882 19358 14910
rect 19254 14877 19386 14882
rect 12261 14518 12393 14523
rect 12289 14490 12313 14518
rect 12341 14490 12365 14518
rect 12261 14485 12393 14490
rect 16923 14518 17055 14523
rect 16951 14490 16975 14518
rect 17003 14490 17027 14518
rect 16923 14485 17055 14490
rect 14592 14126 14724 14131
rect 14620 14098 14644 14126
rect 14672 14098 14696 14126
rect 14592 14093 14724 14098
rect 19254 14126 19386 14131
rect 19282 14098 19306 14126
rect 19334 14098 19358 14126
rect 19254 14093 19386 14098
rect 12261 13734 12393 13739
rect 12289 13706 12313 13734
rect 12341 13706 12365 13734
rect 12261 13701 12393 13706
rect 16923 13734 17055 13739
rect 16951 13706 16975 13734
rect 17003 13706 17027 13734
rect 16923 13701 17055 13706
rect 11046 13426 11130 13454
rect 10710 11073 10738 11079
rect 10710 11047 10711 11073
rect 10737 11047 10738 11073
rect 10710 10906 10738 11047
rect 10878 11074 10906 11079
rect 11046 11074 11074 11079
rect 10878 11027 10906 11046
rect 10990 11073 11074 11074
rect 10990 11047 11047 11073
rect 11073 11047 11074 11073
rect 10990 11046 11074 11047
rect 10710 10873 10738 10878
rect 10990 10905 11018 11046
rect 11046 11041 11074 11046
rect 10990 10879 10991 10905
rect 11017 10879 11018 10905
rect 10990 10873 11018 10879
rect 10710 10794 10738 10799
rect 10934 10794 10962 10799
rect 10710 10793 10850 10794
rect 10710 10767 10711 10793
rect 10737 10767 10850 10793
rect 10710 10766 10850 10767
rect 10710 10761 10738 10766
rect 10654 10458 10682 10463
rect 10598 10457 10682 10458
rect 10598 10431 10655 10457
rect 10681 10431 10682 10457
rect 10598 10430 10682 10431
rect 10654 10425 10682 10430
rect 8862 10375 8863 10401
rect 8889 10375 8890 10401
rect 8862 10369 8890 10375
rect 9422 10401 9450 10407
rect 9422 10375 9423 10401
rect 9449 10375 9450 10401
rect 9422 10346 9450 10375
rect 9422 10313 9450 10318
rect 10822 10401 10850 10766
rect 10934 10747 10962 10766
rect 10822 10375 10823 10401
rect 10849 10375 10850 10401
rect 8862 10290 8890 10295
rect 8862 10094 8890 10262
rect 9930 10206 10062 10211
rect 9958 10178 9982 10206
rect 10010 10178 10034 10206
rect 9930 10173 10062 10178
rect 8694 10066 8722 10071
rect 8862 10066 9002 10094
rect 8694 10019 8722 10038
rect 8806 10009 8834 10015
rect 8806 9983 8807 10009
rect 8833 9983 8834 10009
rect 8638 9702 8722 9730
rect 8022 9591 8023 9617
rect 8049 9591 8050 9617
rect 1134 9529 1162 9534
rect 7742 9562 7770 9567
rect 7854 9562 7882 9567
rect 7770 9561 7882 9562
rect 7770 9535 7855 9561
rect 7881 9535 7882 9561
rect 7770 9534 7882 9535
rect 7742 9515 7770 9534
rect 7854 9529 7882 9534
rect 1022 9506 1050 9511
rect 1022 9459 1050 9478
rect 1246 9505 1274 9511
rect 1246 9479 1247 9505
rect 1273 9479 1274 9505
rect 854 9417 882 9422
rect 1246 9450 1274 9479
rect 1246 9417 1274 9422
rect 5268 9422 5400 9427
rect 5296 9394 5320 9422
rect 5348 9394 5372 9422
rect 5268 9389 5400 9394
rect 1022 9281 1050 9287
rect 1022 9255 1023 9281
rect 1049 9255 1050 9281
rect 854 9225 882 9231
rect 854 9199 855 9225
rect 881 9199 882 9225
rect 854 9114 882 9199
rect 1022 9226 1050 9255
rect 1022 9193 1050 9198
rect 8022 9226 8050 9591
rect 8246 9618 8274 9623
rect 8246 9571 8274 9590
rect 8694 9617 8722 9702
rect 8694 9591 8695 9617
rect 8721 9591 8722 9617
rect 8358 9562 8386 9567
rect 8358 9515 8386 9534
rect 8694 9338 8722 9591
rect 8806 9562 8834 9983
rect 8974 9617 9002 10066
rect 9534 9953 9562 9959
rect 9534 9927 9535 9953
rect 9561 9927 9562 9953
rect 8974 9591 8975 9617
rect 9001 9591 9002 9617
rect 8974 9585 9002 9591
rect 9366 9617 9394 9623
rect 9366 9591 9367 9617
rect 9393 9591 9394 9617
rect 8806 9529 8834 9534
rect 9310 9506 9338 9511
rect 9142 9338 9170 9343
rect 8694 9337 9170 9338
rect 8694 9311 9143 9337
rect 9169 9311 9170 9337
rect 8694 9310 9170 9311
rect 9142 9305 9170 9310
rect 9198 9282 9226 9287
rect 8022 9193 8050 9198
rect 8694 9226 8722 9231
rect 8694 9179 8722 9198
rect 8918 9225 8946 9231
rect 8918 9199 8919 9225
rect 8945 9199 8946 9225
rect 854 9081 882 9086
rect 1246 9169 1274 9175
rect 1246 9143 1247 9169
rect 1273 9143 1274 9169
rect 1246 9114 1274 9143
rect 1246 9081 1274 9086
rect 8414 9169 8442 9175
rect 8414 9143 8415 9169
rect 8441 9143 8442 9169
rect 2937 9030 3069 9035
rect 2965 9002 2989 9030
rect 3017 9002 3041 9030
rect 2937 8997 3069 9002
rect 7599 9030 7731 9035
rect 7627 9002 7651 9030
rect 7679 9002 7703 9030
rect 7599 8997 7731 9002
rect 966 8889 994 8895
rect 966 8863 967 8889
rect 993 8863 994 8889
rect 854 8778 882 8783
rect 854 8553 882 8750
rect 854 8527 855 8553
rect 881 8527 882 8553
rect 854 8521 882 8527
rect 966 8442 994 8863
rect 2142 8833 2170 8839
rect 2142 8807 2143 8833
rect 2169 8807 2170 8833
rect 1246 8778 1274 8783
rect 966 8409 994 8414
rect 1022 8497 1050 8503
rect 1022 8471 1023 8497
rect 1049 8471 1050 8497
rect 1022 8330 1050 8471
rect 1022 8297 1050 8302
rect 1190 8441 1218 8447
rect 1190 8415 1191 8441
rect 1217 8415 1218 8441
rect 1190 8386 1218 8415
rect 1190 8106 1218 8358
rect 1190 8073 1218 8078
rect 1246 8105 1274 8750
rect 1246 8079 1247 8105
rect 1273 8079 1274 8105
rect 1246 8073 1274 8079
rect 1358 8497 1386 8503
rect 1358 8471 1359 8497
rect 1385 8471 1386 8497
rect 910 8049 938 8055
rect 910 8023 911 8049
rect 937 8023 938 8049
rect 910 7770 938 8023
rect 1358 8050 1386 8471
rect 1582 8441 1610 8447
rect 1582 8415 1583 8441
rect 1609 8415 1610 8441
rect 1582 8386 1610 8415
rect 1582 8353 1610 8358
rect 2142 8162 2170 8807
rect 8414 8722 8442 9143
rect 8918 9114 8946 9199
rect 9198 9114 9226 9254
rect 8806 9086 9226 9114
rect 9310 9225 9338 9478
rect 9310 9199 9311 9225
rect 9337 9199 9338 9225
rect 8638 8722 8666 8727
rect 8806 8722 8834 9086
rect 8414 8721 8834 8722
rect 8414 8695 8639 8721
rect 8665 8695 8834 8721
rect 8414 8694 8834 8695
rect 8862 8889 8890 8895
rect 8862 8863 8863 8889
rect 8889 8863 8890 8889
rect 5268 8638 5400 8643
rect 5296 8610 5320 8638
rect 5348 8610 5372 8638
rect 5268 8605 5400 8610
rect 7966 8497 7994 8503
rect 7966 8471 7967 8497
rect 7993 8471 7994 8497
rect 2937 8246 3069 8251
rect 2965 8218 2989 8246
rect 3017 8218 3041 8246
rect 2937 8213 3069 8218
rect 7599 8246 7731 8251
rect 7627 8218 7651 8246
rect 7679 8218 7703 8246
rect 7599 8213 7731 8218
rect 2142 8129 2170 8134
rect 7966 8162 7994 8471
rect 7966 8129 7994 8134
rect 8078 8441 8106 8447
rect 8078 8415 8079 8441
rect 8105 8415 8106 8441
rect 1358 8017 1386 8022
rect 7742 8049 7770 8055
rect 7742 8023 7743 8049
rect 7769 8023 7770 8049
rect 7574 7994 7602 7999
rect 7574 7947 7602 7966
rect 7686 7994 7714 7999
rect 1022 7938 1050 7943
rect 1022 7891 1050 7910
rect 5268 7854 5400 7859
rect 5296 7826 5320 7854
rect 5348 7826 5372 7854
rect 5268 7821 5400 7826
rect 910 7723 938 7742
rect 7686 7713 7714 7966
rect 7686 7687 7687 7713
rect 7713 7687 7714 7713
rect 7686 7681 7714 7687
rect 7742 7714 7770 8023
rect 7966 8050 7994 8055
rect 7966 8003 7994 8022
rect 8078 7993 8106 8415
rect 8638 8330 8666 8694
rect 8638 8297 8666 8302
rect 8582 8050 8610 8055
rect 8470 8049 8610 8050
rect 8470 8023 8583 8049
rect 8609 8023 8610 8049
rect 8470 8022 8610 8023
rect 8078 7967 8079 7993
rect 8105 7967 8106 7993
rect 8078 7961 8106 7967
rect 8302 7994 8330 7999
rect 8302 7947 8330 7966
rect 7910 7770 7938 7775
rect 7910 7769 8162 7770
rect 7910 7743 7911 7769
rect 7937 7743 8162 7769
rect 7910 7742 8162 7743
rect 7910 7737 7938 7742
rect 7742 7681 7770 7686
rect 6902 7657 6930 7663
rect 6902 7631 6903 7657
rect 6929 7631 6930 7657
rect 2937 7462 3069 7467
rect 2965 7434 2989 7462
rect 3017 7434 3041 7462
rect 2937 7429 3069 7434
rect 5268 7070 5400 7075
rect 5296 7042 5320 7070
rect 5348 7042 5372 7070
rect 5268 7037 5400 7042
rect 2937 6678 3069 6683
rect 2965 6650 2989 6678
rect 3017 6650 3041 6678
rect 2937 6645 3069 6650
rect 5268 6286 5400 6291
rect 5296 6258 5320 6286
rect 5348 6258 5372 6286
rect 5268 6253 5400 6258
rect 2937 5894 3069 5899
rect 2965 5866 2989 5894
rect 3017 5866 3041 5894
rect 2937 5861 3069 5866
rect 5268 5502 5400 5507
rect 5296 5474 5320 5502
rect 5348 5474 5372 5502
rect 5268 5469 5400 5474
rect 2937 5110 3069 5115
rect 2965 5082 2989 5110
rect 3017 5082 3041 5110
rect 2937 5077 3069 5082
rect 5268 4718 5400 4723
rect 5296 4690 5320 4718
rect 5348 4690 5372 4718
rect 5268 4685 5400 4690
rect 2937 4326 3069 4331
rect 2965 4298 2989 4326
rect 3017 4298 3041 4326
rect 2937 4293 3069 4298
rect 6902 4214 6930 7631
rect 7294 7657 7322 7663
rect 7294 7631 7295 7657
rect 7321 7631 7322 7657
rect 6902 4186 7042 4214
rect 5268 3934 5400 3939
rect 5296 3906 5320 3934
rect 5348 3906 5372 3934
rect 5268 3901 5400 3906
rect 2937 3542 3069 3547
rect 2965 3514 2989 3542
rect 3017 3514 3041 3542
rect 2937 3509 3069 3514
rect 5268 3150 5400 3155
rect 5296 3122 5320 3150
rect 5348 3122 5372 3150
rect 5268 3117 5400 3122
rect 2937 2758 3069 2763
rect 2965 2730 2989 2758
rect 3017 2730 3041 2758
rect 2937 2725 3069 2730
rect 5268 2366 5400 2371
rect 5296 2338 5320 2366
rect 5348 2338 5372 2366
rect 5268 2333 5400 2338
rect 6734 2282 6762 2287
rect 6734 2281 6930 2282
rect 6734 2255 6735 2281
rect 6761 2255 6930 2281
rect 6734 2254 6930 2255
rect 6734 2249 6762 2254
rect 6846 2169 6874 2175
rect 6846 2143 6847 2169
rect 6873 2143 6874 2169
rect 6510 2114 6538 2119
rect 6510 2067 6538 2086
rect 6846 2114 6874 2143
rect 6902 2170 6930 2254
rect 7014 2281 7042 4186
rect 7014 2255 7015 2281
rect 7041 2255 7042 2281
rect 7014 2249 7042 2255
rect 7294 2282 7322 7631
rect 8022 7657 8050 7663
rect 8022 7631 8023 7657
rect 8049 7631 8050 7657
rect 7599 7462 7731 7467
rect 7627 7434 7651 7462
rect 7679 7434 7703 7462
rect 7599 7429 7731 7434
rect 7294 2249 7322 2254
rect 7350 7210 7378 7215
rect 7350 2281 7378 7182
rect 7599 6678 7731 6683
rect 7627 6650 7651 6678
rect 7679 6650 7703 6678
rect 7599 6645 7731 6650
rect 7854 6034 7882 6039
rect 7798 6006 7854 6034
rect 7599 5894 7731 5899
rect 7627 5866 7651 5894
rect 7679 5866 7703 5894
rect 7599 5861 7731 5866
rect 7599 5110 7731 5115
rect 7627 5082 7651 5110
rect 7679 5082 7703 5110
rect 7599 5077 7731 5082
rect 7599 4326 7731 4331
rect 7627 4298 7651 4326
rect 7679 4298 7703 4326
rect 7599 4293 7731 4298
rect 7599 3542 7731 3547
rect 7627 3514 7651 3542
rect 7679 3514 7703 3542
rect 7599 3509 7731 3514
rect 7599 2758 7731 2763
rect 7627 2730 7651 2758
rect 7679 2730 7703 2758
rect 7599 2725 7731 2730
rect 7798 2674 7826 6006
rect 7854 6001 7882 6006
rect 7686 2646 7826 2674
rect 7350 2255 7351 2281
rect 7377 2255 7378 2281
rect 7350 2249 7378 2255
rect 7406 2561 7434 2567
rect 7406 2535 7407 2561
rect 7433 2535 7434 2561
rect 7182 2170 7210 2175
rect 6902 2169 7210 2170
rect 6902 2143 7183 2169
rect 7209 2143 7210 2169
rect 6902 2142 7210 2143
rect 7406 2170 7434 2535
rect 7686 2281 7714 2646
rect 7742 2450 7770 2455
rect 7742 2449 7882 2450
rect 7742 2423 7743 2449
rect 7769 2423 7882 2449
rect 7742 2422 7882 2423
rect 7742 2417 7770 2422
rect 7686 2255 7687 2281
rect 7713 2255 7714 2281
rect 7686 2249 7714 2255
rect 7854 2225 7882 2422
rect 8022 2281 8050 7631
rect 8134 7574 8162 7742
rect 8246 7714 8274 7719
rect 8246 7657 8274 7686
rect 8246 7631 8247 7657
rect 8273 7631 8274 7657
rect 8246 7625 8274 7631
rect 8414 7601 8442 7607
rect 8414 7575 8415 7601
rect 8441 7575 8442 7601
rect 8134 7546 8218 7574
rect 8190 7265 8218 7546
rect 8190 7239 8191 7265
rect 8217 7239 8218 7265
rect 8190 7233 8218 7239
rect 8078 7154 8106 7159
rect 8078 7153 8162 7154
rect 8078 7127 8079 7153
rect 8105 7127 8162 7153
rect 8078 7126 8162 7127
rect 8078 7121 8106 7126
rect 8022 2255 8023 2281
rect 8049 2255 8050 2281
rect 8022 2249 8050 2255
rect 8078 2449 8106 2455
rect 8078 2423 8079 2449
rect 8105 2423 8106 2449
rect 7854 2199 7855 2225
rect 7881 2199 7882 2225
rect 7574 2170 7602 2175
rect 7406 2169 7602 2170
rect 7406 2143 7575 2169
rect 7601 2143 7602 2169
rect 7406 2142 7602 2143
rect 2937 1974 3069 1979
rect 2965 1946 2989 1974
rect 3017 1946 3041 1974
rect 2937 1941 3069 1946
rect 6678 1834 6706 1839
rect 6398 1833 6706 1834
rect 6398 1807 6679 1833
rect 6705 1807 6706 1833
rect 6398 1806 6706 1807
rect 5268 1582 5400 1587
rect 5296 1554 5320 1582
rect 5348 1554 5372 1582
rect 5268 1549 5400 1554
rect 6398 400 6426 1806
rect 6678 1801 6706 1806
rect 6846 1442 6874 2086
rect 7182 1778 7210 2142
rect 6734 1414 6874 1442
rect 7070 1750 7210 1778
rect 6734 400 6762 1414
rect 7070 400 7098 1750
rect 7518 1554 7546 2142
rect 7574 2137 7602 2142
rect 7599 1974 7731 1979
rect 7627 1946 7651 1974
rect 7679 1946 7703 1974
rect 7599 1941 7731 1946
rect 7798 1778 7826 1797
rect 7798 1745 7826 1750
rect 7854 1694 7882 2199
rect 7406 1526 7546 1554
rect 7742 1666 7882 1694
rect 8022 1722 8050 1741
rect 8022 1689 8050 1694
rect 8078 1694 8106 2423
rect 8134 1778 8162 7126
rect 8414 6034 8442 7575
rect 8414 6001 8442 6006
rect 8470 5922 8498 8022
rect 8582 8017 8610 8022
rect 8862 7714 8890 8863
rect 9030 8833 9058 9086
rect 9030 8807 9031 8833
rect 9057 8807 9058 8833
rect 9030 8801 9058 8807
rect 9310 8834 9338 9199
rect 9366 9226 9394 9591
rect 9534 9506 9562 9927
rect 9926 9674 9954 9679
rect 9926 9627 9954 9646
rect 10822 9674 10850 10375
rect 11046 10402 11074 10407
rect 11102 10402 11130 13426
rect 11158 13426 11242 13454
rect 11158 10794 11186 13426
rect 14592 13342 14724 13347
rect 14620 13314 14644 13342
rect 14672 13314 14696 13342
rect 14592 13309 14724 13314
rect 19254 13342 19386 13347
rect 19282 13314 19306 13342
rect 19334 13314 19358 13342
rect 19254 13309 19386 13314
rect 12261 12950 12393 12955
rect 12289 12922 12313 12950
rect 12341 12922 12365 12950
rect 12261 12917 12393 12922
rect 16923 12950 17055 12955
rect 16951 12922 16975 12950
rect 17003 12922 17027 12950
rect 16923 12917 17055 12922
rect 14592 12558 14724 12563
rect 14620 12530 14644 12558
rect 14672 12530 14696 12558
rect 14592 12525 14724 12530
rect 19254 12558 19386 12563
rect 19282 12530 19306 12558
rect 19334 12530 19358 12558
rect 19254 12525 19386 12530
rect 11214 12362 11242 12367
rect 11214 11129 11242 12334
rect 17822 12362 17850 12367
rect 17822 12315 17850 12334
rect 18998 12249 19026 12255
rect 18998 12223 18999 12249
rect 19025 12223 19026 12249
rect 12261 12166 12393 12171
rect 12289 12138 12313 12166
rect 12341 12138 12365 12166
rect 12261 12133 12393 12138
rect 16923 12166 17055 12171
rect 16951 12138 16975 12166
rect 17003 12138 17027 12166
rect 16923 12133 17055 12138
rect 18998 12138 19026 12223
rect 18998 12105 19026 12110
rect 19110 11913 19138 11919
rect 19110 11887 19111 11913
rect 19137 11887 19138 11913
rect 18830 11858 18858 11863
rect 18942 11858 18970 11863
rect 18830 11811 18858 11830
rect 18886 11857 18970 11858
rect 18886 11831 18943 11857
rect 18969 11831 18970 11857
rect 18886 11830 18970 11831
rect 14592 11774 14724 11779
rect 14620 11746 14644 11774
rect 14672 11746 14696 11774
rect 14592 11741 14724 11746
rect 11214 11103 11215 11129
rect 11241 11103 11242 11129
rect 11214 11097 11242 11103
rect 12054 11634 12082 11639
rect 11158 10761 11186 10766
rect 11214 10906 11242 10911
rect 11046 10401 11130 10402
rect 11046 10375 11047 10401
rect 11073 10375 11130 10401
rect 11046 10374 11130 10375
rect 11046 10369 11074 10374
rect 11158 10346 11186 10351
rect 11214 10346 11242 10878
rect 11158 10345 11242 10346
rect 11158 10319 11159 10345
rect 11185 10319 11242 10345
rect 11158 10318 11242 10319
rect 11326 10793 11354 10799
rect 11326 10767 11327 10793
rect 11353 10767 11354 10793
rect 11326 10402 11354 10767
rect 11606 10794 11634 10799
rect 11606 10747 11634 10766
rect 12054 10793 12082 11606
rect 18830 11521 18858 11527
rect 18830 11495 18831 11521
rect 18857 11495 18858 11521
rect 18830 11466 18858 11495
rect 18830 11433 18858 11438
rect 12261 11382 12393 11387
rect 12289 11354 12313 11382
rect 12341 11354 12365 11382
rect 12261 11349 12393 11354
rect 16923 11382 17055 11387
rect 16951 11354 16975 11382
rect 17003 11354 17027 11382
rect 16923 11349 17055 11354
rect 18830 11130 18858 11135
rect 18830 11083 18858 11102
rect 17822 11074 17850 11079
rect 14592 10990 14724 10995
rect 14620 10962 14644 10990
rect 14672 10962 14696 10990
rect 14592 10957 14724 10962
rect 12054 10767 12055 10793
rect 12081 10767 12082 10793
rect 12054 10761 12082 10767
rect 17822 10793 17850 11046
rect 17822 10767 17823 10793
rect 17849 10767 17850 10793
rect 17822 10761 17850 10767
rect 12261 10598 12393 10603
rect 12289 10570 12313 10598
rect 12341 10570 12365 10598
rect 12261 10565 12393 10570
rect 16923 10598 17055 10603
rect 16951 10570 16975 10598
rect 17003 10570 17027 10598
rect 16923 10565 17055 10570
rect 18270 10458 18298 10463
rect 18270 10411 18298 10430
rect 11382 10402 11410 10407
rect 11326 10401 11410 10402
rect 11326 10375 11383 10401
rect 11409 10375 11410 10401
rect 11326 10374 11410 10375
rect 11158 10313 11186 10318
rect 11326 10094 11354 10374
rect 11382 10369 11410 10374
rect 11718 10402 11746 10407
rect 11718 10355 11746 10374
rect 12222 10401 12250 10407
rect 12222 10375 12223 10401
rect 12249 10375 12250 10401
rect 12222 10346 12250 10375
rect 18886 10402 18914 11830
rect 18942 11825 18970 11830
rect 19110 11858 19138 11887
rect 19110 11825 19138 11830
rect 19254 11774 19386 11779
rect 19282 11746 19306 11774
rect 19334 11746 19358 11774
rect 19254 11741 19386 11746
rect 18942 11634 18970 11639
rect 18942 11587 18970 11606
rect 19110 11577 19138 11583
rect 19110 11551 19111 11577
rect 19137 11551 19138 11577
rect 19110 11466 19138 11551
rect 19110 11433 19138 11438
rect 19110 11130 19138 11135
rect 19110 11083 19138 11102
rect 18942 11073 18970 11079
rect 18942 11047 18943 11073
rect 18969 11047 18970 11073
rect 18942 10906 18970 11047
rect 19254 10990 19386 10995
rect 19282 10962 19306 10990
rect 19334 10962 19358 10990
rect 19254 10957 19386 10962
rect 18942 10873 18970 10878
rect 18998 10794 19026 10799
rect 18998 10737 19026 10766
rect 18998 10711 18999 10737
rect 19025 10711 19026 10737
rect 18998 10705 19026 10711
rect 18886 10369 18914 10374
rect 19110 10458 19138 10463
rect 19110 10401 19138 10430
rect 19110 10375 19111 10401
rect 19137 10375 19138 10401
rect 19110 10369 19138 10375
rect 12222 10313 12250 10318
rect 18774 10346 18802 10351
rect 18942 10346 18970 10351
rect 18774 10345 18858 10346
rect 18774 10319 18775 10345
rect 18801 10319 18858 10345
rect 18774 10318 18858 10319
rect 18774 10313 18802 10318
rect 18606 10289 18634 10295
rect 18606 10263 18607 10289
rect 18633 10263 18634 10289
rect 14592 10206 14724 10211
rect 14620 10178 14644 10206
rect 14672 10178 14696 10206
rect 14592 10173 14724 10178
rect 18606 10094 18634 10263
rect 9646 9506 9674 9511
rect 9534 9505 9674 9506
rect 9534 9479 9647 9505
rect 9673 9479 9674 9505
rect 9534 9478 9674 9479
rect 9646 9282 9674 9478
rect 10094 9506 10122 9511
rect 10094 9459 10122 9478
rect 10262 9506 10290 9511
rect 10262 9459 10290 9478
rect 9930 9422 10062 9427
rect 9958 9394 9982 9422
rect 10010 9394 10034 9422
rect 9930 9389 10062 9394
rect 9646 9249 9674 9254
rect 9366 9193 9394 9198
rect 10822 9225 10850 9646
rect 11270 10066 11354 10094
rect 18550 10066 18634 10094
rect 18830 10122 18858 10318
rect 18942 10299 18970 10318
rect 19254 10206 19386 10211
rect 19282 10178 19306 10206
rect 19334 10178 19358 10206
rect 19254 10173 19386 10178
rect 18830 10089 18858 10094
rect 18942 10066 18970 10071
rect 11158 9506 11186 9511
rect 11102 9505 11186 9506
rect 11102 9479 11159 9505
rect 11185 9479 11186 9505
rect 11102 9478 11186 9479
rect 11102 9337 11130 9478
rect 11158 9473 11186 9478
rect 11270 9506 11298 10066
rect 12261 9814 12393 9819
rect 12289 9786 12313 9814
rect 12341 9786 12365 9814
rect 12261 9781 12393 9786
rect 16923 9814 17055 9819
rect 16951 9786 16975 9814
rect 17003 9786 17027 9814
rect 16923 9781 17055 9786
rect 11102 9311 11103 9337
rect 11129 9311 11130 9337
rect 11102 9305 11130 9311
rect 10822 9199 10823 9225
rect 10849 9199 10850 9225
rect 10598 9170 10626 9175
rect 10598 9123 10626 9142
rect 9590 8834 9618 8839
rect 9310 8833 9618 8834
rect 9310 8807 9591 8833
rect 9617 8807 9618 8833
rect 9310 8806 9618 8807
rect 9086 8050 9114 8055
rect 8862 7574 8890 7686
rect 8974 8049 9114 8050
rect 8974 8023 9087 8049
rect 9113 8023 9114 8049
rect 8974 8022 9114 8023
rect 8862 7546 8946 7574
rect 8918 7265 8946 7546
rect 8918 7239 8919 7265
rect 8945 7239 8946 7265
rect 8918 7233 8946 7239
rect 8750 7210 8778 7215
rect 8750 7163 8778 7182
rect 8358 5894 8498 5922
rect 8358 4634 8386 5894
rect 8974 5194 9002 8022
rect 9086 8017 9114 8022
rect 9254 7938 9282 7943
rect 9142 7602 9170 7607
rect 8246 4606 8386 4634
rect 8806 5166 9002 5194
rect 9086 7601 9170 7602
rect 9086 7575 9143 7601
rect 9169 7575 9170 7601
rect 9086 7574 9170 7575
rect 8190 2282 8218 2287
rect 8190 2235 8218 2254
rect 8134 1745 8162 1750
rect 8190 1722 8218 1727
rect 8246 1722 8274 4606
rect 8358 2449 8386 2455
rect 8358 2423 8359 2449
rect 8385 2423 8386 2449
rect 8190 1721 8274 1722
rect 8190 1695 8191 1721
rect 8217 1695 8274 1721
rect 8190 1694 8274 1695
rect 8302 2169 8330 2175
rect 8302 2143 8303 2169
rect 8329 2143 8330 2169
rect 8078 1666 8162 1694
rect 8190 1689 8218 1694
rect 7406 400 7434 1526
rect 7742 400 7770 1666
rect 8134 1554 8162 1666
rect 8302 1554 8330 2143
rect 8358 1722 8386 2423
rect 8638 1777 8666 1783
rect 8638 1751 8639 1777
rect 8665 1751 8666 1777
rect 8358 1666 8442 1694
rect 8078 1526 8330 1554
rect 8078 400 8106 1526
rect 8414 400 8442 1666
rect 8638 1274 8666 1751
rect 8750 1722 8778 1727
rect 8806 1722 8834 5166
rect 8750 1721 8834 1722
rect 8750 1695 8751 1721
rect 8777 1695 8834 1721
rect 8750 1694 8834 1695
rect 8862 2113 8890 2119
rect 8862 2087 8863 2113
rect 8889 2087 8890 2113
rect 8750 1689 8778 1694
rect 8862 1274 8890 2087
rect 8638 1246 8890 1274
rect 8974 1777 9002 1783
rect 8974 1751 8975 1777
rect 9001 1751 9002 1777
rect 8974 1274 9002 1751
rect 9086 1721 9114 7574
rect 9142 7569 9170 7574
rect 9198 7265 9226 7271
rect 9198 7239 9199 7265
rect 9225 7239 9226 7265
rect 9198 5922 9226 7239
rect 9254 7209 9282 7910
rect 9310 7714 9338 7719
rect 9310 7657 9338 7686
rect 9310 7631 9311 7657
rect 9337 7631 9338 7657
rect 9310 7625 9338 7631
rect 9254 7183 9255 7209
rect 9281 7183 9282 7209
rect 9254 7177 9282 7183
rect 9198 5894 9282 5922
rect 9086 1695 9087 1721
rect 9113 1695 9114 1721
rect 9086 1689 9114 1695
rect 9198 2113 9226 2119
rect 9198 2087 9199 2113
rect 9225 2087 9226 2113
rect 9198 1274 9226 2087
rect 9254 1721 9282 5894
rect 9422 2282 9450 8806
rect 9590 8801 9618 8806
rect 10822 8833 10850 9199
rect 11046 9225 11074 9231
rect 11046 9199 11047 9225
rect 11073 9199 11074 9225
rect 11046 8946 11074 9199
rect 11270 9226 11298 9478
rect 11326 9590 11578 9618
rect 11326 9505 11354 9590
rect 11326 9479 11327 9505
rect 11353 9479 11354 9505
rect 11326 9473 11354 9479
rect 11494 9505 11522 9511
rect 11494 9479 11495 9505
rect 11521 9479 11522 9505
rect 11326 9226 11354 9231
rect 11270 9225 11466 9226
rect 11270 9199 11327 9225
rect 11353 9199 11466 9225
rect 11270 9198 11466 9199
rect 11326 9193 11354 9198
rect 11046 8913 11074 8918
rect 10822 8807 10823 8833
rect 10849 8807 10850 8833
rect 10822 8801 10850 8807
rect 11102 8833 11130 8839
rect 11102 8807 11103 8833
rect 11129 8807 11130 8833
rect 10654 8778 10682 8783
rect 10654 8731 10682 8750
rect 9478 8721 9506 8727
rect 9478 8695 9479 8721
rect 9505 8695 9506 8721
rect 9478 7994 9506 8695
rect 9930 8638 10062 8643
rect 9958 8610 9982 8638
rect 10010 8610 10034 8638
rect 9930 8605 10062 8610
rect 11102 8386 11130 8807
rect 11438 8833 11466 9198
rect 11438 8807 11439 8833
rect 11465 8807 11466 8833
rect 11438 8801 11466 8807
rect 11158 8722 11186 8727
rect 11494 8722 11522 9479
rect 11158 8721 11522 8722
rect 11158 8695 11159 8721
rect 11185 8695 11522 8721
rect 11158 8694 11522 8695
rect 11158 8689 11186 8694
rect 11102 8353 11130 8358
rect 9478 7658 9506 7966
rect 9702 7937 9730 7943
rect 9702 7911 9703 7937
rect 9729 7911 9730 7937
rect 9646 7770 9674 7775
rect 9702 7770 9730 7911
rect 9646 7769 9730 7770
rect 9646 7743 9647 7769
rect 9673 7743 9730 7769
rect 9646 7742 9730 7743
rect 9870 7937 9898 7943
rect 9870 7911 9871 7937
rect 9897 7911 9898 7937
rect 9870 7770 9898 7911
rect 10038 7938 10066 7957
rect 10038 7905 10066 7910
rect 10206 7938 10234 7943
rect 10206 7891 10234 7910
rect 9930 7854 10062 7859
rect 9958 7826 9982 7854
rect 10010 7826 10034 7854
rect 9930 7821 10062 7826
rect 9646 7737 9674 7742
rect 9870 7737 9898 7742
rect 9478 7265 9506 7630
rect 9478 7239 9479 7265
rect 9505 7239 9506 7265
rect 9478 7233 9506 7239
rect 9590 7657 9618 7663
rect 9590 7631 9591 7657
rect 9617 7631 9618 7657
rect 9422 2249 9450 2254
rect 9534 2114 9562 2119
rect 9254 1695 9255 1721
rect 9281 1695 9282 1721
rect 9254 1689 9282 1695
rect 9422 2113 9562 2114
rect 9422 2087 9535 2113
rect 9561 2087 9562 2113
rect 9422 2086 9562 2087
rect 9422 1777 9450 2086
rect 9534 2081 9562 2086
rect 9422 1751 9423 1777
rect 9449 1751 9450 1777
rect 8974 1246 9226 1274
rect 8750 400 8778 1246
rect 9086 400 9114 1246
rect 9422 400 9450 1751
rect 9590 1721 9618 7631
rect 9870 7658 9898 7663
rect 9870 7611 9898 7630
rect 10262 7658 10290 7663
rect 10262 7657 10346 7658
rect 10262 7631 10263 7657
rect 10289 7631 10346 7657
rect 10262 7630 10346 7631
rect 10262 7625 10290 7630
rect 10318 7574 10346 7630
rect 10710 7657 10738 7663
rect 10710 7631 10711 7657
rect 10737 7631 10738 7657
rect 10710 7574 10738 7631
rect 10318 7546 10570 7574
rect 9870 7265 9898 7271
rect 9870 7239 9871 7265
rect 9897 7239 9898 7265
rect 9870 2506 9898 7239
rect 10318 7265 10346 7271
rect 10318 7239 10319 7265
rect 10345 7239 10346 7265
rect 9930 7070 10062 7075
rect 9958 7042 9982 7070
rect 10010 7042 10034 7070
rect 9930 7037 10062 7042
rect 9930 6286 10062 6291
rect 9958 6258 9982 6286
rect 10010 6258 10034 6286
rect 9930 6253 10062 6258
rect 10318 5922 10346 7239
rect 10318 5889 10346 5894
rect 9930 5502 10062 5507
rect 9958 5474 9982 5502
rect 10010 5474 10034 5502
rect 9930 5469 10062 5474
rect 9930 4718 10062 4723
rect 9958 4690 9982 4718
rect 10010 4690 10034 4718
rect 9930 4685 10062 4690
rect 9930 3934 10062 3939
rect 9958 3906 9982 3934
rect 10010 3906 10034 3934
rect 9930 3901 10062 3906
rect 9930 3150 10062 3155
rect 9958 3122 9982 3150
rect 10010 3122 10034 3150
rect 9930 3117 10062 3122
rect 9870 2473 9898 2478
rect 9930 2366 10062 2371
rect 9958 2338 9982 2366
rect 10010 2338 10034 2366
rect 9930 2333 10062 2338
rect 9926 2282 9954 2287
rect 9870 2114 9898 2119
rect 9590 1695 9591 1721
rect 9617 1695 9618 1721
rect 9590 1689 9618 1695
rect 9758 2113 9898 2114
rect 9758 2087 9871 2113
rect 9897 2087 9898 2113
rect 9758 2086 9898 2087
rect 9758 1777 9786 2086
rect 9870 2081 9898 2086
rect 9758 1751 9759 1777
rect 9785 1751 9786 1777
rect 9758 400 9786 1751
rect 9926 1721 9954 2254
rect 10150 2114 10178 2119
rect 9926 1695 9927 1721
rect 9953 1695 9954 1721
rect 9926 1689 9954 1695
rect 10094 2113 10178 2114
rect 10094 2087 10151 2113
rect 10177 2087 10178 2113
rect 10094 2086 10178 2087
rect 10094 1777 10122 2086
rect 10150 2081 10178 2086
rect 10430 2113 10458 2119
rect 10430 2087 10431 2113
rect 10457 2087 10458 2113
rect 10094 1751 10095 1777
rect 10121 1751 10122 1777
rect 9930 1582 10062 1587
rect 9958 1554 9982 1582
rect 10010 1554 10034 1582
rect 9930 1549 10062 1554
rect 10094 400 10122 1751
rect 10430 1274 10458 2087
rect 10542 1721 10570 7546
rect 10654 7546 10738 7574
rect 10654 1946 10682 7546
rect 11550 6818 11578 9590
rect 11662 9505 11690 9511
rect 11662 9479 11663 9505
rect 11689 9479 11690 9505
rect 11662 9338 11690 9479
rect 11662 9305 11690 9310
rect 12166 9506 12194 9511
rect 11718 9226 11746 9231
rect 11718 9179 11746 9198
rect 12166 9225 12194 9478
rect 14592 9422 14724 9427
rect 14620 9394 14644 9422
rect 14672 9394 14696 9422
rect 14592 9389 14724 9394
rect 12166 9199 12167 9225
rect 12193 9199 12194 9225
rect 12166 9193 12194 9199
rect 17822 9338 17850 9343
rect 12670 9170 12698 9175
rect 12670 9123 12698 9142
rect 12950 9169 12978 9175
rect 12950 9143 12951 9169
rect 12977 9143 12978 9169
rect 12261 9030 12393 9035
rect 12289 9002 12313 9030
rect 12341 9002 12365 9030
rect 12261 8997 12393 9002
rect 12950 8946 12978 9143
rect 16923 9030 17055 9035
rect 16951 9002 16975 9030
rect 17003 9002 17027 9030
rect 16923 8997 17055 9002
rect 12950 8913 12978 8918
rect 12222 8890 12250 8895
rect 11718 8834 11746 8839
rect 11718 8787 11746 8806
rect 12222 8833 12250 8862
rect 12222 8807 12223 8833
rect 12249 8807 12250 8833
rect 12222 8801 12250 8807
rect 14592 8638 14724 8643
rect 14620 8610 14644 8638
rect 14672 8610 14696 8638
rect 14592 8605 14724 8610
rect 12261 8246 12393 8251
rect 12289 8218 12313 8246
rect 12341 8218 12365 8246
rect 12261 8213 12393 8218
rect 16923 8246 17055 8251
rect 16951 8218 16975 8246
rect 17003 8218 17027 8246
rect 16923 8213 17055 8218
rect 12614 7938 12642 7943
rect 11550 6785 11578 6790
rect 12166 7770 12194 7775
rect 11214 5922 11242 5927
rect 10766 2114 10794 2119
rect 10766 2113 11018 2114
rect 10766 2087 10767 2113
rect 10793 2087 11018 2113
rect 10766 2086 11018 2087
rect 10766 2081 10794 2086
rect 10654 1918 10906 1946
rect 10542 1695 10543 1721
rect 10569 1695 10570 1721
rect 10542 1689 10570 1695
rect 10654 1777 10682 1783
rect 10654 1751 10655 1777
rect 10681 1751 10682 1777
rect 10654 1274 10682 1751
rect 10430 1246 10682 1274
rect 10766 1722 10794 1727
rect 10430 400 10458 1246
rect 10766 400 10794 1694
rect 10878 1721 10906 1918
rect 10878 1695 10879 1721
rect 10905 1695 10906 1721
rect 10878 1689 10906 1695
rect 10990 1777 11018 2086
rect 10990 1751 10991 1777
rect 11017 1751 11018 1777
rect 10990 1722 11018 1751
rect 10990 1689 11018 1694
rect 11102 2113 11130 2119
rect 11102 2087 11103 2113
rect 11129 2087 11130 2113
rect 11102 1274 11130 2087
rect 11214 1721 11242 5894
rect 11382 2506 11410 2511
rect 11214 1695 11215 1721
rect 11241 1695 11242 1721
rect 11214 1689 11242 1695
rect 11326 1777 11354 1783
rect 11326 1751 11327 1777
rect 11353 1751 11354 1777
rect 11326 1274 11354 1751
rect 11382 1694 11410 2478
rect 11438 2114 11466 2119
rect 11438 2113 11690 2114
rect 11438 2087 11439 2113
rect 11465 2087 11690 2113
rect 11438 2086 11690 2087
rect 11438 2081 11466 2086
rect 11662 1777 11690 2086
rect 12110 2058 12138 2063
rect 11662 1751 11663 1777
rect 11689 1751 11690 1777
rect 11382 1666 11578 1694
rect 11550 1665 11578 1666
rect 11550 1639 11551 1665
rect 11577 1639 11578 1665
rect 11550 1633 11578 1639
rect 11662 1274 11690 1751
rect 11102 1246 11354 1274
rect 11438 1246 11690 1274
rect 11774 1834 11802 1839
rect 11102 400 11130 1246
rect 11438 400 11466 1246
rect 11774 400 11802 1806
rect 12110 400 12138 2030
rect 12166 1778 12194 7742
rect 12261 7462 12393 7467
rect 12289 7434 12313 7462
rect 12341 7434 12365 7462
rect 12261 7429 12393 7434
rect 12261 6678 12393 6683
rect 12289 6650 12313 6678
rect 12341 6650 12365 6678
rect 12261 6645 12393 6650
rect 12261 5894 12393 5899
rect 12289 5866 12313 5894
rect 12341 5866 12365 5894
rect 12261 5861 12393 5866
rect 12261 5110 12393 5115
rect 12289 5082 12313 5110
rect 12341 5082 12365 5110
rect 12261 5077 12393 5082
rect 12261 4326 12393 4331
rect 12289 4298 12313 4326
rect 12341 4298 12365 4326
rect 12261 4293 12393 4298
rect 12261 3542 12393 3547
rect 12289 3514 12313 3542
rect 12341 3514 12365 3542
rect 12261 3509 12393 3514
rect 12261 2758 12393 2763
rect 12289 2730 12313 2758
rect 12341 2730 12365 2758
rect 12261 2725 12393 2730
rect 12614 2169 12642 7910
rect 14592 7854 14724 7859
rect 14620 7826 14644 7854
rect 14672 7826 14696 7854
rect 14592 7821 14724 7826
rect 17822 7657 17850 9310
rect 18550 9226 18578 10066
rect 18886 10065 18970 10066
rect 18886 10039 18943 10065
rect 18969 10039 18970 10065
rect 18886 10038 18970 10039
rect 18606 9953 18634 9959
rect 18606 9927 18607 9953
rect 18633 9927 18634 9953
rect 18606 9786 18634 9927
rect 18606 9753 18634 9758
rect 18830 9562 18858 9567
rect 18830 9515 18858 9534
rect 18550 9193 18578 9198
rect 18830 9169 18858 9175
rect 18830 9143 18831 9169
rect 18857 9143 18858 9169
rect 18830 9114 18858 9143
rect 18886 9170 18914 10038
rect 18942 10033 18970 10038
rect 19110 10009 19138 10015
rect 19110 9983 19111 10009
rect 19137 9983 19138 10009
rect 19110 9786 19138 9983
rect 19110 9753 19138 9758
rect 19110 9561 19138 9567
rect 19110 9535 19111 9561
rect 19137 9535 19138 9561
rect 18942 9506 18970 9511
rect 18942 9459 18970 9478
rect 19110 9506 19138 9535
rect 19110 9473 19138 9478
rect 19254 9422 19386 9427
rect 19282 9394 19306 9422
rect 19334 9394 19358 9422
rect 19254 9389 19386 9394
rect 18886 9137 18914 9142
rect 18942 9281 18970 9287
rect 18942 9255 18943 9281
rect 18969 9255 18970 9281
rect 18830 9081 18858 9086
rect 18942 8946 18970 9255
rect 19110 9225 19138 9231
rect 19110 9199 19111 9225
rect 19137 9199 19138 9225
rect 19110 9114 19138 9199
rect 19110 9081 19138 9086
rect 18886 8918 18970 8946
rect 18998 8946 19026 8951
rect 18606 8890 18634 8895
rect 18270 8778 18298 8783
rect 18270 8731 18298 8750
rect 18606 8777 18634 8862
rect 18606 8751 18607 8777
rect 18633 8751 18634 8777
rect 18606 8745 18634 8751
rect 18774 8777 18802 8783
rect 18774 8751 18775 8777
rect 18801 8751 18802 8777
rect 18774 8442 18802 8751
rect 18886 8722 18914 8918
rect 18942 8834 18970 8839
rect 18942 8777 18970 8806
rect 18942 8751 18943 8777
rect 18969 8751 18970 8777
rect 18942 8745 18970 8751
rect 18886 8689 18914 8694
rect 18774 8395 18802 8414
rect 18942 8497 18970 8503
rect 18942 8471 18943 8497
rect 18969 8471 18970 8497
rect 18942 8386 18970 8471
rect 18942 8353 18970 8358
rect 18998 8050 19026 8918
rect 19110 8778 19138 8783
rect 19110 8731 19138 8750
rect 19254 8638 19386 8643
rect 19282 8610 19306 8638
rect 19334 8610 19358 8638
rect 19254 8605 19386 8610
rect 19110 8441 19138 8447
rect 19110 8415 19111 8441
rect 19137 8415 19138 8441
rect 19110 8106 19138 8415
rect 19166 8106 19194 8111
rect 19110 8078 19166 8106
rect 19166 8059 19194 8078
rect 17822 7631 17823 7657
rect 17849 7631 17850 7657
rect 17822 7625 17850 7631
rect 18942 8022 19026 8050
rect 16923 7462 17055 7467
rect 16951 7434 16975 7462
rect 17003 7434 17027 7462
rect 16923 7429 17055 7434
rect 18830 7434 18858 7439
rect 18830 7321 18858 7406
rect 18830 7295 18831 7321
rect 18857 7295 18858 7321
rect 18830 7289 18858 7295
rect 18942 7209 18970 8022
rect 19254 7854 19386 7859
rect 19282 7826 19306 7854
rect 19334 7826 19358 7854
rect 19254 7821 19386 7826
rect 18998 7770 19026 7775
rect 18998 7601 19026 7742
rect 18998 7575 18999 7601
rect 19025 7575 19026 7601
rect 18998 7569 19026 7575
rect 19110 7434 19138 7439
rect 19110 7265 19138 7406
rect 19110 7239 19111 7265
rect 19137 7239 19138 7265
rect 19110 7233 19138 7239
rect 18942 7183 18943 7209
rect 18969 7183 18970 7209
rect 18942 7177 18970 7183
rect 14592 7070 14724 7075
rect 14620 7042 14644 7070
rect 14672 7042 14696 7070
rect 14592 7037 14724 7042
rect 19254 7070 19386 7075
rect 19282 7042 19306 7070
rect 19334 7042 19358 7070
rect 19254 7037 19386 7042
rect 18998 6986 19026 6991
rect 17878 6873 17906 6879
rect 17878 6847 17879 6873
rect 17905 6847 17906 6873
rect 17654 6818 17682 6823
rect 17654 6771 17682 6790
rect 17878 6818 17906 6847
rect 17878 6785 17906 6790
rect 18998 6817 19026 6958
rect 18998 6791 18999 6817
rect 19025 6791 19026 6817
rect 18998 6785 19026 6791
rect 16923 6678 17055 6683
rect 16951 6650 16975 6678
rect 17003 6650 17027 6678
rect 16923 6645 17055 6650
rect 14592 6286 14724 6291
rect 14620 6258 14644 6286
rect 14672 6258 14696 6286
rect 14592 6253 14724 6258
rect 19254 6286 19386 6291
rect 19282 6258 19306 6286
rect 19334 6258 19358 6286
rect 19254 6253 19386 6258
rect 16923 5894 17055 5899
rect 16951 5866 16975 5894
rect 17003 5866 17027 5894
rect 16923 5861 17055 5866
rect 14592 5502 14724 5507
rect 14620 5474 14644 5502
rect 14672 5474 14696 5502
rect 14592 5469 14724 5474
rect 19254 5502 19386 5507
rect 19282 5474 19306 5502
rect 19334 5474 19358 5502
rect 19254 5469 19386 5474
rect 16923 5110 17055 5115
rect 16951 5082 16975 5110
rect 17003 5082 17027 5110
rect 16923 5077 17055 5082
rect 14592 4718 14724 4723
rect 14620 4690 14644 4718
rect 14672 4690 14696 4718
rect 14592 4685 14724 4690
rect 19254 4718 19386 4723
rect 19282 4690 19306 4718
rect 19334 4690 19358 4718
rect 19254 4685 19386 4690
rect 16923 4326 17055 4331
rect 16951 4298 16975 4326
rect 17003 4298 17027 4326
rect 16923 4293 17055 4298
rect 14592 3934 14724 3939
rect 14620 3906 14644 3934
rect 14672 3906 14696 3934
rect 14592 3901 14724 3906
rect 19254 3934 19386 3939
rect 19282 3906 19306 3934
rect 19334 3906 19358 3934
rect 19254 3901 19386 3906
rect 16923 3542 17055 3547
rect 16951 3514 16975 3542
rect 17003 3514 17027 3542
rect 16923 3509 17055 3514
rect 14592 3150 14724 3155
rect 14620 3122 14644 3150
rect 14672 3122 14696 3150
rect 14592 3117 14724 3122
rect 19254 3150 19386 3155
rect 19282 3122 19306 3150
rect 19334 3122 19358 3150
rect 19254 3117 19386 3122
rect 16923 2758 17055 2763
rect 16951 2730 16975 2758
rect 17003 2730 17027 2758
rect 16923 2725 17055 2730
rect 14592 2366 14724 2371
rect 14620 2338 14644 2366
rect 14672 2338 14696 2366
rect 14592 2333 14724 2338
rect 19254 2366 19386 2371
rect 19282 2338 19306 2366
rect 19334 2338 19358 2366
rect 19254 2333 19386 2338
rect 12614 2143 12615 2169
rect 12641 2143 12642 2169
rect 12614 2137 12642 2143
rect 13118 2058 13146 2063
rect 13118 2011 13146 2030
rect 12261 1974 12393 1979
rect 12289 1946 12313 1974
rect 12341 1946 12365 1974
rect 12261 1941 12393 1946
rect 16923 1974 17055 1979
rect 16951 1946 16975 1974
rect 17003 1946 17027 1974
rect 16923 1941 17055 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 12278 1778 12306 1783
rect 12166 1777 12306 1778
rect 12166 1751 12279 1777
rect 12305 1751 12306 1777
rect 12166 1750 12306 1751
rect 12278 1745 12306 1750
rect 14592 1582 14724 1587
rect 14620 1554 14644 1582
rect 14672 1554 14696 1582
rect 14592 1549 14724 1554
rect 19254 1582 19386 1587
rect 19282 1554 19306 1582
rect 19334 1554 19358 1582
rect 19254 1549 19386 1554
rect 6384 0 6440 400
rect 6720 0 6776 400
rect 7056 0 7112 400
rect 7392 0 7448 400
rect 7728 0 7784 400
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 9744 0 9800 400
rect 10080 0 10136 400
rect 10416 0 10472 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 11424 0 11480 400
rect 11760 0 11816 400
rect 12096 0 12152 400
<< via2 >>
rect 2937 18437 2965 18438
rect 2937 18411 2938 18437
rect 2938 18411 2964 18437
rect 2964 18411 2965 18437
rect 2937 18410 2965 18411
rect 2989 18437 3017 18438
rect 2989 18411 2990 18437
rect 2990 18411 3016 18437
rect 3016 18411 3017 18437
rect 2989 18410 3017 18411
rect 3041 18437 3069 18438
rect 3041 18411 3042 18437
rect 3042 18411 3068 18437
rect 3068 18411 3069 18437
rect 3041 18410 3069 18411
rect 7599 18437 7627 18438
rect 7599 18411 7600 18437
rect 7600 18411 7626 18437
rect 7626 18411 7627 18437
rect 7599 18410 7627 18411
rect 7651 18437 7679 18438
rect 7651 18411 7652 18437
rect 7652 18411 7678 18437
rect 7678 18411 7679 18437
rect 7651 18410 7679 18411
rect 7703 18437 7731 18438
rect 7703 18411 7704 18437
rect 7704 18411 7730 18437
rect 7730 18411 7731 18437
rect 7703 18410 7731 18411
rect 5268 18045 5296 18046
rect 5268 18019 5269 18045
rect 5269 18019 5295 18045
rect 5295 18019 5296 18045
rect 5268 18018 5296 18019
rect 5320 18045 5348 18046
rect 5320 18019 5321 18045
rect 5321 18019 5347 18045
rect 5347 18019 5348 18045
rect 5320 18018 5348 18019
rect 5372 18045 5400 18046
rect 5372 18019 5373 18045
rect 5373 18019 5399 18045
rect 5399 18019 5400 18045
rect 5372 18018 5400 18019
rect 7518 17961 7546 17962
rect 7518 17935 7519 17961
rect 7519 17935 7545 17961
rect 7545 17935 7546 17961
rect 7518 17934 7546 17935
rect 8414 18326 8442 18354
rect 7854 17934 7882 17962
rect 2937 17653 2965 17654
rect 2937 17627 2938 17653
rect 2938 17627 2964 17653
rect 2964 17627 2965 17653
rect 2937 17626 2965 17627
rect 2989 17653 3017 17654
rect 2989 17627 2990 17653
rect 2990 17627 3016 17653
rect 3016 17627 3017 17653
rect 2989 17626 3017 17627
rect 3041 17653 3069 17654
rect 3041 17627 3042 17653
rect 3042 17627 3068 17653
rect 3068 17627 3069 17653
rect 3041 17626 3069 17627
rect 7599 17653 7627 17654
rect 7599 17627 7600 17653
rect 7600 17627 7626 17653
rect 7626 17627 7627 17653
rect 7599 17626 7627 17627
rect 7651 17653 7679 17654
rect 7651 17627 7652 17653
rect 7652 17627 7678 17653
rect 7678 17627 7679 17653
rect 7651 17626 7679 17627
rect 7703 17653 7731 17654
rect 7703 17627 7704 17653
rect 7704 17627 7730 17653
rect 7730 17627 7731 17653
rect 7703 17626 7731 17627
rect 5268 17261 5296 17262
rect 5268 17235 5269 17261
rect 5269 17235 5295 17261
rect 5295 17235 5296 17261
rect 5268 17234 5296 17235
rect 5320 17261 5348 17262
rect 5320 17235 5321 17261
rect 5321 17235 5347 17261
rect 5347 17235 5348 17261
rect 5320 17234 5348 17235
rect 5372 17261 5400 17262
rect 5372 17235 5373 17261
rect 5373 17235 5399 17261
rect 5399 17235 5400 17261
rect 5372 17234 5400 17235
rect 2937 16869 2965 16870
rect 2937 16843 2938 16869
rect 2938 16843 2964 16869
rect 2964 16843 2965 16869
rect 2937 16842 2965 16843
rect 2989 16869 3017 16870
rect 2989 16843 2990 16869
rect 2990 16843 3016 16869
rect 3016 16843 3017 16869
rect 2989 16842 3017 16843
rect 3041 16869 3069 16870
rect 3041 16843 3042 16869
rect 3042 16843 3068 16869
rect 3068 16843 3069 16869
rect 3041 16842 3069 16843
rect 7599 16869 7627 16870
rect 7599 16843 7600 16869
rect 7600 16843 7626 16869
rect 7626 16843 7627 16869
rect 7599 16842 7627 16843
rect 7651 16869 7679 16870
rect 7651 16843 7652 16869
rect 7652 16843 7678 16869
rect 7678 16843 7679 16869
rect 7651 16842 7679 16843
rect 7703 16869 7731 16870
rect 7703 16843 7704 16869
rect 7704 16843 7730 16869
rect 7730 16843 7731 16869
rect 7703 16842 7731 16843
rect 5268 16477 5296 16478
rect 5268 16451 5269 16477
rect 5269 16451 5295 16477
rect 5295 16451 5296 16477
rect 5268 16450 5296 16451
rect 5320 16477 5348 16478
rect 5320 16451 5321 16477
rect 5321 16451 5347 16477
rect 5347 16451 5348 16477
rect 5320 16450 5348 16451
rect 5372 16477 5400 16478
rect 5372 16451 5373 16477
rect 5373 16451 5399 16477
rect 5399 16451 5400 16477
rect 5372 16450 5400 16451
rect 2937 16085 2965 16086
rect 2937 16059 2938 16085
rect 2938 16059 2964 16085
rect 2964 16059 2965 16085
rect 2937 16058 2965 16059
rect 2989 16085 3017 16086
rect 2989 16059 2990 16085
rect 2990 16059 3016 16085
rect 3016 16059 3017 16085
rect 2989 16058 3017 16059
rect 3041 16085 3069 16086
rect 3041 16059 3042 16085
rect 3042 16059 3068 16085
rect 3068 16059 3069 16085
rect 3041 16058 3069 16059
rect 7599 16085 7627 16086
rect 7599 16059 7600 16085
rect 7600 16059 7626 16085
rect 7626 16059 7627 16085
rect 7599 16058 7627 16059
rect 7651 16085 7679 16086
rect 7651 16059 7652 16085
rect 7652 16059 7678 16085
rect 7678 16059 7679 16085
rect 7651 16058 7679 16059
rect 7703 16085 7731 16086
rect 7703 16059 7704 16085
rect 7704 16059 7730 16085
rect 7730 16059 7731 16085
rect 7703 16058 7731 16059
rect 5268 15693 5296 15694
rect 5268 15667 5269 15693
rect 5269 15667 5295 15693
rect 5295 15667 5296 15693
rect 5268 15666 5296 15667
rect 5320 15693 5348 15694
rect 5320 15667 5321 15693
rect 5321 15667 5347 15693
rect 5347 15667 5348 15693
rect 5320 15666 5348 15667
rect 5372 15693 5400 15694
rect 5372 15667 5373 15693
rect 5373 15667 5399 15693
rect 5399 15667 5400 15693
rect 5372 15666 5400 15667
rect 2937 15301 2965 15302
rect 2937 15275 2938 15301
rect 2938 15275 2964 15301
rect 2964 15275 2965 15301
rect 2937 15274 2965 15275
rect 2989 15301 3017 15302
rect 2989 15275 2990 15301
rect 2990 15275 3016 15301
rect 3016 15275 3017 15301
rect 2989 15274 3017 15275
rect 3041 15301 3069 15302
rect 3041 15275 3042 15301
rect 3042 15275 3068 15301
rect 3068 15275 3069 15301
rect 3041 15274 3069 15275
rect 7599 15301 7627 15302
rect 7599 15275 7600 15301
rect 7600 15275 7626 15301
rect 7626 15275 7627 15301
rect 7599 15274 7627 15275
rect 7651 15301 7679 15302
rect 7651 15275 7652 15301
rect 7652 15275 7678 15301
rect 7678 15275 7679 15301
rect 7651 15274 7679 15275
rect 7703 15301 7731 15302
rect 7703 15275 7704 15301
rect 7704 15275 7730 15301
rect 7730 15275 7731 15301
rect 7703 15274 7731 15275
rect 8302 15078 8330 15106
rect 8022 14966 8050 14994
rect 8414 14966 8442 14994
rect 5268 14909 5296 14910
rect 5268 14883 5269 14909
rect 5269 14883 5295 14909
rect 5295 14883 5296 14909
rect 5268 14882 5296 14883
rect 5320 14909 5348 14910
rect 5320 14883 5321 14909
rect 5321 14883 5347 14909
rect 5347 14883 5348 14909
rect 5320 14882 5348 14883
rect 5372 14909 5400 14910
rect 5372 14883 5373 14909
rect 5373 14883 5399 14909
rect 5399 14883 5400 14909
rect 5372 14882 5400 14883
rect 2937 14517 2965 14518
rect 2937 14491 2938 14517
rect 2938 14491 2964 14517
rect 2964 14491 2965 14517
rect 2937 14490 2965 14491
rect 2989 14517 3017 14518
rect 2989 14491 2990 14517
rect 2990 14491 3016 14517
rect 3016 14491 3017 14517
rect 2989 14490 3017 14491
rect 3041 14517 3069 14518
rect 3041 14491 3042 14517
rect 3042 14491 3068 14517
rect 3068 14491 3069 14517
rect 3041 14490 3069 14491
rect 7599 14517 7627 14518
rect 7599 14491 7600 14517
rect 7600 14491 7626 14517
rect 7626 14491 7627 14517
rect 7599 14490 7627 14491
rect 7651 14517 7679 14518
rect 7651 14491 7652 14517
rect 7652 14491 7678 14517
rect 7678 14491 7679 14517
rect 7651 14490 7679 14491
rect 7703 14517 7731 14518
rect 7703 14491 7704 14517
rect 7704 14491 7730 14517
rect 7730 14491 7731 14517
rect 7703 14490 7731 14491
rect 5268 14125 5296 14126
rect 5268 14099 5269 14125
rect 5269 14099 5295 14125
rect 5295 14099 5296 14125
rect 5268 14098 5296 14099
rect 5320 14125 5348 14126
rect 5320 14099 5321 14125
rect 5321 14099 5347 14125
rect 5347 14099 5348 14125
rect 5320 14098 5348 14099
rect 5372 14125 5400 14126
rect 5372 14099 5373 14125
rect 5373 14099 5399 14125
rect 5399 14099 5400 14125
rect 5372 14098 5400 14099
rect 2937 13733 2965 13734
rect 2937 13707 2938 13733
rect 2938 13707 2964 13733
rect 2964 13707 2965 13733
rect 2937 13706 2965 13707
rect 2989 13733 3017 13734
rect 2989 13707 2990 13733
rect 2990 13707 3016 13733
rect 3016 13707 3017 13733
rect 2989 13706 3017 13707
rect 3041 13733 3069 13734
rect 3041 13707 3042 13733
rect 3042 13707 3068 13733
rect 3068 13707 3069 13733
rect 3041 13706 3069 13707
rect 7599 13733 7627 13734
rect 7599 13707 7600 13733
rect 7600 13707 7626 13733
rect 7626 13707 7627 13733
rect 7599 13706 7627 13707
rect 7651 13733 7679 13734
rect 7651 13707 7652 13733
rect 7652 13707 7678 13733
rect 7678 13707 7679 13733
rect 7651 13706 7679 13707
rect 7703 13733 7731 13734
rect 7703 13707 7704 13733
rect 7704 13707 7730 13733
rect 7730 13707 7731 13733
rect 7703 13706 7731 13707
rect 5268 13341 5296 13342
rect 5268 13315 5269 13341
rect 5269 13315 5295 13341
rect 5295 13315 5296 13341
rect 5268 13314 5296 13315
rect 5320 13341 5348 13342
rect 5320 13315 5321 13341
rect 5321 13315 5347 13341
rect 5347 13315 5348 13341
rect 5320 13314 5348 13315
rect 5372 13341 5400 13342
rect 5372 13315 5373 13341
rect 5373 13315 5399 13341
rect 5399 13315 5400 13341
rect 5372 13314 5400 13315
rect 966 12782 994 12810
rect 854 12446 882 12474
rect 1022 12417 1050 12418
rect 1022 12391 1023 12417
rect 1023 12391 1049 12417
rect 1049 12391 1050 12417
rect 1022 12390 1050 12391
rect 854 12110 882 12138
rect 1022 11857 1050 11858
rect 1022 11831 1023 11857
rect 1023 11831 1049 11857
rect 1049 11831 1050 11857
rect 1022 11830 1050 11831
rect 854 11774 882 11802
rect 854 11438 882 11466
rect 1022 11158 1050 11186
rect 854 11129 882 11130
rect 854 11103 855 11129
rect 855 11103 881 11129
rect 881 11103 882 11129
rect 854 11102 882 11103
rect 1022 10849 1050 10850
rect 1022 10823 1023 10849
rect 1023 10823 1049 10849
rect 1049 10823 1050 10849
rect 1022 10822 1050 10823
rect 854 10710 882 10738
rect 854 10430 882 10458
rect 1078 10318 1106 10346
rect 1022 10289 1050 10290
rect 1022 10263 1023 10289
rect 1023 10263 1049 10289
rect 1049 10263 1050 10289
rect 1022 10262 1050 10263
rect 854 10094 882 10122
rect 966 9897 994 9898
rect 966 9871 967 9897
rect 967 9871 993 9897
rect 993 9871 994 9897
rect 966 9870 994 9871
rect 1246 12446 1274 12474
rect 1246 12110 1274 12138
rect 1246 11774 1274 11802
rect 1246 11438 1274 11466
rect 1246 11102 1274 11130
rect 1358 11073 1386 11074
rect 1358 11047 1359 11073
rect 1359 11047 1385 11073
rect 1385 11047 1386 11073
rect 1358 11046 1386 11047
rect 1190 10766 1218 10794
rect 1582 10766 1610 10794
rect 1470 10737 1498 10738
rect 1470 10711 1471 10737
rect 1471 10711 1497 10737
rect 1497 10711 1498 10737
rect 1470 10710 1498 10711
rect 1246 10094 1274 10122
rect 2937 12949 2965 12950
rect 2937 12923 2938 12949
rect 2938 12923 2964 12949
rect 2964 12923 2965 12949
rect 2937 12922 2965 12923
rect 2989 12949 3017 12950
rect 2989 12923 2990 12949
rect 2990 12923 3016 12949
rect 3016 12923 3017 12949
rect 2989 12922 3017 12923
rect 3041 12949 3069 12950
rect 3041 12923 3042 12949
rect 3042 12923 3068 12949
rect 3068 12923 3069 12949
rect 3041 12922 3069 12923
rect 7599 12949 7627 12950
rect 7599 12923 7600 12949
rect 7600 12923 7626 12949
rect 7626 12923 7627 12949
rect 7599 12922 7627 12923
rect 7651 12949 7679 12950
rect 7651 12923 7652 12949
rect 7652 12923 7678 12949
rect 7678 12923 7679 12949
rect 7651 12922 7679 12923
rect 7703 12949 7731 12950
rect 7703 12923 7704 12949
rect 7704 12923 7730 12949
rect 7730 12923 7731 12949
rect 7703 12922 7731 12923
rect 5268 12557 5296 12558
rect 5268 12531 5269 12557
rect 5269 12531 5295 12557
rect 5295 12531 5296 12557
rect 5268 12530 5296 12531
rect 5320 12557 5348 12558
rect 5320 12531 5321 12557
rect 5321 12531 5347 12557
rect 5347 12531 5348 12557
rect 5320 12530 5348 12531
rect 5372 12557 5400 12558
rect 5372 12531 5373 12557
rect 5373 12531 5399 12557
rect 5399 12531 5400 12557
rect 5372 12530 5400 12531
rect 8022 12390 8050 12418
rect 2937 12165 2965 12166
rect 2937 12139 2938 12165
rect 2938 12139 2964 12165
rect 2964 12139 2965 12165
rect 2937 12138 2965 12139
rect 2989 12165 3017 12166
rect 2989 12139 2990 12165
rect 2990 12139 3016 12165
rect 3016 12139 3017 12165
rect 2989 12138 3017 12139
rect 3041 12165 3069 12166
rect 3041 12139 3042 12165
rect 3042 12139 3068 12165
rect 3068 12139 3069 12165
rect 3041 12138 3069 12139
rect 7599 12165 7627 12166
rect 7599 12139 7600 12165
rect 7600 12139 7626 12165
rect 7626 12139 7627 12165
rect 7599 12138 7627 12139
rect 7651 12165 7679 12166
rect 7651 12139 7652 12165
rect 7652 12139 7678 12165
rect 7678 12139 7679 12165
rect 7651 12138 7679 12139
rect 7703 12165 7731 12166
rect 7703 12139 7704 12165
rect 7704 12139 7730 12165
rect 7730 12139 7731 12165
rect 7703 12138 7731 12139
rect 8022 11830 8050 11858
rect 5268 11773 5296 11774
rect 5268 11747 5269 11773
rect 5269 11747 5295 11773
rect 5295 11747 5296 11773
rect 5268 11746 5296 11747
rect 5320 11773 5348 11774
rect 5320 11747 5321 11773
rect 5321 11747 5347 11773
rect 5347 11747 5348 11773
rect 5320 11746 5348 11747
rect 5372 11773 5400 11774
rect 5372 11747 5373 11773
rect 5373 11747 5399 11773
rect 5399 11747 5400 11773
rect 5372 11746 5400 11747
rect 2937 11381 2965 11382
rect 2937 11355 2938 11381
rect 2938 11355 2964 11381
rect 2964 11355 2965 11381
rect 2937 11354 2965 11355
rect 2989 11381 3017 11382
rect 2989 11355 2990 11381
rect 2990 11355 3016 11381
rect 3016 11355 3017 11381
rect 2989 11354 3017 11355
rect 3041 11381 3069 11382
rect 3041 11355 3042 11381
rect 3042 11355 3068 11381
rect 3068 11355 3069 11381
rect 3041 11354 3069 11355
rect 7599 11381 7627 11382
rect 7599 11355 7600 11381
rect 7600 11355 7626 11381
rect 7626 11355 7627 11381
rect 7599 11354 7627 11355
rect 7651 11381 7679 11382
rect 7651 11355 7652 11381
rect 7652 11355 7678 11381
rect 7678 11355 7679 11381
rect 7651 11354 7679 11355
rect 7703 11381 7731 11382
rect 7703 11355 7704 11381
rect 7704 11355 7730 11381
rect 7730 11355 7731 11381
rect 7703 11354 7731 11355
rect 7854 11158 7882 11186
rect 5268 10989 5296 10990
rect 5268 10963 5269 10989
rect 5269 10963 5295 10989
rect 5295 10963 5296 10989
rect 5268 10962 5296 10963
rect 5320 10989 5348 10990
rect 5320 10963 5321 10989
rect 5321 10963 5347 10989
rect 5347 10963 5348 10989
rect 5320 10962 5348 10963
rect 5372 10989 5400 10990
rect 5372 10963 5373 10989
rect 5373 10963 5399 10989
rect 5399 10963 5400 10989
rect 5372 10962 5400 10963
rect 2937 10597 2965 10598
rect 2937 10571 2938 10597
rect 2938 10571 2964 10597
rect 2964 10571 2965 10597
rect 2937 10570 2965 10571
rect 2989 10597 3017 10598
rect 2989 10571 2990 10597
rect 2990 10571 3016 10597
rect 3016 10571 3017 10597
rect 2989 10570 3017 10571
rect 3041 10597 3069 10598
rect 3041 10571 3042 10597
rect 3042 10571 3068 10597
rect 3068 10571 3069 10597
rect 3041 10570 3069 10571
rect 7599 10597 7627 10598
rect 7599 10571 7600 10597
rect 7600 10571 7626 10597
rect 7626 10571 7627 10597
rect 7599 10570 7627 10571
rect 7651 10597 7679 10598
rect 7651 10571 7652 10597
rect 7652 10571 7678 10597
rect 7678 10571 7679 10597
rect 7651 10570 7679 10571
rect 7703 10597 7731 10598
rect 7703 10571 7704 10597
rect 7704 10571 7730 10597
rect 7730 10571 7731 10597
rect 7703 10570 7731 10571
rect 9030 18353 9058 18354
rect 9030 18327 9031 18353
rect 9031 18327 9057 18353
rect 9057 18327 9058 18353
rect 9030 18326 9058 18327
rect 8694 15078 8722 15106
rect 8526 11857 8554 11858
rect 8526 11831 8527 11857
rect 8527 11831 8553 11857
rect 8553 11831 8554 11857
rect 8526 11830 8554 11831
rect 8806 11830 8834 11858
rect 9478 17934 9506 17962
rect 9930 18045 9958 18046
rect 9930 18019 9931 18045
rect 9931 18019 9957 18045
rect 9957 18019 9958 18045
rect 9930 18018 9958 18019
rect 9982 18045 10010 18046
rect 9982 18019 9983 18045
rect 9983 18019 10009 18045
rect 10009 18019 10010 18045
rect 9982 18018 10010 18019
rect 10034 18045 10062 18046
rect 10034 18019 10035 18045
rect 10035 18019 10061 18045
rect 10061 18019 10062 18045
rect 10034 18018 10062 18019
rect 9870 17961 9898 17962
rect 9870 17935 9871 17961
rect 9871 17935 9897 17961
rect 9897 17935 9898 17961
rect 9870 17934 9898 17935
rect 9930 17261 9958 17262
rect 9930 17235 9931 17261
rect 9931 17235 9957 17261
rect 9957 17235 9958 17261
rect 9930 17234 9958 17235
rect 9982 17261 10010 17262
rect 9982 17235 9983 17261
rect 9983 17235 10009 17261
rect 10009 17235 10010 17261
rect 9982 17234 10010 17235
rect 10034 17261 10062 17262
rect 10034 17235 10035 17261
rect 10035 17235 10061 17261
rect 10061 17235 10062 17261
rect 10034 17234 10062 17235
rect 9930 16477 9958 16478
rect 9930 16451 9931 16477
rect 9931 16451 9957 16477
rect 9957 16451 9958 16477
rect 9930 16450 9958 16451
rect 9982 16477 10010 16478
rect 9982 16451 9983 16477
rect 9983 16451 10009 16477
rect 10009 16451 10010 16477
rect 9982 16450 10010 16451
rect 10034 16477 10062 16478
rect 10034 16451 10035 16477
rect 10035 16451 10061 16477
rect 10061 16451 10062 16477
rect 10034 16450 10062 16451
rect 9930 15693 9958 15694
rect 9930 15667 9931 15693
rect 9931 15667 9957 15693
rect 9957 15667 9958 15693
rect 9930 15666 9958 15667
rect 9982 15693 10010 15694
rect 9982 15667 9983 15693
rect 9983 15667 10009 15693
rect 10009 15667 10010 15693
rect 9982 15666 10010 15667
rect 10034 15693 10062 15694
rect 10034 15667 10035 15693
rect 10035 15667 10061 15693
rect 10061 15667 10062 15693
rect 10034 15666 10062 15667
rect 9930 14909 9958 14910
rect 9930 14883 9931 14909
rect 9931 14883 9957 14909
rect 9957 14883 9958 14909
rect 9930 14882 9958 14883
rect 9982 14909 10010 14910
rect 9982 14883 9983 14909
rect 9983 14883 10009 14909
rect 10009 14883 10010 14909
rect 9982 14882 10010 14883
rect 10034 14909 10062 14910
rect 10034 14883 10035 14909
rect 10035 14883 10061 14909
rect 10061 14883 10062 14909
rect 10034 14882 10062 14883
rect 12261 18437 12289 18438
rect 12261 18411 12262 18437
rect 12262 18411 12288 18437
rect 12288 18411 12289 18437
rect 12261 18410 12289 18411
rect 12313 18437 12341 18438
rect 12313 18411 12314 18437
rect 12314 18411 12340 18437
rect 12340 18411 12341 18437
rect 12313 18410 12341 18411
rect 12365 18437 12393 18438
rect 12365 18411 12366 18437
rect 12366 18411 12392 18437
rect 12392 18411 12393 18437
rect 12365 18410 12393 18411
rect 16923 18437 16951 18438
rect 16923 18411 16924 18437
rect 16924 18411 16950 18437
rect 16950 18411 16951 18437
rect 16923 18410 16951 18411
rect 16975 18437 17003 18438
rect 16975 18411 16976 18437
rect 16976 18411 17002 18437
rect 17002 18411 17003 18437
rect 16975 18410 17003 18411
rect 17027 18437 17055 18438
rect 17027 18411 17028 18437
rect 17028 18411 17054 18437
rect 17054 18411 17055 18437
rect 17027 18410 17055 18411
rect 10374 14686 10402 14714
rect 9930 14125 9958 14126
rect 9930 14099 9931 14125
rect 9931 14099 9957 14125
rect 9957 14099 9958 14125
rect 9930 14098 9958 14099
rect 9982 14125 10010 14126
rect 9982 14099 9983 14125
rect 9983 14099 10009 14125
rect 10009 14099 10010 14125
rect 9982 14098 10010 14099
rect 10034 14125 10062 14126
rect 10034 14099 10035 14125
rect 10035 14099 10061 14125
rect 10061 14099 10062 14125
rect 10034 14098 10062 14099
rect 7742 10345 7770 10346
rect 7742 10319 7743 10345
rect 7743 10319 7769 10345
rect 7769 10319 7770 10345
rect 7742 10318 7770 10319
rect 5268 10205 5296 10206
rect 5268 10179 5269 10205
rect 5269 10179 5295 10205
rect 5295 10179 5296 10205
rect 5268 10178 5296 10179
rect 5320 10205 5348 10206
rect 5320 10179 5321 10205
rect 5321 10179 5347 10205
rect 5347 10179 5348 10205
rect 5320 10178 5348 10179
rect 5372 10205 5400 10206
rect 5372 10179 5373 10205
rect 5373 10179 5399 10205
rect 5399 10179 5400 10205
rect 5372 10178 5400 10179
rect 8246 10822 8274 10850
rect 9930 13341 9958 13342
rect 9930 13315 9931 13341
rect 9931 13315 9957 13341
rect 9957 13315 9958 13341
rect 9930 13314 9958 13315
rect 9982 13341 10010 13342
rect 9982 13315 9983 13341
rect 9983 13315 10009 13341
rect 10009 13315 10010 13341
rect 9982 13314 10010 13315
rect 10034 13341 10062 13342
rect 10034 13315 10035 13341
rect 10035 13315 10061 13341
rect 10061 13315 10062 13341
rect 10034 13314 10062 13315
rect 9930 12557 9958 12558
rect 9930 12531 9931 12557
rect 9931 12531 9957 12557
rect 9957 12531 9958 12557
rect 9930 12530 9958 12531
rect 9982 12557 10010 12558
rect 9982 12531 9983 12557
rect 9983 12531 10009 12557
rect 10009 12531 10010 12557
rect 9982 12530 10010 12531
rect 10034 12557 10062 12558
rect 10034 12531 10035 12557
rect 10035 12531 10061 12557
rect 10061 12531 10062 12557
rect 10034 12530 10062 12531
rect 9930 11773 9958 11774
rect 9930 11747 9931 11773
rect 9931 11747 9957 11773
rect 9957 11747 9958 11773
rect 9930 11746 9958 11747
rect 9982 11773 10010 11774
rect 9982 11747 9983 11773
rect 9983 11747 10009 11773
rect 10009 11747 10010 11773
rect 9982 11746 10010 11747
rect 10034 11773 10062 11774
rect 10034 11747 10035 11773
rect 10035 11747 10061 11773
rect 10061 11747 10062 11773
rect 10034 11746 10062 11747
rect 10598 14686 10626 14714
rect 2422 10038 2450 10066
rect 2142 10009 2170 10010
rect 2142 9983 2143 10009
rect 2143 9983 2169 10009
rect 2169 9983 2170 10009
rect 2142 9982 2170 9983
rect 2937 9813 2965 9814
rect 2937 9787 2938 9813
rect 2938 9787 2964 9813
rect 2964 9787 2965 9813
rect 2937 9786 2965 9787
rect 2989 9813 3017 9814
rect 2989 9787 2990 9813
rect 2990 9787 3016 9813
rect 3016 9787 3017 9813
rect 2989 9786 3017 9787
rect 3041 9813 3069 9814
rect 3041 9787 3042 9813
rect 3042 9787 3068 9813
rect 3068 9787 3069 9813
rect 3041 9786 3069 9787
rect 7599 9813 7627 9814
rect 7599 9787 7600 9813
rect 7600 9787 7626 9813
rect 7626 9787 7627 9813
rect 7599 9786 7627 9787
rect 7651 9813 7679 9814
rect 7651 9787 7652 9813
rect 7652 9787 7678 9813
rect 7678 9787 7679 9813
rect 7651 9786 7679 9787
rect 7703 9813 7731 9814
rect 7703 9787 7704 9813
rect 7704 9787 7730 9813
rect 7730 9787 7731 9813
rect 7703 9786 7731 9787
rect 8246 10065 8274 10066
rect 8246 10039 8247 10065
rect 8247 10039 8273 10065
rect 8273 10039 8274 10065
rect 8246 10038 8274 10039
rect 8862 11046 8890 11074
rect 9930 10989 9958 10990
rect 9930 10963 9931 10989
rect 9931 10963 9957 10989
rect 9957 10963 9958 10989
rect 9930 10962 9958 10963
rect 9982 10989 10010 10990
rect 9982 10963 9983 10989
rect 9983 10963 10009 10989
rect 10009 10963 10010 10989
rect 9982 10962 10010 10963
rect 10034 10989 10062 10990
rect 10034 10963 10035 10989
rect 10035 10963 10061 10989
rect 10061 10963 10062 10989
rect 10034 10962 10062 10963
rect 14592 18045 14620 18046
rect 14592 18019 14593 18045
rect 14593 18019 14619 18045
rect 14619 18019 14620 18045
rect 14592 18018 14620 18019
rect 14644 18045 14672 18046
rect 14644 18019 14645 18045
rect 14645 18019 14671 18045
rect 14671 18019 14672 18045
rect 14644 18018 14672 18019
rect 14696 18045 14724 18046
rect 14696 18019 14697 18045
rect 14697 18019 14723 18045
rect 14723 18019 14724 18045
rect 14696 18018 14724 18019
rect 19254 18045 19282 18046
rect 19254 18019 19255 18045
rect 19255 18019 19281 18045
rect 19281 18019 19282 18045
rect 19254 18018 19282 18019
rect 19306 18045 19334 18046
rect 19306 18019 19307 18045
rect 19307 18019 19333 18045
rect 19333 18019 19334 18045
rect 19306 18018 19334 18019
rect 19358 18045 19386 18046
rect 19358 18019 19359 18045
rect 19359 18019 19385 18045
rect 19385 18019 19386 18045
rect 19358 18018 19386 18019
rect 12261 17653 12289 17654
rect 12261 17627 12262 17653
rect 12262 17627 12288 17653
rect 12288 17627 12289 17653
rect 12261 17626 12289 17627
rect 12313 17653 12341 17654
rect 12313 17627 12314 17653
rect 12314 17627 12340 17653
rect 12340 17627 12341 17653
rect 12313 17626 12341 17627
rect 12365 17653 12393 17654
rect 12365 17627 12366 17653
rect 12366 17627 12392 17653
rect 12392 17627 12393 17653
rect 12365 17626 12393 17627
rect 16923 17653 16951 17654
rect 16923 17627 16924 17653
rect 16924 17627 16950 17653
rect 16950 17627 16951 17653
rect 16923 17626 16951 17627
rect 16975 17653 17003 17654
rect 16975 17627 16976 17653
rect 16976 17627 17002 17653
rect 17002 17627 17003 17653
rect 16975 17626 17003 17627
rect 17027 17653 17055 17654
rect 17027 17627 17028 17653
rect 17028 17627 17054 17653
rect 17054 17627 17055 17653
rect 17027 17626 17055 17627
rect 14592 17261 14620 17262
rect 14592 17235 14593 17261
rect 14593 17235 14619 17261
rect 14619 17235 14620 17261
rect 14592 17234 14620 17235
rect 14644 17261 14672 17262
rect 14644 17235 14645 17261
rect 14645 17235 14671 17261
rect 14671 17235 14672 17261
rect 14644 17234 14672 17235
rect 14696 17261 14724 17262
rect 14696 17235 14697 17261
rect 14697 17235 14723 17261
rect 14723 17235 14724 17261
rect 14696 17234 14724 17235
rect 19254 17261 19282 17262
rect 19254 17235 19255 17261
rect 19255 17235 19281 17261
rect 19281 17235 19282 17261
rect 19254 17234 19282 17235
rect 19306 17261 19334 17262
rect 19306 17235 19307 17261
rect 19307 17235 19333 17261
rect 19333 17235 19334 17261
rect 19306 17234 19334 17235
rect 19358 17261 19386 17262
rect 19358 17235 19359 17261
rect 19359 17235 19385 17261
rect 19385 17235 19386 17261
rect 19358 17234 19386 17235
rect 12261 16869 12289 16870
rect 12261 16843 12262 16869
rect 12262 16843 12288 16869
rect 12288 16843 12289 16869
rect 12261 16842 12289 16843
rect 12313 16869 12341 16870
rect 12313 16843 12314 16869
rect 12314 16843 12340 16869
rect 12340 16843 12341 16869
rect 12313 16842 12341 16843
rect 12365 16869 12393 16870
rect 12365 16843 12366 16869
rect 12366 16843 12392 16869
rect 12392 16843 12393 16869
rect 12365 16842 12393 16843
rect 16923 16869 16951 16870
rect 16923 16843 16924 16869
rect 16924 16843 16950 16869
rect 16950 16843 16951 16869
rect 16923 16842 16951 16843
rect 16975 16869 17003 16870
rect 16975 16843 16976 16869
rect 16976 16843 17002 16869
rect 17002 16843 17003 16869
rect 16975 16842 17003 16843
rect 17027 16869 17055 16870
rect 17027 16843 17028 16869
rect 17028 16843 17054 16869
rect 17054 16843 17055 16869
rect 17027 16842 17055 16843
rect 14592 16477 14620 16478
rect 14592 16451 14593 16477
rect 14593 16451 14619 16477
rect 14619 16451 14620 16477
rect 14592 16450 14620 16451
rect 14644 16477 14672 16478
rect 14644 16451 14645 16477
rect 14645 16451 14671 16477
rect 14671 16451 14672 16477
rect 14644 16450 14672 16451
rect 14696 16477 14724 16478
rect 14696 16451 14697 16477
rect 14697 16451 14723 16477
rect 14723 16451 14724 16477
rect 14696 16450 14724 16451
rect 19254 16477 19282 16478
rect 19254 16451 19255 16477
rect 19255 16451 19281 16477
rect 19281 16451 19282 16477
rect 19254 16450 19282 16451
rect 19306 16477 19334 16478
rect 19306 16451 19307 16477
rect 19307 16451 19333 16477
rect 19333 16451 19334 16477
rect 19306 16450 19334 16451
rect 19358 16477 19386 16478
rect 19358 16451 19359 16477
rect 19359 16451 19385 16477
rect 19385 16451 19386 16477
rect 19358 16450 19386 16451
rect 12261 16085 12289 16086
rect 12261 16059 12262 16085
rect 12262 16059 12288 16085
rect 12288 16059 12289 16085
rect 12261 16058 12289 16059
rect 12313 16085 12341 16086
rect 12313 16059 12314 16085
rect 12314 16059 12340 16085
rect 12340 16059 12341 16085
rect 12313 16058 12341 16059
rect 12365 16085 12393 16086
rect 12365 16059 12366 16085
rect 12366 16059 12392 16085
rect 12392 16059 12393 16085
rect 12365 16058 12393 16059
rect 16923 16085 16951 16086
rect 16923 16059 16924 16085
rect 16924 16059 16950 16085
rect 16950 16059 16951 16085
rect 16923 16058 16951 16059
rect 16975 16085 17003 16086
rect 16975 16059 16976 16085
rect 16976 16059 17002 16085
rect 17002 16059 17003 16085
rect 16975 16058 17003 16059
rect 17027 16085 17055 16086
rect 17027 16059 17028 16085
rect 17028 16059 17054 16085
rect 17054 16059 17055 16085
rect 17027 16058 17055 16059
rect 14592 15693 14620 15694
rect 14592 15667 14593 15693
rect 14593 15667 14619 15693
rect 14619 15667 14620 15693
rect 14592 15666 14620 15667
rect 14644 15693 14672 15694
rect 14644 15667 14645 15693
rect 14645 15667 14671 15693
rect 14671 15667 14672 15693
rect 14644 15666 14672 15667
rect 14696 15693 14724 15694
rect 14696 15667 14697 15693
rect 14697 15667 14723 15693
rect 14723 15667 14724 15693
rect 14696 15666 14724 15667
rect 19254 15693 19282 15694
rect 19254 15667 19255 15693
rect 19255 15667 19281 15693
rect 19281 15667 19282 15693
rect 19254 15666 19282 15667
rect 19306 15693 19334 15694
rect 19306 15667 19307 15693
rect 19307 15667 19333 15693
rect 19333 15667 19334 15693
rect 19306 15666 19334 15667
rect 19358 15693 19386 15694
rect 19358 15667 19359 15693
rect 19359 15667 19385 15693
rect 19385 15667 19386 15693
rect 19358 15666 19386 15667
rect 12261 15301 12289 15302
rect 12261 15275 12262 15301
rect 12262 15275 12288 15301
rect 12288 15275 12289 15301
rect 12261 15274 12289 15275
rect 12313 15301 12341 15302
rect 12313 15275 12314 15301
rect 12314 15275 12340 15301
rect 12340 15275 12341 15301
rect 12313 15274 12341 15275
rect 12365 15301 12393 15302
rect 12365 15275 12366 15301
rect 12366 15275 12392 15301
rect 12392 15275 12393 15301
rect 12365 15274 12393 15275
rect 16923 15301 16951 15302
rect 16923 15275 16924 15301
rect 16924 15275 16950 15301
rect 16950 15275 16951 15301
rect 16923 15274 16951 15275
rect 16975 15301 17003 15302
rect 16975 15275 16976 15301
rect 16976 15275 17002 15301
rect 17002 15275 17003 15301
rect 16975 15274 17003 15275
rect 17027 15301 17055 15302
rect 17027 15275 17028 15301
rect 17028 15275 17054 15301
rect 17054 15275 17055 15301
rect 17027 15274 17055 15275
rect 14592 14909 14620 14910
rect 14592 14883 14593 14909
rect 14593 14883 14619 14909
rect 14619 14883 14620 14909
rect 14592 14882 14620 14883
rect 14644 14909 14672 14910
rect 14644 14883 14645 14909
rect 14645 14883 14671 14909
rect 14671 14883 14672 14909
rect 14644 14882 14672 14883
rect 14696 14909 14724 14910
rect 14696 14883 14697 14909
rect 14697 14883 14723 14909
rect 14723 14883 14724 14909
rect 14696 14882 14724 14883
rect 19254 14909 19282 14910
rect 19254 14883 19255 14909
rect 19255 14883 19281 14909
rect 19281 14883 19282 14909
rect 19254 14882 19282 14883
rect 19306 14909 19334 14910
rect 19306 14883 19307 14909
rect 19307 14883 19333 14909
rect 19333 14883 19334 14909
rect 19306 14882 19334 14883
rect 19358 14909 19386 14910
rect 19358 14883 19359 14909
rect 19359 14883 19385 14909
rect 19385 14883 19386 14909
rect 19358 14882 19386 14883
rect 12261 14517 12289 14518
rect 12261 14491 12262 14517
rect 12262 14491 12288 14517
rect 12288 14491 12289 14517
rect 12261 14490 12289 14491
rect 12313 14517 12341 14518
rect 12313 14491 12314 14517
rect 12314 14491 12340 14517
rect 12340 14491 12341 14517
rect 12313 14490 12341 14491
rect 12365 14517 12393 14518
rect 12365 14491 12366 14517
rect 12366 14491 12392 14517
rect 12392 14491 12393 14517
rect 12365 14490 12393 14491
rect 16923 14517 16951 14518
rect 16923 14491 16924 14517
rect 16924 14491 16950 14517
rect 16950 14491 16951 14517
rect 16923 14490 16951 14491
rect 16975 14517 17003 14518
rect 16975 14491 16976 14517
rect 16976 14491 17002 14517
rect 17002 14491 17003 14517
rect 16975 14490 17003 14491
rect 17027 14517 17055 14518
rect 17027 14491 17028 14517
rect 17028 14491 17054 14517
rect 17054 14491 17055 14517
rect 17027 14490 17055 14491
rect 14592 14125 14620 14126
rect 14592 14099 14593 14125
rect 14593 14099 14619 14125
rect 14619 14099 14620 14125
rect 14592 14098 14620 14099
rect 14644 14125 14672 14126
rect 14644 14099 14645 14125
rect 14645 14099 14671 14125
rect 14671 14099 14672 14125
rect 14644 14098 14672 14099
rect 14696 14125 14724 14126
rect 14696 14099 14697 14125
rect 14697 14099 14723 14125
rect 14723 14099 14724 14125
rect 14696 14098 14724 14099
rect 19254 14125 19282 14126
rect 19254 14099 19255 14125
rect 19255 14099 19281 14125
rect 19281 14099 19282 14125
rect 19254 14098 19282 14099
rect 19306 14125 19334 14126
rect 19306 14099 19307 14125
rect 19307 14099 19333 14125
rect 19333 14099 19334 14125
rect 19306 14098 19334 14099
rect 19358 14125 19386 14126
rect 19358 14099 19359 14125
rect 19359 14099 19385 14125
rect 19385 14099 19386 14125
rect 19358 14098 19386 14099
rect 12261 13733 12289 13734
rect 12261 13707 12262 13733
rect 12262 13707 12288 13733
rect 12288 13707 12289 13733
rect 12261 13706 12289 13707
rect 12313 13733 12341 13734
rect 12313 13707 12314 13733
rect 12314 13707 12340 13733
rect 12340 13707 12341 13733
rect 12313 13706 12341 13707
rect 12365 13733 12393 13734
rect 12365 13707 12366 13733
rect 12366 13707 12392 13733
rect 12392 13707 12393 13733
rect 12365 13706 12393 13707
rect 16923 13733 16951 13734
rect 16923 13707 16924 13733
rect 16924 13707 16950 13733
rect 16950 13707 16951 13733
rect 16923 13706 16951 13707
rect 16975 13733 17003 13734
rect 16975 13707 16976 13733
rect 16976 13707 17002 13733
rect 17002 13707 17003 13733
rect 16975 13706 17003 13707
rect 17027 13733 17055 13734
rect 17027 13707 17028 13733
rect 17028 13707 17054 13733
rect 17054 13707 17055 13733
rect 17027 13706 17055 13707
rect 10878 11073 10906 11074
rect 10878 11047 10879 11073
rect 10879 11047 10905 11073
rect 10905 11047 10906 11073
rect 10878 11046 10906 11047
rect 10710 10878 10738 10906
rect 9422 10318 9450 10346
rect 10934 10793 10962 10794
rect 10934 10767 10935 10793
rect 10935 10767 10961 10793
rect 10961 10767 10962 10793
rect 10934 10766 10962 10767
rect 8862 10262 8890 10290
rect 9930 10205 9958 10206
rect 9930 10179 9931 10205
rect 9931 10179 9957 10205
rect 9957 10179 9958 10205
rect 9930 10178 9958 10179
rect 9982 10205 10010 10206
rect 9982 10179 9983 10205
rect 9983 10179 10009 10205
rect 10009 10179 10010 10205
rect 9982 10178 10010 10179
rect 10034 10205 10062 10206
rect 10034 10179 10035 10205
rect 10035 10179 10061 10205
rect 10061 10179 10062 10205
rect 10034 10178 10062 10179
rect 8694 10065 8722 10066
rect 8694 10039 8695 10065
rect 8695 10039 8721 10065
rect 8721 10039 8722 10065
rect 8694 10038 8722 10039
rect 1134 9534 1162 9562
rect 7742 9561 7770 9562
rect 7742 9535 7743 9561
rect 7743 9535 7769 9561
rect 7769 9535 7770 9561
rect 7742 9534 7770 9535
rect 1022 9505 1050 9506
rect 1022 9479 1023 9505
rect 1023 9479 1049 9505
rect 1049 9479 1050 9505
rect 1022 9478 1050 9479
rect 854 9422 882 9450
rect 1246 9422 1274 9450
rect 5268 9421 5296 9422
rect 5268 9395 5269 9421
rect 5269 9395 5295 9421
rect 5295 9395 5296 9421
rect 5268 9394 5296 9395
rect 5320 9421 5348 9422
rect 5320 9395 5321 9421
rect 5321 9395 5347 9421
rect 5347 9395 5348 9421
rect 5320 9394 5348 9395
rect 5372 9421 5400 9422
rect 5372 9395 5373 9421
rect 5373 9395 5399 9421
rect 5399 9395 5400 9421
rect 5372 9394 5400 9395
rect 1022 9198 1050 9226
rect 8246 9617 8274 9618
rect 8246 9591 8247 9617
rect 8247 9591 8273 9617
rect 8273 9591 8274 9617
rect 8246 9590 8274 9591
rect 8358 9561 8386 9562
rect 8358 9535 8359 9561
rect 8359 9535 8385 9561
rect 8385 9535 8386 9561
rect 8358 9534 8386 9535
rect 8806 9534 8834 9562
rect 9310 9478 9338 9506
rect 9198 9254 9226 9282
rect 8022 9198 8050 9226
rect 8694 9225 8722 9226
rect 8694 9199 8695 9225
rect 8695 9199 8721 9225
rect 8721 9199 8722 9225
rect 8694 9198 8722 9199
rect 854 9086 882 9114
rect 1246 9086 1274 9114
rect 2937 9029 2965 9030
rect 2937 9003 2938 9029
rect 2938 9003 2964 9029
rect 2964 9003 2965 9029
rect 2937 9002 2965 9003
rect 2989 9029 3017 9030
rect 2989 9003 2990 9029
rect 2990 9003 3016 9029
rect 3016 9003 3017 9029
rect 2989 9002 3017 9003
rect 3041 9029 3069 9030
rect 3041 9003 3042 9029
rect 3042 9003 3068 9029
rect 3068 9003 3069 9029
rect 3041 9002 3069 9003
rect 7599 9029 7627 9030
rect 7599 9003 7600 9029
rect 7600 9003 7626 9029
rect 7626 9003 7627 9029
rect 7599 9002 7627 9003
rect 7651 9029 7679 9030
rect 7651 9003 7652 9029
rect 7652 9003 7678 9029
rect 7678 9003 7679 9029
rect 7651 9002 7679 9003
rect 7703 9029 7731 9030
rect 7703 9003 7704 9029
rect 7704 9003 7730 9029
rect 7730 9003 7731 9029
rect 7703 9002 7731 9003
rect 854 8750 882 8778
rect 1246 8750 1274 8778
rect 966 8414 994 8442
rect 1022 8302 1050 8330
rect 1190 8358 1218 8386
rect 1190 8078 1218 8106
rect 1582 8358 1610 8386
rect 5268 8637 5296 8638
rect 5268 8611 5269 8637
rect 5269 8611 5295 8637
rect 5295 8611 5296 8637
rect 5268 8610 5296 8611
rect 5320 8637 5348 8638
rect 5320 8611 5321 8637
rect 5321 8611 5347 8637
rect 5347 8611 5348 8637
rect 5320 8610 5348 8611
rect 5372 8637 5400 8638
rect 5372 8611 5373 8637
rect 5373 8611 5399 8637
rect 5399 8611 5400 8637
rect 5372 8610 5400 8611
rect 2937 8245 2965 8246
rect 2937 8219 2938 8245
rect 2938 8219 2964 8245
rect 2964 8219 2965 8245
rect 2937 8218 2965 8219
rect 2989 8245 3017 8246
rect 2989 8219 2990 8245
rect 2990 8219 3016 8245
rect 3016 8219 3017 8245
rect 2989 8218 3017 8219
rect 3041 8245 3069 8246
rect 3041 8219 3042 8245
rect 3042 8219 3068 8245
rect 3068 8219 3069 8245
rect 3041 8218 3069 8219
rect 7599 8245 7627 8246
rect 7599 8219 7600 8245
rect 7600 8219 7626 8245
rect 7626 8219 7627 8245
rect 7599 8218 7627 8219
rect 7651 8245 7679 8246
rect 7651 8219 7652 8245
rect 7652 8219 7678 8245
rect 7678 8219 7679 8245
rect 7651 8218 7679 8219
rect 7703 8245 7731 8246
rect 7703 8219 7704 8245
rect 7704 8219 7730 8245
rect 7730 8219 7731 8245
rect 7703 8218 7731 8219
rect 2142 8134 2170 8162
rect 7966 8134 7994 8162
rect 1358 8022 1386 8050
rect 7574 7993 7602 7994
rect 7574 7967 7575 7993
rect 7575 7967 7601 7993
rect 7601 7967 7602 7993
rect 7574 7966 7602 7967
rect 7686 7966 7714 7994
rect 1022 7937 1050 7938
rect 1022 7911 1023 7937
rect 1023 7911 1049 7937
rect 1049 7911 1050 7937
rect 1022 7910 1050 7911
rect 5268 7853 5296 7854
rect 5268 7827 5269 7853
rect 5269 7827 5295 7853
rect 5295 7827 5296 7853
rect 5268 7826 5296 7827
rect 5320 7853 5348 7854
rect 5320 7827 5321 7853
rect 5321 7827 5347 7853
rect 5347 7827 5348 7853
rect 5320 7826 5348 7827
rect 5372 7853 5400 7854
rect 5372 7827 5373 7853
rect 5373 7827 5399 7853
rect 5399 7827 5400 7853
rect 5372 7826 5400 7827
rect 910 7769 938 7770
rect 910 7743 911 7769
rect 911 7743 937 7769
rect 937 7743 938 7769
rect 910 7742 938 7743
rect 7966 8049 7994 8050
rect 7966 8023 7967 8049
rect 7967 8023 7993 8049
rect 7993 8023 7994 8049
rect 7966 8022 7994 8023
rect 8638 8302 8666 8330
rect 8302 7993 8330 7994
rect 8302 7967 8303 7993
rect 8303 7967 8329 7993
rect 8329 7967 8330 7993
rect 8302 7966 8330 7967
rect 7742 7686 7770 7714
rect 2937 7461 2965 7462
rect 2937 7435 2938 7461
rect 2938 7435 2964 7461
rect 2964 7435 2965 7461
rect 2937 7434 2965 7435
rect 2989 7461 3017 7462
rect 2989 7435 2990 7461
rect 2990 7435 3016 7461
rect 3016 7435 3017 7461
rect 2989 7434 3017 7435
rect 3041 7461 3069 7462
rect 3041 7435 3042 7461
rect 3042 7435 3068 7461
rect 3068 7435 3069 7461
rect 3041 7434 3069 7435
rect 5268 7069 5296 7070
rect 5268 7043 5269 7069
rect 5269 7043 5295 7069
rect 5295 7043 5296 7069
rect 5268 7042 5296 7043
rect 5320 7069 5348 7070
rect 5320 7043 5321 7069
rect 5321 7043 5347 7069
rect 5347 7043 5348 7069
rect 5320 7042 5348 7043
rect 5372 7069 5400 7070
rect 5372 7043 5373 7069
rect 5373 7043 5399 7069
rect 5399 7043 5400 7069
rect 5372 7042 5400 7043
rect 2937 6677 2965 6678
rect 2937 6651 2938 6677
rect 2938 6651 2964 6677
rect 2964 6651 2965 6677
rect 2937 6650 2965 6651
rect 2989 6677 3017 6678
rect 2989 6651 2990 6677
rect 2990 6651 3016 6677
rect 3016 6651 3017 6677
rect 2989 6650 3017 6651
rect 3041 6677 3069 6678
rect 3041 6651 3042 6677
rect 3042 6651 3068 6677
rect 3068 6651 3069 6677
rect 3041 6650 3069 6651
rect 5268 6285 5296 6286
rect 5268 6259 5269 6285
rect 5269 6259 5295 6285
rect 5295 6259 5296 6285
rect 5268 6258 5296 6259
rect 5320 6285 5348 6286
rect 5320 6259 5321 6285
rect 5321 6259 5347 6285
rect 5347 6259 5348 6285
rect 5320 6258 5348 6259
rect 5372 6285 5400 6286
rect 5372 6259 5373 6285
rect 5373 6259 5399 6285
rect 5399 6259 5400 6285
rect 5372 6258 5400 6259
rect 2937 5893 2965 5894
rect 2937 5867 2938 5893
rect 2938 5867 2964 5893
rect 2964 5867 2965 5893
rect 2937 5866 2965 5867
rect 2989 5893 3017 5894
rect 2989 5867 2990 5893
rect 2990 5867 3016 5893
rect 3016 5867 3017 5893
rect 2989 5866 3017 5867
rect 3041 5893 3069 5894
rect 3041 5867 3042 5893
rect 3042 5867 3068 5893
rect 3068 5867 3069 5893
rect 3041 5866 3069 5867
rect 5268 5501 5296 5502
rect 5268 5475 5269 5501
rect 5269 5475 5295 5501
rect 5295 5475 5296 5501
rect 5268 5474 5296 5475
rect 5320 5501 5348 5502
rect 5320 5475 5321 5501
rect 5321 5475 5347 5501
rect 5347 5475 5348 5501
rect 5320 5474 5348 5475
rect 5372 5501 5400 5502
rect 5372 5475 5373 5501
rect 5373 5475 5399 5501
rect 5399 5475 5400 5501
rect 5372 5474 5400 5475
rect 2937 5109 2965 5110
rect 2937 5083 2938 5109
rect 2938 5083 2964 5109
rect 2964 5083 2965 5109
rect 2937 5082 2965 5083
rect 2989 5109 3017 5110
rect 2989 5083 2990 5109
rect 2990 5083 3016 5109
rect 3016 5083 3017 5109
rect 2989 5082 3017 5083
rect 3041 5109 3069 5110
rect 3041 5083 3042 5109
rect 3042 5083 3068 5109
rect 3068 5083 3069 5109
rect 3041 5082 3069 5083
rect 5268 4717 5296 4718
rect 5268 4691 5269 4717
rect 5269 4691 5295 4717
rect 5295 4691 5296 4717
rect 5268 4690 5296 4691
rect 5320 4717 5348 4718
rect 5320 4691 5321 4717
rect 5321 4691 5347 4717
rect 5347 4691 5348 4717
rect 5320 4690 5348 4691
rect 5372 4717 5400 4718
rect 5372 4691 5373 4717
rect 5373 4691 5399 4717
rect 5399 4691 5400 4717
rect 5372 4690 5400 4691
rect 2937 4325 2965 4326
rect 2937 4299 2938 4325
rect 2938 4299 2964 4325
rect 2964 4299 2965 4325
rect 2937 4298 2965 4299
rect 2989 4325 3017 4326
rect 2989 4299 2990 4325
rect 2990 4299 3016 4325
rect 3016 4299 3017 4325
rect 2989 4298 3017 4299
rect 3041 4325 3069 4326
rect 3041 4299 3042 4325
rect 3042 4299 3068 4325
rect 3068 4299 3069 4325
rect 3041 4298 3069 4299
rect 5268 3933 5296 3934
rect 5268 3907 5269 3933
rect 5269 3907 5295 3933
rect 5295 3907 5296 3933
rect 5268 3906 5296 3907
rect 5320 3933 5348 3934
rect 5320 3907 5321 3933
rect 5321 3907 5347 3933
rect 5347 3907 5348 3933
rect 5320 3906 5348 3907
rect 5372 3933 5400 3934
rect 5372 3907 5373 3933
rect 5373 3907 5399 3933
rect 5399 3907 5400 3933
rect 5372 3906 5400 3907
rect 2937 3541 2965 3542
rect 2937 3515 2938 3541
rect 2938 3515 2964 3541
rect 2964 3515 2965 3541
rect 2937 3514 2965 3515
rect 2989 3541 3017 3542
rect 2989 3515 2990 3541
rect 2990 3515 3016 3541
rect 3016 3515 3017 3541
rect 2989 3514 3017 3515
rect 3041 3541 3069 3542
rect 3041 3515 3042 3541
rect 3042 3515 3068 3541
rect 3068 3515 3069 3541
rect 3041 3514 3069 3515
rect 5268 3149 5296 3150
rect 5268 3123 5269 3149
rect 5269 3123 5295 3149
rect 5295 3123 5296 3149
rect 5268 3122 5296 3123
rect 5320 3149 5348 3150
rect 5320 3123 5321 3149
rect 5321 3123 5347 3149
rect 5347 3123 5348 3149
rect 5320 3122 5348 3123
rect 5372 3149 5400 3150
rect 5372 3123 5373 3149
rect 5373 3123 5399 3149
rect 5399 3123 5400 3149
rect 5372 3122 5400 3123
rect 2937 2757 2965 2758
rect 2937 2731 2938 2757
rect 2938 2731 2964 2757
rect 2964 2731 2965 2757
rect 2937 2730 2965 2731
rect 2989 2757 3017 2758
rect 2989 2731 2990 2757
rect 2990 2731 3016 2757
rect 3016 2731 3017 2757
rect 2989 2730 3017 2731
rect 3041 2757 3069 2758
rect 3041 2731 3042 2757
rect 3042 2731 3068 2757
rect 3068 2731 3069 2757
rect 3041 2730 3069 2731
rect 5268 2365 5296 2366
rect 5268 2339 5269 2365
rect 5269 2339 5295 2365
rect 5295 2339 5296 2365
rect 5268 2338 5296 2339
rect 5320 2365 5348 2366
rect 5320 2339 5321 2365
rect 5321 2339 5347 2365
rect 5347 2339 5348 2365
rect 5320 2338 5348 2339
rect 5372 2365 5400 2366
rect 5372 2339 5373 2365
rect 5373 2339 5399 2365
rect 5399 2339 5400 2365
rect 5372 2338 5400 2339
rect 6510 2113 6538 2114
rect 6510 2087 6511 2113
rect 6511 2087 6537 2113
rect 6537 2087 6538 2113
rect 6510 2086 6538 2087
rect 7599 7461 7627 7462
rect 7599 7435 7600 7461
rect 7600 7435 7626 7461
rect 7626 7435 7627 7461
rect 7599 7434 7627 7435
rect 7651 7461 7679 7462
rect 7651 7435 7652 7461
rect 7652 7435 7678 7461
rect 7678 7435 7679 7461
rect 7651 7434 7679 7435
rect 7703 7461 7731 7462
rect 7703 7435 7704 7461
rect 7704 7435 7730 7461
rect 7730 7435 7731 7461
rect 7703 7434 7731 7435
rect 7294 2254 7322 2282
rect 7350 7182 7378 7210
rect 7599 6677 7627 6678
rect 7599 6651 7600 6677
rect 7600 6651 7626 6677
rect 7626 6651 7627 6677
rect 7599 6650 7627 6651
rect 7651 6677 7679 6678
rect 7651 6651 7652 6677
rect 7652 6651 7678 6677
rect 7678 6651 7679 6677
rect 7651 6650 7679 6651
rect 7703 6677 7731 6678
rect 7703 6651 7704 6677
rect 7704 6651 7730 6677
rect 7730 6651 7731 6677
rect 7703 6650 7731 6651
rect 7854 6006 7882 6034
rect 7599 5893 7627 5894
rect 7599 5867 7600 5893
rect 7600 5867 7626 5893
rect 7626 5867 7627 5893
rect 7599 5866 7627 5867
rect 7651 5893 7679 5894
rect 7651 5867 7652 5893
rect 7652 5867 7678 5893
rect 7678 5867 7679 5893
rect 7651 5866 7679 5867
rect 7703 5893 7731 5894
rect 7703 5867 7704 5893
rect 7704 5867 7730 5893
rect 7730 5867 7731 5893
rect 7703 5866 7731 5867
rect 7599 5109 7627 5110
rect 7599 5083 7600 5109
rect 7600 5083 7626 5109
rect 7626 5083 7627 5109
rect 7599 5082 7627 5083
rect 7651 5109 7679 5110
rect 7651 5083 7652 5109
rect 7652 5083 7678 5109
rect 7678 5083 7679 5109
rect 7651 5082 7679 5083
rect 7703 5109 7731 5110
rect 7703 5083 7704 5109
rect 7704 5083 7730 5109
rect 7730 5083 7731 5109
rect 7703 5082 7731 5083
rect 7599 4325 7627 4326
rect 7599 4299 7600 4325
rect 7600 4299 7626 4325
rect 7626 4299 7627 4325
rect 7599 4298 7627 4299
rect 7651 4325 7679 4326
rect 7651 4299 7652 4325
rect 7652 4299 7678 4325
rect 7678 4299 7679 4325
rect 7651 4298 7679 4299
rect 7703 4325 7731 4326
rect 7703 4299 7704 4325
rect 7704 4299 7730 4325
rect 7730 4299 7731 4325
rect 7703 4298 7731 4299
rect 7599 3541 7627 3542
rect 7599 3515 7600 3541
rect 7600 3515 7626 3541
rect 7626 3515 7627 3541
rect 7599 3514 7627 3515
rect 7651 3541 7679 3542
rect 7651 3515 7652 3541
rect 7652 3515 7678 3541
rect 7678 3515 7679 3541
rect 7651 3514 7679 3515
rect 7703 3541 7731 3542
rect 7703 3515 7704 3541
rect 7704 3515 7730 3541
rect 7730 3515 7731 3541
rect 7703 3514 7731 3515
rect 7599 2757 7627 2758
rect 7599 2731 7600 2757
rect 7600 2731 7626 2757
rect 7626 2731 7627 2757
rect 7599 2730 7627 2731
rect 7651 2757 7679 2758
rect 7651 2731 7652 2757
rect 7652 2731 7678 2757
rect 7678 2731 7679 2757
rect 7651 2730 7679 2731
rect 7703 2757 7731 2758
rect 7703 2731 7704 2757
rect 7704 2731 7730 2757
rect 7730 2731 7731 2757
rect 7703 2730 7731 2731
rect 8246 7686 8274 7714
rect 6846 2086 6874 2114
rect 2937 1973 2965 1974
rect 2937 1947 2938 1973
rect 2938 1947 2964 1973
rect 2964 1947 2965 1973
rect 2937 1946 2965 1947
rect 2989 1973 3017 1974
rect 2989 1947 2990 1973
rect 2990 1947 3016 1973
rect 3016 1947 3017 1973
rect 2989 1946 3017 1947
rect 3041 1973 3069 1974
rect 3041 1947 3042 1973
rect 3042 1947 3068 1973
rect 3068 1947 3069 1973
rect 3041 1946 3069 1947
rect 5268 1581 5296 1582
rect 5268 1555 5269 1581
rect 5269 1555 5295 1581
rect 5295 1555 5296 1581
rect 5268 1554 5296 1555
rect 5320 1581 5348 1582
rect 5320 1555 5321 1581
rect 5321 1555 5347 1581
rect 5347 1555 5348 1581
rect 5320 1554 5348 1555
rect 5372 1581 5400 1582
rect 5372 1555 5373 1581
rect 5373 1555 5399 1581
rect 5399 1555 5400 1581
rect 5372 1554 5400 1555
rect 7599 1973 7627 1974
rect 7599 1947 7600 1973
rect 7600 1947 7626 1973
rect 7626 1947 7627 1973
rect 7599 1946 7627 1947
rect 7651 1973 7679 1974
rect 7651 1947 7652 1973
rect 7652 1947 7678 1973
rect 7678 1947 7679 1973
rect 7651 1946 7679 1947
rect 7703 1973 7731 1974
rect 7703 1947 7704 1973
rect 7704 1947 7730 1973
rect 7730 1947 7731 1973
rect 7703 1946 7731 1947
rect 7798 1777 7826 1778
rect 7798 1751 7799 1777
rect 7799 1751 7825 1777
rect 7825 1751 7826 1777
rect 7798 1750 7826 1751
rect 8022 1721 8050 1722
rect 8022 1695 8023 1721
rect 8023 1695 8049 1721
rect 8049 1695 8050 1721
rect 8022 1694 8050 1695
rect 8414 6006 8442 6034
rect 9926 9673 9954 9674
rect 9926 9647 9927 9673
rect 9927 9647 9953 9673
rect 9953 9647 9954 9673
rect 9926 9646 9954 9647
rect 14592 13341 14620 13342
rect 14592 13315 14593 13341
rect 14593 13315 14619 13341
rect 14619 13315 14620 13341
rect 14592 13314 14620 13315
rect 14644 13341 14672 13342
rect 14644 13315 14645 13341
rect 14645 13315 14671 13341
rect 14671 13315 14672 13341
rect 14644 13314 14672 13315
rect 14696 13341 14724 13342
rect 14696 13315 14697 13341
rect 14697 13315 14723 13341
rect 14723 13315 14724 13341
rect 14696 13314 14724 13315
rect 19254 13341 19282 13342
rect 19254 13315 19255 13341
rect 19255 13315 19281 13341
rect 19281 13315 19282 13341
rect 19254 13314 19282 13315
rect 19306 13341 19334 13342
rect 19306 13315 19307 13341
rect 19307 13315 19333 13341
rect 19333 13315 19334 13341
rect 19306 13314 19334 13315
rect 19358 13341 19386 13342
rect 19358 13315 19359 13341
rect 19359 13315 19385 13341
rect 19385 13315 19386 13341
rect 19358 13314 19386 13315
rect 12261 12949 12289 12950
rect 12261 12923 12262 12949
rect 12262 12923 12288 12949
rect 12288 12923 12289 12949
rect 12261 12922 12289 12923
rect 12313 12949 12341 12950
rect 12313 12923 12314 12949
rect 12314 12923 12340 12949
rect 12340 12923 12341 12949
rect 12313 12922 12341 12923
rect 12365 12949 12393 12950
rect 12365 12923 12366 12949
rect 12366 12923 12392 12949
rect 12392 12923 12393 12949
rect 12365 12922 12393 12923
rect 16923 12949 16951 12950
rect 16923 12923 16924 12949
rect 16924 12923 16950 12949
rect 16950 12923 16951 12949
rect 16923 12922 16951 12923
rect 16975 12949 17003 12950
rect 16975 12923 16976 12949
rect 16976 12923 17002 12949
rect 17002 12923 17003 12949
rect 16975 12922 17003 12923
rect 17027 12949 17055 12950
rect 17027 12923 17028 12949
rect 17028 12923 17054 12949
rect 17054 12923 17055 12949
rect 17027 12922 17055 12923
rect 14592 12557 14620 12558
rect 14592 12531 14593 12557
rect 14593 12531 14619 12557
rect 14619 12531 14620 12557
rect 14592 12530 14620 12531
rect 14644 12557 14672 12558
rect 14644 12531 14645 12557
rect 14645 12531 14671 12557
rect 14671 12531 14672 12557
rect 14644 12530 14672 12531
rect 14696 12557 14724 12558
rect 14696 12531 14697 12557
rect 14697 12531 14723 12557
rect 14723 12531 14724 12557
rect 14696 12530 14724 12531
rect 19254 12557 19282 12558
rect 19254 12531 19255 12557
rect 19255 12531 19281 12557
rect 19281 12531 19282 12557
rect 19254 12530 19282 12531
rect 19306 12557 19334 12558
rect 19306 12531 19307 12557
rect 19307 12531 19333 12557
rect 19333 12531 19334 12557
rect 19306 12530 19334 12531
rect 19358 12557 19386 12558
rect 19358 12531 19359 12557
rect 19359 12531 19385 12557
rect 19385 12531 19386 12557
rect 19358 12530 19386 12531
rect 11214 12334 11242 12362
rect 17822 12361 17850 12362
rect 17822 12335 17823 12361
rect 17823 12335 17849 12361
rect 17849 12335 17850 12361
rect 17822 12334 17850 12335
rect 12261 12165 12289 12166
rect 12261 12139 12262 12165
rect 12262 12139 12288 12165
rect 12288 12139 12289 12165
rect 12261 12138 12289 12139
rect 12313 12165 12341 12166
rect 12313 12139 12314 12165
rect 12314 12139 12340 12165
rect 12340 12139 12341 12165
rect 12313 12138 12341 12139
rect 12365 12165 12393 12166
rect 12365 12139 12366 12165
rect 12366 12139 12392 12165
rect 12392 12139 12393 12165
rect 12365 12138 12393 12139
rect 16923 12165 16951 12166
rect 16923 12139 16924 12165
rect 16924 12139 16950 12165
rect 16950 12139 16951 12165
rect 16923 12138 16951 12139
rect 16975 12165 17003 12166
rect 16975 12139 16976 12165
rect 16976 12139 17002 12165
rect 17002 12139 17003 12165
rect 16975 12138 17003 12139
rect 17027 12165 17055 12166
rect 17027 12139 17028 12165
rect 17028 12139 17054 12165
rect 17054 12139 17055 12165
rect 17027 12138 17055 12139
rect 18998 12110 19026 12138
rect 18830 11857 18858 11858
rect 18830 11831 18831 11857
rect 18831 11831 18857 11857
rect 18857 11831 18858 11857
rect 18830 11830 18858 11831
rect 14592 11773 14620 11774
rect 14592 11747 14593 11773
rect 14593 11747 14619 11773
rect 14619 11747 14620 11773
rect 14592 11746 14620 11747
rect 14644 11773 14672 11774
rect 14644 11747 14645 11773
rect 14645 11747 14671 11773
rect 14671 11747 14672 11773
rect 14644 11746 14672 11747
rect 14696 11773 14724 11774
rect 14696 11747 14697 11773
rect 14697 11747 14723 11773
rect 14723 11747 14724 11773
rect 14696 11746 14724 11747
rect 12054 11606 12082 11634
rect 11158 10766 11186 10794
rect 11214 10878 11242 10906
rect 11606 10793 11634 10794
rect 11606 10767 11607 10793
rect 11607 10767 11633 10793
rect 11633 10767 11634 10793
rect 11606 10766 11634 10767
rect 18830 11438 18858 11466
rect 12261 11381 12289 11382
rect 12261 11355 12262 11381
rect 12262 11355 12288 11381
rect 12288 11355 12289 11381
rect 12261 11354 12289 11355
rect 12313 11381 12341 11382
rect 12313 11355 12314 11381
rect 12314 11355 12340 11381
rect 12340 11355 12341 11381
rect 12313 11354 12341 11355
rect 12365 11381 12393 11382
rect 12365 11355 12366 11381
rect 12366 11355 12392 11381
rect 12392 11355 12393 11381
rect 12365 11354 12393 11355
rect 16923 11381 16951 11382
rect 16923 11355 16924 11381
rect 16924 11355 16950 11381
rect 16950 11355 16951 11381
rect 16923 11354 16951 11355
rect 16975 11381 17003 11382
rect 16975 11355 16976 11381
rect 16976 11355 17002 11381
rect 17002 11355 17003 11381
rect 16975 11354 17003 11355
rect 17027 11381 17055 11382
rect 17027 11355 17028 11381
rect 17028 11355 17054 11381
rect 17054 11355 17055 11381
rect 17027 11354 17055 11355
rect 18830 11129 18858 11130
rect 18830 11103 18831 11129
rect 18831 11103 18857 11129
rect 18857 11103 18858 11129
rect 18830 11102 18858 11103
rect 17822 11046 17850 11074
rect 14592 10989 14620 10990
rect 14592 10963 14593 10989
rect 14593 10963 14619 10989
rect 14619 10963 14620 10989
rect 14592 10962 14620 10963
rect 14644 10989 14672 10990
rect 14644 10963 14645 10989
rect 14645 10963 14671 10989
rect 14671 10963 14672 10989
rect 14644 10962 14672 10963
rect 14696 10989 14724 10990
rect 14696 10963 14697 10989
rect 14697 10963 14723 10989
rect 14723 10963 14724 10989
rect 14696 10962 14724 10963
rect 12261 10597 12289 10598
rect 12261 10571 12262 10597
rect 12262 10571 12288 10597
rect 12288 10571 12289 10597
rect 12261 10570 12289 10571
rect 12313 10597 12341 10598
rect 12313 10571 12314 10597
rect 12314 10571 12340 10597
rect 12340 10571 12341 10597
rect 12313 10570 12341 10571
rect 12365 10597 12393 10598
rect 12365 10571 12366 10597
rect 12366 10571 12392 10597
rect 12392 10571 12393 10597
rect 12365 10570 12393 10571
rect 16923 10597 16951 10598
rect 16923 10571 16924 10597
rect 16924 10571 16950 10597
rect 16950 10571 16951 10597
rect 16923 10570 16951 10571
rect 16975 10597 17003 10598
rect 16975 10571 16976 10597
rect 16976 10571 17002 10597
rect 17002 10571 17003 10597
rect 16975 10570 17003 10571
rect 17027 10597 17055 10598
rect 17027 10571 17028 10597
rect 17028 10571 17054 10597
rect 17054 10571 17055 10597
rect 17027 10570 17055 10571
rect 18270 10457 18298 10458
rect 18270 10431 18271 10457
rect 18271 10431 18297 10457
rect 18297 10431 18298 10457
rect 18270 10430 18298 10431
rect 11718 10401 11746 10402
rect 11718 10375 11719 10401
rect 11719 10375 11745 10401
rect 11745 10375 11746 10401
rect 11718 10374 11746 10375
rect 19110 11830 19138 11858
rect 19254 11773 19282 11774
rect 19254 11747 19255 11773
rect 19255 11747 19281 11773
rect 19281 11747 19282 11773
rect 19254 11746 19282 11747
rect 19306 11773 19334 11774
rect 19306 11747 19307 11773
rect 19307 11747 19333 11773
rect 19333 11747 19334 11773
rect 19306 11746 19334 11747
rect 19358 11773 19386 11774
rect 19358 11747 19359 11773
rect 19359 11747 19385 11773
rect 19385 11747 19386 11773
rect 19358 11746 19386 11747
rect 18942 11633 18970 11634
rect 18942 11607 18943 11633
rect 18943 11607 18969 11633
rect 18969 11607 18970 11633
rect 18942 11606 18970 11607
rect 19110 11438 19138 11466
rect 19110 11129 19138 11130
rect 19110 11103 19111 11129
rect 19111 11103 19137 11129
rect 19137 11103 19138 11129
rect 19110 11102 19138 11103
rect 19254 10989 19282 10990
rect 19254 10963 19255 10989
rect 19255 10963 19281 10989
rect 19281 10963 19282 10989
rect 19254 10962 19282 10963
rect 19306 10989 19334 10990
rect 19306 10963 19307 10989
rect 19307 10963 19333 10989
rect 19333 10963 19334 10989
rect 19306 10962 19334 10963
rect 19358 10989 19386 10990
rect 19358 10963 19359 10989
rect 19359 10963 19385 10989
rect 19385 10963 19386 10989
rect 19358 10962 19386 10963
rect 18942 10878 18970 10906
rect 18998 10766 19026 10794
rect 18886 10374 18914 10402
rect 19110 10430 19138 10458
rect 12222 10318 12250 10346
rect 14592 10205 14620 10206
rect 14592 10179 14593 10205
rect 14593 10179 14619 10205
rect 14619 10179 14620 10205
rect 14592 10178 14620 10179
rect 14644 10205 14672 10206
rect 14644 10179 14645 10205
rect 14645 10179 14671 10205
rect 14671 10179 14672 10205
rect 14644 10178 14672 10179
rect 14696 10205 14724 10206
rect 14696 10179 14697 10205
rect 14697 10179 14723 10205
rect 14723 10179 14724 10205
rect 14696 10178 14724 10179
rect 10822 9646 10850 9674
rect 10094 9505 10122 9506
rect 10094 9479 10095 9505
rect 10095 9479 10121 9505
rect 10121 9479 10122 9505
rect 10094 9478 10122 9479
rect 10262 9505 10290 9506
rect 10262 9479 10263 9505
rect 10263 9479 10289 9505
rect 10289 9479 10290 9505
rect 10262 9478 10290 9479
rect 9930 9421 9958 9422
rect 9930 9395 9931 9421
rect 9931 9395 9957 9421
rect 9957 9395 9958 9421
rect 9930 9394 9958 9395
rect 9982 9421 10010 9422
rect 9982 9395 9983 9421
rect 9983 9395 10009 9421
rect 10009 9395 10010 9421
rect 9982 9394 10010 9395
rect 10034 9421 10062 9422
rect 10034 9395 10035 9421
rect 10035 9395 10061 9421
rect 10061 9395 10062 9421
rect 10034 9394 10062 9395
rect 9646 9254 9674 9282
rect 9366 9198 9394 9226
rect 18942 10345 18970 10346
rect 18942 10319 18943 10345
rect 18943 10319 18969 10345
rect 18969 10319 18970 10345
rect 18942 10318 18970 10319
rect 19254 10205 19282 10206
rect 19254 10179 19255 10205
rect 19255 10179 19281 10205
rect 19281 10179 19282 10205
rect 19254 10178 19282 10179
rect 19306 10205 19334 10206
rect 19306 10179 19307 10205
rect 19307 10179 19333 10205
rect 19333 10179 19334 10205
rect 19306 10178 19334 10179
rect 19358 10205 19386 10206
rect 19358 10179 19359 10205
rect 19359 10179 19385 10205
rect 19385 10179 19386 10205
rect 19358 10178 19386 10179
rect 18830 10121 18858 10122
rect 18830 10095 18831 10121
rect 18831 10095 18857 10121
rect 18857 10095 18858 10121
rect 18830 10094 18858 10095
rect 12261 9813 12289 9814
rect 12261 9787 12262 9813
rect 12262 9787 12288 9813
rect 12288 9787 12289 9813
rect 12261 9786 12289 9787
rect 12313 9813 12341 9814
rect 12313 9787 12314 9813
rect 12314 9787 12340 9813
rect 12340 9787 12341 9813
rect 12313 9786 12341 9787
rect 12365 9813 12393 9814
rect 12365 9787 12366 9813
rect 12366 9787 12392 9813
rect 12392 9787 12393 9813
rect 12365 9786 12393 9787
rect 16923 9813 16951 9814
rect 16923 9787 16924 9813
rect 16924 9787 16950 9813
rect 16950 9787 16951 9813
rect 16923 9786 16951 9787
rect 16975 9813 17003 9814
rect 16975 9787 16976 9813
rect 16976 9787 17002 9813
rect 17002 9787 17003 9813
rect 16975 9786 17003 9787
rect 17027 9813 17055 9814
rect 17027 9787 17028 9813
rect 17028 9787 17054 9813
rect 17054 9787 17055 9813
rect 17027 9786 17055 9787
rect 11270 9478 11298 9506
rect 10598 9169 10626 9170
rect 10598 9143 10599 9169
rect 10599 9143 10625 9169
rect 10625 9143 10626 9169
rect 10598 9142 10626 9143
rect 8862 7686 8890 7714
rect 8750 7209 8778 7210
rect 8750 7183 8751 7209
rect 8751 7183 8777 7209
rect 8777 7183 8778 7209
rect 8750 7182 8778 7183
rect 9254 7910 9282 7938
rect 8190 2281 8218 2282
rect 8190 2255 8191 2281
rect 8191 2255 8217 2281
rect 8217 2255 8218 2281
rect 8190 2254 8218 2255
rect 8134 1750 8162 1778
rect 8358 1694 8386 1722
rect 9310 7686 9338 7714
rect 11046 8918 11074 8946
rect 10654 8777 10682 8778
rect 10654 8751 10655 8777
rect 10655 8751 10681 8777
rect 10681 8751 10682 8777
rect 10654 8750 10682 8751
rect 9930 8637 9958 8638
rect 9930 8611 9931 8637
rect 9931 8611 9957 8637
rect 9957 8611 9958 8637
rect 9930 8610 9958 8611
rect 9982 8637 10010 8638
rect 9982 8611 9983 8637
rect 9983 8611 10009 8637
rect 10009 8611 10010 8637
rect 9982 8610 10010 8611
rect 10034 8637 10062 8638
rect 10034 8611 10035 8637
rect 10035 8611 10061 8637
rect 10061 8611 10062 8637
rect 10034 8610 10062 8611
rect 11102 8358 11130 8386
rect 9478 7966 9506 7994
rect 10038 7937 10066 7938
rect 10038 7911 10039 7937
rect 10039 7911 10065 7937
rect 10065 7911 10066 7937
rect 10038 7910 10066 7911
rect 10206 7937 10234 7938
rect 10206 7911 10207 7937
rect 10207 7911 10233 7937
rect 10233 7911 10234 7937
rect 10206 7910 10234 7911
rect 9930 7853 9958 7854
rect 9930 7827 9931 7853
rect 9931 7827 9957 7853
rect 9957 7827 9958 7853
rect 9930 7826 9958 7827
rect 9982 7853 10010 7854
rect 9982 7827 9983 7853
rect 9983 7827 10009 7853
rect 10009 7827 10010 7853
rect 9982 7826 10010 7827
rect 10034 7853 10062 7854
rect 10034 7827 10035 7853
rect 10035 7827 10061 7853
rect 10061 7827 10062 7853
rect 10034 7826 10062 7827
rect 9870 7742 9898 7770
rect 9478 7630 9506 7658
rect 9422 2254 9450 2282
rect 9870 7657 9898 7658
rect 9870 7631 9871 7657
rect 9871 7631 9897 7657
rect 9897 7631 9898 7657
rect 9870 7630 9898 7631
rect 9930 7069 9958 7070
rect 9930 7043 9931 7069
rect 9931 7043 9957 7069
rect 9957 7043 9958 7069
rect 9930 7042 9958 7043
rect 9982 7069 10010 7070
rect 9982 7043 9983 7069
rect 9983 7043 10009 7069
rect 10009 7043 10010 7069
rect 9982 7042 10010 7043
rect 10034 7069 10062 7070
rect 10034 7043 10035 7069
rect 10035 7043 10061 7069
rect 10061 7043 10062 7069
rect 10034 7042 10062 7043
rect 9930 6285 9958 6286
rect 9930 6259 9931 6285
rect 9931 6259 9957 6285
rect 9957 6259 9958 6285
rect 9930 6258 9958 6259
rect 9982 6285 10010 6286
rect 9982 6259 9983 6285
rect 9983 6259 10009 6285
rect 10009 6259 10010 6285
rect 9982 6258 10010 6259
rect 10034 6285 10062 6286
rect 10034 6259 10035 6285
rect 10035 6259 10061 6285
rect 10061 6259 10062 6285
rect 10034 6258 10062 6259
rect 10318 5894 10346 5922
rect 9930 5501 9958 5502
rect 9930 5475 9931 5501
rect 9931 5475 9957 5501
rect 9957 5475 9958 5501
rect 9930 5474 9958 5475
rect 9982 5501 10010 5502
rect 9982 5475 9983 5501
rect 9983 5475 10009 5501
rect 10009 5475 10010 5501
rect 9982 5474 10010 5475
rect 10034 5501 10062 5502
rect 10034 5475 10035 5501
rect 10035 5475 10061 5501
rect 10061 5475 10062 5501
rect 10034 5474 10062 5475
rect 9930 4717 9958 4718
rect 9930 4691 9931 4717
rect 9931 4691 9957 4717
rect 9957 4691 9958 4717
rect 9930 4690 9958 4691
rect 9982 4717 10010 4718
rect 9982 4691 9983 4717
rect 9983 4691 10009 4717
rect 10009 4691 10010 4717
rect 9982 4690 10010 4691
rect 10034 4717 10062 4718
rect 10034 4691 10035 4717
rect 10035 4691 10061 4717
rect 10061 4691 10062 4717
rect 10034 4690 10062 4691
rect 9930 3933 9958 3934
rect 9930 3907 9931 3933
rect 9931 3907 9957 3933
rect 9957 3907 9958 3933
rect 9930 3906 9958 3907
rect 9982 3933 10010 3934
rect 9982 3907 9983 3933
rect 9983 3907 10009 3933
rect 10009 3907 10010 3933
rect 9982 3906 10010 3907
rect 10034 3933 10062 3934
rect 10034 3907 10035 3933
rect 10035 3907 10061 3933
rect 10061 3907 10062 3933
rect 10034 3906 10062 3907
rect 9930 3149 9958 3150
rect 9930 3123 9931 3149
rect 9931 3123 9957 3149
rect 9957 3123 9958 3149
rect 9930 3122 9958 3123
rect 9982 3149 10010 3150
rect 9982 3123 9983 3149
rect 9983 3123 10009 3149
rect 10009 3123 10010 3149
rect 9982 3122 10010 3123
rect 10034 3149 10062 3150
rect 10034 3123 10035 3149
rect 10035 3123 10061 3149
rect 10061 3123 10062 3149
rect 10034 3122 10062 3123
rect 9870 2478 9898 2506
rect 9930 2365 9958 2366
rect 9930 2339 9931 2365
rect 9931 2339 9957 2365
rect 9957 2339 9958 2365
rect 9930 2338 9958 2339
rect 9982 2365 10010 2366
rect 9982 2339 9983 2365
rect 9983 2339 10009 2365
rect 10009 2339 10010 2365
rect 9982 2338 10010 2339
rect 10034 2365 10062 2366
rect 10034 2339 10035 2365
rect 10035 2339 10061 2365
rect 10061 2339 10062 2365
rect 10034 2338 10062 2339
rect 9926 2254 9954 2282
rect 9930 1581 9958 1582
rect 9930 1555 9931 1581
rect 9931 1555 9957 1581
rect 9957 1555 9958 1581
rect 9930 1554 9958 1555
rect 9982 1581 10010 1582
rect 9982 1555 9983 1581
rect 9983 1555 10009 1581
rect 10009 1555 10010 1581
rect 9982 1554 10010 1555
rect 10034 1581 10062 1582
rect 10034 1555 10035 1581
rect 10035 1555 10061 1581
rect 10061 1555 10062 1581
rect 10034 1554 10062 1555
rect 11662 9310 11690 9338
rect 12166 9478 12194 9506
rect 11718 9225 11746 9226
rect 11718 9199 11719 9225
rect 11719 9199 11745 9225
rect 11745 9199 11746 9225
rect 11718 9198 11746 9199
rect 14592 9421 14620 9422
rect 14592 9395 14593 9421
rect 14593 9395 14619 9421
rect 14619 9395 14620 9421
rect 14592 9394 14620 9395
rect 14644 9421 14672 9422
rect 14644 9395 14645 9421
rect 14645 9395 14671 9421
rect 14671 9395 14672 9421
rect 14644 9394 14672 9395
rect 14696 9421 14724 9422
rect 14696 9395 14697 9421
rect 14697 9395 14723 9421
rect 14723 9395 14724 9421
rect 14696 9394 14724 9395
rect 17822 9310 17850 9338
rect 12670 9169 12698 9170
rect 12670 9143 12671 9169
rect 12671 9143 12697 9169
rect 12697 9143 12698 9169
rect 12670 9142 12698 9143
rect 12261 9029 12289 9030
rect 12261 9003 12262 9029
rect 12262 9003 12288 9029
rect 12288 9003 12289 9029
rect 12261 9002 12289 9003
rect 12313 9029 12341 9030
rect 12313 9003 12314 9029
rect 12314 9003 12340 9029
rect 12340 9003 12341 9029
rect 12313 9002 12341 9003
rect 12365 9029 12393 9030
rect 12365 9003 12366 9029
rect 12366 9003 12392 9029
rect 12392 9003 12393 9029
rect 12365 9002 12393 9003
rect 16923 9029 16951 9030
rect 16923 9003 16924 9029
rect 16924 9003 16950 9029
rect 16950 9003 16951 9029
rect 16923 9002 16951 9003
rect 16975 9029 17003 9030
rect 16975 9003 16976 9029
rect 16976 9003 17002 9029
rect 17002 9003 17003 9029
rect 16975 9002 17003 9003
rect 17027 9029 17055 9030
rect 17027 9003 17028 9029
rect 17028 9003 17054 9029
rect 17054 9003 17055 9029
rect 17027 9002 17055 9003
rect 12950 8918 12978 8946
rect 12222 8862 12250 8890
rect 11718 8833 11746 8834
rect 11718 8807 11719 8833
rect 11719 8807 11745 8833
rect 11745 8807 11746 8833
rect 11718 8806 11746 8807
rect 14592 8637 14620 8638
rect 14592 8611 14593 8637
rect 14593 8611 14619 8637
rect 14619 8611 14620 8637
rect 14592 8610 14620 8611
rect 14644 8637 14672 8638
rect 14644 8611 14645 8637
rect 14645 8611 14671 8637
rect 14671 8611 14672 8637
rect 14644 8610 14672 8611
rect 14696 8637 14724 8638
rect 14696 8611 14697 8637
rect 14697 8611 14723 8637
rect 14723 8611 14724 8637
rect 14696 8610 14724 8611
rect 12261 8245 12289 8246
rect 12261 8219 12262 8245
rect 12262 8219 12288 8245
rect 12288 8219 12289 8245
rect 12261 8218 12289 8219
rect 12313 8245 12341 8246
rect 12313 8219 12314 8245
rect 12314 8219 12340 8245
rect 12340 8219 12341 8245
rect 12313 8218 12341 8219
rect 12365 8245 12393 8246
rect 12365 8219 12366 8245
rect 12366 8219 12392 8245
rect 12392 8219 12393 8245
rect 12365 8218 12393 8219
rect 16923 8245 16951 8246
rect 16923 8219 16924 8245
rect 16924 8219 16950 8245
rect 16950 8219 16951 8245
rect 16923 8218 16951 8219
rect 16975 8245 17003 8246
rect 16975 8219 16976 8245
rect 16976 8219 17002 8245
rect 17002 8219 17003 8245
rect 16975 8218 17003 8219
rect 17027 8245 17055 8246
rect 17027 8219 17028 8245
rect 17028 8219 17054 8245
rect 17054 8219 17055 8245
rect 17027 8218 17055 8219
rect 12614 7910 12642 7938
rect 11550 6790 11578 6818
rect 12166 7742 12194 7770
rect 11214 5894 11242 5922
rect 10766 1694 10794 1722
rect 10990 1694 11018 1722
rect 11382 2478 11410 2506
rect 12110 2030 12138 2058
rect 11774 1806 11802 1834
rect 12261 7461 12289 7462
rect 12261 7435 12262 7461
rect 12262 7435 12288 7461
rect 12288 7435 12289 7461
rect 12261 7434 12289 7435
rect 12313 7461 12341 7462
rect 12313 7435 12314 7461
rect 12314 7435 12340 7461
rect 12340 7435 12341 7461
rect 12313 7434 12341 7435
rect 12365 7461 12393 7462
rect 12365 7435 12366 7461
rect 12366 7435 12392 7461
rect 12392 7435 12393 7461
rect 12365 7434 12393 7435
rect 12261 6677 12289 6678
rect 12261 6651 12262 6677
rect 12262 6651 12288 6677
rect 12288 6651 12289 6677
rect 12261 6650 12289 6651
rect 12313 6677 12341 6678
rect 12313 6651 12314 6677
rect 12314 6651 12340 6677
rect 12340 6651 12341 6677
rect 12313 6650 12341 6651
rect 12365 6677 12393 6678
rect 12365 6651 12366 6677
rect 12366 6651 12392 6677
rect 12392 6651 12393 6677
rect 12365 6650 12393 6651
rect 12261 5893 12289 5894
rect 12261 5867 12262 5893
rect 12262 5867 12288 5893
rect 12288 5867 12289 5893
rect 12261 5866 12289 5867
rect 12313 5893 12341 5894
rect 12313 5867 12314 5893
rect 12314 5867 12340 5893
rect 12340 5867 12341 5893
rect 12313 5866 12341 5867
rect 12365 5893 12393 5894
rect 12365 5867 12366 5893
rect 12366 5867 12392 5893
rect 12392 5867 12393 5893
rect 12365 5866 12393 5867
rect 12261 5109 12289 5110
rect 12261 5083 12262 5109
rect 12262 5083 12288 5109
rect 12288 5083 12289 5109
rect 12261 5082 12289 5083
rect 12313 5109 12341 5110
rect 12313 5083 12314 5109
rect 12314 5083 12340 5109
rect 12340 5083 12341 5109
rect 12313 5082 12341 5083
rect 12365 5109 12393 5110
rect 12365 5083 12366 5109
rect 12366 5083 12392 5109
rect 12392 5083 12393 5109
rect 12365 5082 12393 5083
rect 12261 4325 12289 4326
rect 12261 4299 12262 4325
rect 12262 4299 12288 4325
rect 12288 4299 12289 4325
rect 12261 4298 12289 4299
rect 12313 4325 12341 4326
rect 12313 4299 12314 4325
rect 12314 4299 12340 4325
rect 12340 4299 12341 4325
rect 12313 4298 12341 4299
rect 12365 4325 12393 4326
rect 12365 4299 12366 4325
rect 12366 4299 12392 4325
rect 12392 4299 12393 4325
rect 12365 4298 12393 4299
rect 12261 3541 12289 3542
rect 12261 3515 12262 3541
rect 12262 3515 12288 3541
rect 12288 3515 12289 3541
rect 12261 3514 12289 3515
rect 12313 3541 12341 3542
rect 12313 3515 12314 3541
rect 12314 3515 12340 3541
rect 12340 3515 12341 3541
rect 12313 3514 12341 3515
rect 12365 3541 12393 3542
rect 12365 3515 12366 3541
rect 12366 3515 12392 3541
rect 12392 3515 12393 3541
rect 12365 3514 12393 3515
rect 12261 2757 12289 2758
rect 12261 2731 12262 2757
rect 12262 2731 12288 2757
rect 12288 2731 12289 2757
rect 12261 2730 12289 2731
rect 12313 2757 12341 2758
rect 12313 2731 12314 2757
rect 12314 2731 12340 2757
rect 12340 2731 12341 2757
rect 12313 2730 12341 2731
rect 12365 2757 12393 2758
rect 12365 2731 12366 2757
rect 12366 2731 12392 2757
rect 12392 2731 12393 2757
rect 12365 2730 12393 2731
rect 14592 7853 14620 7854
rect 14592 7827 14593 7853
rect 14593 7827 14619 7853
rect 14619 7827 14620 7853
rect 14592 7826 14620 7827
rect 14644 7853 14672 7854
rect 14644 7827 14645 7853
rect 14645 7827 14671 7853
rect 14671 7827 14672 7853
rect 14644 7826 14672 7827
rect 14696 7853 14724 7854
rect 14696 7827 14697 7853
rect 14697 7827 14723 7853
rect 14723 7827 14724 7853
rect 14696 7826 14724 7827
rect 18606 9758 18634 9786
rect 18830 9561 18858 9562
rect 18830 9535 18831 9561
rect 18831 9535 18857 9561
rect 18857 9535 18858 9561
rect 18830 9534 18858 9535
rect 18550 9198 18578 9226
rect 19110 9758 19138 9786
rect 18942 9505 18970 9506
rect 18942 9479 18943 9505
rect 18943 9479 18969 9505
rect 18969 9479 18970 9505
rect 18942 9478 18970 9479
rect 19110 9478 19138 9506
rect 19254 9421 19282 9422
rect 19254 9395 19255 9421
rect 19255 9395 19281 9421
rect 19281 9395 19282 9421
rect 19254 9394 19282 9395
rect 19306 9421 19334 9422
rect 19306 9395 19307 9421
rect 19307 9395 19333 9421
rect 19333 9395 19334 9421
rect 19306 9394 19334 9395
rect 19358 9421 19386 9422
rect 19358 9395 19359 9421
rect 19359 9395 19385 9421
rect 19385 9395 19386 9421
rect 19358 9394 19386 9395
rect 18886 9142 18914 9170
rect 18830 9086 18858 9114
rect 19110 9086 19138 9114
rect 18998 8918 19026 8946
rect 18606 8862 18634 8890
rect 18270 8777 18298 8778
rect 18270 8751 18271 8777
rect 18271 8751 18297 8777
rect 18297 8751 18298 8777
rect 18270 8750 18298 8751
rect 18942 8806 18970 8834
rect 18886 8694 18914 8722
rect 18774 8441 18802 8442
rect 18774 8415 18775 8441
rect 18775 8415 18801 8441
rect 18801 8415 18802 8441
rect 18774 8414 18802 8415
rect 18942 8358 18970 8386
rect 19110 8777 19138 8778
rect 19110 8751 19111 8777
rect 19111 8751 19137 8777
rect 19137 8751 19138 8777
rect 19110 8750 19138 8751
rect 19254 8637 19282 8638
rect 19254 8611 19255 8637
rect 19255 8611 19281 8637
rect 19281 8611 19282 8637
rect 19254 8610 19282 8611
rect 19306 8637 19334 8638
rect 19306 8611 19307 8637
rect 19307 8611 19333 8637
rect 19333 8611 19334 8637
rect 19306 8610 19334 8611
rect 19358 8637 19386 8638
rect 19358 8611 19359 8637
rect 19359 8611 19385 8637
rect 19385 8611 19386 8637
rect 19358 8610 19386 8611
rect 19166 8105 19194 8106
rect 19166 8079 19167 8105
rect 19167 8079 19193 8105
rect 19193 8079 19194 8105
rect 19166 8078 19194 8079
rect 16923 7461 16951 7462
rect 16923 7435 16924 7461
rect 16924 7435 16950 7461
rect 16950 7435 16951 7461
rect 16923 7434 16951 7435
rect 16975 7461 17003 7462
rect 16975 7435 16976 7461
rect 16976 7435 17002 7461
rect 17002 7435 17003 7461
rect 16975 7434 17003 7435
rect 17027 7461 17055 7462
rect 17027 7435 17028 7461
rect 17028 7435 17054 7461
rect 17054 7435 17055 7461
rect 17027 7434 17055 7435
rect 18830 7406 18858 7434
rect 19254 7853 19282 7854
rect 19254 7827 19255 7853
rect 19255 7827 19281 7853
rect 19281 7827 19282 7853
rect 19254 7826 19282 7827
rect 19306 7853 19334 7854
rect 19306 7827 19307 7853
rect 19307 7827 19333 7853
rect 19333 7827 19334 7853
rect 19306 7826 19334 7827
rect 19358 7853 19386 7854
rect 19358 7827 19359 7853
rect 19359 7827 19385 7853
rect 19385 7827 19386 7853
rect 19358 7826 19386 7827
rect 18998 7742 19026 7770
rect 19110 7406 19138 7434
rect 14592 7069 14620 7070
rect 14592 7043 14593 7069
rect 14593 7043 14619 7069
rect 14619 7043 14620 7069
rect 14592 7042 14620 7043
rect 14644 7069 14672 7070
rect 14644 7043 14645 7069
rect 14645 7043 14671 7069
rect 14671 7043 14672 7069
rect 14644 7042 14672 7043
rect 14696 7069 14724 7070
rect 14696 7043 14697 7069
rect 14697 7043 14723 7069
rect 14723 7043 14724 7069
rect 14696 7042 14724 7043
rect 19254 7069 19282 7070
rect 19254 7043 19255 7069
rect 19255 7043 19281 7069
rect 19281 7043 19282 7069
rect 19254 7042 19282 7043
rect 19306 7069 19334 7070
rect 19306 7043 19307 7069
rect 19307 7043 19333 7069
rect 19333 7043 19334 7069
rect 19306 7042 19334 7043
rect 19358 7069 19386 7070
rect 19358 7043 19359 7069
rect 19359 7043 19385 7069
rect 19385 7043 19386 7069
rect 19358 7042 19386 7043
rect 18998 6958 19026 6986
rect 17654 6817 17682 6818
rect 17654 6791 17655 6817
rect 17655 6791 17681 6817
rect 17681 6791 17682 6817
rect 17654 6790 17682 6791
rect 17878 6790 17906 6818
rect 16923 6677 16951 6678
rect 16923 6651 16924 6677
rect 16924 6651 16950 6677
rect 16950 6651 16951 6677
rect 16923 6650 16951 6651
rect 16975 6677 17003 6678
rect 16975 6651 16976 6677
rect 16976 6651 17002 6677
rect 17002 6651 17003 6677
rect 16975 6650 17003 6651
rect 17027 6677 17055 6678
rect 17027 6651 17028 6677
rect 17028 6651 17054 6677
rect 17054 6651 17055 6677
rect 17027 6650 17055 6651
rect 14592 6285 14620 6286
rect 14592 6259 14593 6285
rect 14593 6259 14619 6285
rect 14619 6259 14620 6285
rect 14592 6258 14620 6259
rect 14644 6285 14672 6286
rect 14644 6259 14645 6285
rect 14645 6259 14671 6285
rect 14671 6259 14672 6285
rect 14644 6258 14672 6259
rect 14696 6285 14724 6286
rect 14696 6259 14697 6285
rect 14697 6259 14723 6285
rect 14723 6259 14724 6285
rect 14696 6258 14724 6259
rect 19254 6285 19282 6286
rect 19254 6259 19255 6285
rect 19255 6259 19281 6285
rect 19281 6259 19282 6285
rect 19254 6258 19282 6259
rect 19306 6285 19334 6286
rect 19306 6259 19307 6285
rect 19307 6259 19333 6285
rect 19333 6259 19334 6285
rect 19306 6258 19334 6259
rect 19358 6285 19386 6286
rect 19358 6259 19359 6285
rect 19359 6259 19385 6285
rect 19385 6259 19386 6285
rect 19358 6258 19386 6259
rect 16923 5893 16951 5894
rect 16923 5867 16924 5893
rect 16924 5867 16950 5893
rect 16950 5867 16951 5893
rect 16923 5866 16951 5867
rect 16975 5893 17003 5894
rect 16975 5867 16976 5893
rect 16976 5867 17002 5893
rect 17002 5867 17003 5893
rect 16975 5866 17003 5867
rect 17027 5893 17055 5894
rect 17027 5867 17028 5893
rect 17028 5867 17054 5893
rect 17054 5867 17055 5893
rect 17027 5866 17055 5867
rect 14592 5501 14620 5502
rect 14592 5475 14593 5501
rect 14593 5475 14619 5501
rect 14619 5475 14620 5501
rect 14592 5474 14620 5475
rect 14644 5501 14672 5502
rect 14644 5475 14645 5501
rect 14645 5475 14671 5501
rect 14671 5475 14672 5501
rect 14644 5474 14672 5475
rect 14696 5501 14724 5502
rect 14696 5475 14697 5501
rect 14697 5475 14723 5501
rect 14723 5475 14724 5501
rect 14696 5474 14724 5475
rect 19254 5501 19282 5502
rect 19254 5475 19255 5501
rect 19255 5475 19281 5501
rect 19281 5475 19282 5501
rect 19254 5474 19282 5475
rect 19306 5501 19334 5502
rect 19306 5475 19307 5501
rect 19307 5475 19333 5501
rect 19333 5475 19334 5501
rect 19306 5474 19334 5475
rect 19358 5501 19386 5502
rect 19358 5475 19359 5501
rect 19359 5475 19385 5501
rect 19385 5475 19386 5501
rect 19358 5474 19386 5475
rect 16923 5109 16951 5110
rect 16923 5083 16924 5109
rect 16924 5083 16950 5109
rect 16950 5083 16951 5109
rect 16923 5082 16951 5083
rect 16975 5109 17003 5110
rect 16975 5083 16976 5109
rect 16976 5083 17002 5109
rect 17002 5083 17003 5109
rect 16975 5082 17003 5083
rect 17027 5109 17055 5110
rect 17027 5083 17028 5109
rect 17028 5083 17054 5109
rect 17054 5083 17055 5109
rect 17027 5082 17055 5083
rect 14592 4717 14620 4718
rect 14592 4691 14593 4717
rect 14593 4691 14619 4717
rect 14619 4691 14620 4717
rect 14592 4690 14620 4691
rect 14644 4717 14672 4718
rect 14644 4691 14645 4717
rect 14645 4691 14671 4717
rect 14671 4691 14672 4717
rect 14644 4690 14672 4691
rect 14696 4717 14724 4718
rect 14696 4691 14697 4717
rect 14697 4691 14723 4717
rect 14723 4691 14724 4717
rect 14696 4690 14724 4691
rect 19254 4717 19282 4718
rect 19254 4691 19255 4717
rect 19255 4691 19281 4717
rect 19281 4691 19282 4717
rect 19254 4690 19282 4691
rect 19306 4717 19334 4718
rect 19306 4691 19307 4717
rect 19307 4691 19333 4717
rect 19333 4691 19334 4717
rect 19306 4690 19334 4691
rect 19358 4717 19386 4718
rect 19358 4691 19359 4717
rect 19359 4691 19385 4717
rect 19385 4691 19386 4717
rect 19358 4690 19386 4691
rect 16923 4325 16951 4326
rect 16923 4299 16924 4325
rect 16924 4299 16950 4325
rect 16950 4299 16951 4325
rect 16923 4298 16951 4299
rect 16975 4325 17003 4326
rect 16975 4299 16976 4325
rect 16976 4299 17002 4325
rect 17002 4299 17003 4325
rect 16975 4298 17003 4299
rect 17027 4325 17055 4326
rect 17027 4299 17028 4325
rect 17028 4299 17054 4325
rect 17054 4299 17055 4325
rect 17027 4298 17055 4299
rect 14592 3933 14620 3934
rect 14592 3907 14593 3933
rect 14593 3907 14619 3933
rect 14619 3907 14620 3933
rect 14592 3906 14620 3907
rect 14644 3933 14672 3934
rect 14644 3907 14645 3933
rect 14645 3907 14671 3933
rect 14671 3907 14672 3933
rect 14644 3906 14672 3907
rect 14696 3933 14724 3934
rect 14696 3907 14697 3933
rect 14697 3907 14723 3933
rect 14723 3907 14724 3933
rect 14696 3906 14724 3907
rect 19254 3933 19282 3934
rect 19254 3907 19255 3933
rect 19255 3907 19281 3933
rect 19281 3907 19282 3933
rect 19254 3906 19282 3907
rect 19306 3933 19334 3934
rect 19306 3907 19307 3933
rect 19307 3907 19333 3933
rect 19333 3907 19334 3933
rect 19306 3906 19334 3907
rect 19358 3933 19386 3934
rect 19358 3907 19359 3933
rect 19359 3907 19385 3933
rect 19385 3907 19386 3933
rect 19358 3906 19386 3907
rect 16923 3541 16951 3542
rect 16923 3515 16924 3541
rect 16924 3515 16950 3541
rect 16950 3515 16951 3541
rect 16923 3514 16951 3515
rect 16975 3541 17003 3542
rect 16975 3515 16976 3541
rect 16976 3515 17002 3541
rect 17002 3515 17003 3541
rect 16975 3514 17003 3515
rect 17027 3541 17055 3542
rect 17027 3515 17028 3541
rect 17028 3515 17054 3541
rect 17054 3515 17055 3541
rect 17027 3514 17055 3515
rect 14592 3149 14620 3150
rect 14592 3123 14593 3149
rect 14593 3123 14619 3149
rect 14619 3123 14620 3149
rect 14592 3122 14620 3123
rect 14644 3149 14672 3150
rect 14644 3123 14645 3149
rect 14645 3123 14671 3149
rect 14671 3123 14672 3149
rect 14644 3122 14672 3123
rect 14696 3149 14724 3150
rect 14696 3123 14697 3149
rect 14697 3123 14723 3149
rect 14723 3123 14724 3149
rect 14696 3122 14724 3123
rect 19254 3149 19282 3150
rect 19254 3123 19255 3149
rect 19255 3123 19281 3149
rect 19281 3123 19282 3149
rect 19254 3122 19282 3123
rect 19306 3149 19334 3150
rect 19306 3123 19307 3149
rect 19307 3123 19333 3149
rect 19333 3123 19334 3149
rect 19306 3122 19334 3123
rect 19358 3149 19386 3150
rect 19358 3123 19359 3149
rect 19359 3123 19385 3149
rect 19385 3123 19386 3149
rect 19358 3122 19386 3123
rect 16923 2757 16951 2758
rect 16923 2731 16924 2757
rect 16924 2731 16950 2757
rect 16950 2731 16951 2757
rect 16923 2730 16951 2731
rect 16975 2757 17003 2758
rect 16975 2731 16976 2757
rect 16976 2731 17002 2757
rect 17002 2731 17003 2757
rect 16975 2730 17003 2731
rect 17027 2757 17055 2758
rect 17027 2731 17028 2757
rect 17028 2731 17054 2757
rect 17054 2731 17055 2757
rect 17027 2730 17055 2731
rect 14592 2365 14620 2366
rect 14592 2339 14593 2365
rect 14593 2339 14619 2365
rect 14619 2339 14620 2365
rect 14592 2338 14620 2339
rect 14644 2365 14672 2366
rect 14644 2339 14645 2365
rect 14645 2339 14671 2365
rect 14671 2339 14672 2365
rect 14644 2338 14672 2339
rect 14696 2365 14724 2366
rect 14696 2339 14697 2365
rect 14697 2339 14723 2365
rect 14723 2339 14724 2365
rect 14696 2338 14724 2339
rect 19254 2365 19282 2366
rect 19254 2339 19255 2365
rect 19255 2339 19281 2365
rect 19281 2339 19282 2365
rect 19254 2338 19282 2339
rect 19306 2365 19334 2366
rect 19306 2339 19307 2365
rect 19307 2339 19333 2365
rect 19333 2339 19334 2365
rect 19306 2338 19334 2339
rect 19358 2365 19386 2366
rect 19358 2339 19359 2365
rect 19359 2339 19385 2365
rect 19385 2339 19386 2365
rect 19358 2338 19386 2339
rect 13118 2057 13146 2058
rect 13118 2031 13119 2057
rect 13119 2031 13145 2057
rect 13145 2031 13146 2057
rect 13118 2030 13146 2031
rect 12261 1973 12289 1974
rect 12261 1947 12262 1973
rect 12262 1947 12288 1973
rect 12288 1947 12289 1973
rect 12261 1946 12289 1947
rect 12313 1973 12341 1974
rect 12313 1947 12314 1973
rect 12314 1947 12340 1973
rect 12340 1947 12341 1973
rect 12313 1946 12341 1947
rect 12365 1973 12393 1974
rect 12365 1947 12366 1973
rect 12366 1947 12392 1973
rect 12392 1947 12393 1973
rect 12365 1946 12393 1947
rect 16923 1973 16951 1974
rect 16923 1947 16924 1973
rect 16924 1947 16950 1973
rect 16950 1947 16951 1973
rect 16923 1946 16951 1947
rect 16975 1973 17003 1974
rect 16975 1947 16976 1973
rect 16976 1947 17002 1973
rect 17002 1947 17003 1973
rect 16975 1946 17003 1947
rect 17027 1973 17055 1974
rect 17027 1947 17028 1973
rect 17028 1947 17054 1973
rect 17054 1947 17055 1973
rect 17027 1946 17055 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
rect 14592 1581 14620 1582
rect 14592 1555 14593 1581
rect 14593 1555 14619 1581
rect 14619 1555 14620 1581
rect 14592 1554 14620 1555
rect 14644 1581 14672 1582
rect 14644 1555 14645 1581
rect 14645 1555 14671 1581
rect 14671 1555 14672 1581
rect 14644 1554 14672 1555
rect 14696 1581 14724 1582
rect 14696 1555 14697 1581
rect 14697 1555 14723 1581
rect 14723 1555 14724 1581
rect 14696 1554 14724 1555
rect 19254 1581 19282 1582
rect 19254 1555 19255 1581
rect 19255 1555 19281 1581
rect 19281 1555 19282 1581
rect 19254 1554 19282 1555
rect 19306 1581 19334 1582
rect 19306 1555 19307 1581
rect 19307 1555 19333 1581
rect 19333 1555 19334 1581
rect 19306 1554 19334 1555
rect 19358 1581 19386 1582
rect 19358 1555 19359 1581
rect 19359 1555 19385 1581
rect 19385 1555 19386 1581
rect 19358 1554 19386 1555
<< metal3 >>
rect 2932 18410 2937 18438
rect 2965 18410 2989 18438
rect 3017 18410 3041 18438
rect 3069 18410 3074 18438
rect 7594 18410 7599 18438
rect 7627 18410 7651 18438
rect 7679 18410 7703 18438
rect 7731 18410 7736 18438
rect 12256 18410 12261 18438
rect 12289 18410 12313 18438
rect 12341 18410 12365 18438
rect 12393 18410 12398 18438
rect 16918 18410 16923 18438
rect 16951 18410 16975 18438
rect 17003 18410 17027 18438
rect 17055 18410 17060 18438
rect 8409 18326 8414 18354
rect 8442 18326 9030 18354
rect 9058 18326 9063 18354
rect 5263 18018 5268 18046
rect 5296 18018 5320 18046
rect 5348 18018 5372 18046
rect 5400 18018 5405 18046
rect 9925 18018 9930 18046
rect 9958 18018 9982 18046
rect 10010 18018 10034 18046
rect 10062 18018 10067 18046
rect 14587 18018 14592 18046
rect 14620 18018 14644 18046
rect 14672 18018 14696 18046
rect 14724 18018 14729 18046
rect 19249 18018 19254 18046
rect 19282 18018 19306 18046
rect 19334 18018 19358 18046
rect 19386 18018 19391 18046
rect 7513 17934 7518 17962
rect 7546 17934 7854 17962
rect 7882 17934 7887 17962
rect 9473 17934 9478 17962
rect 9506 17934 9870 17962
rect 9898 17934 9903 17962
rect 2932 17626 2937 17654
rect 2965 17626 2989 17654
rect 3017 17626 3041 17654
rect 3069 17626 3074 17654
rect 7594 17626 7599 17654
rect 7627 17626 7651 17654
rect 7679 17626 7703 17654
rect 7731 17626 7736 17654
rect 12256 17626 12261 17654
rect 12289 17626 12313 17654
rect 12341 17626 12365 17654
rect 12393 17626 12398 17654
rect 16918 17626 16923 17654
rect 16951 17626 16975 17654
rect 17003 17626 17027 17654
rect 17055 17626 17060 17654
rect 5263 17234 5268 17262
rect 5296 17234 5320 17262
rect 5348 17234 5372 17262
rect 5400 17234 5405 17262
rect 9925 17234 9930 17262
rect 9958 17234 9982 17262
rect 10010 17234 10034 17262
rect 10062 17234 10067 17262
rect 14587 17234 14592 17262
rect 14620 17234 14644 17262
rect 14672 17234 14696 17262
rect 14724 17234 14729 17262
rect 19249 17234 19254 17262
rect 19282 17234 19306 17262
rect 19334 17234 19358 17262
rect 19386 17234 19391 17262
rect 2932 16842 2937 16870
rect 2965 16842 2989 16870
rect 3017 16842 3041 16870
rect 3069 16842 3074 16870
rect 7594 16842 7599 16870
rect 7627 16842 7651 16870
rect 7679 16842 7703 16870
rect 7731 16842 7736 16870
rect 12256 16842 12261 16870
rect 12289 16842 12313 16870
rect 12341 16842 12365 16870
rect 12393 16842 12398 16870
rect 16918 16842 16923 16870
rect 16951 16842 16975 16870
rect 17003 16842 17027 16870
rect 17055 16842 17060 16870
rect 5263 16450 5268 16478
rect 5296 16450 5320 16478
rect 5348 16450 5372 16478
rect 5400 16450 5405 16478
rect 9925 16450 9930 16478
rect 9958 16450 9982 16478
rect 10010 16450 10034 16478
rect 10062 16450 10067 16478
rect 14587 16450 14592 16478
rect 14620 16450 14644 16478
rect 14672 16450 14696 16478
rect 14724 16450 14729 16478
rect 19249 16450 19254 16478
rect 19282 16450 19306 16478
rect 19334 16450 19358 16478
rect 19386 16450 19391 16478
rect 2932 16058 2937 16086
rect 2965 16058 2989 16086
rect 3017 16058 3041 16086
rect 3069 16058 3074 16086
rect 7594 16058 7599 16086
rect 7627 16058 7651 16086
rect 7679 16058 7703 16086
rect 7731 16058 7736 16086
rect 12256 16058 12261 16086
rect 12289 16058 12313 16086
rect 12341 16058 12365 16086
rect 12393 16058 12398 16086
rect 16918 16058 16923 16086
rect 16951 16058 16975 16086
rect 17003 16058 17027 16086
rect 17055 16058 17060 16086
rect 5263 15666 5268 15694
rect 5296 15666 5320 15694
rect 5348 15666 5372 15694
rect 5400 15666 5405 15694
rect 9925 15666 9930 15694
rect 9958 15666 9982 15694
rect 10010 15666 10034 15694
rect 10062 15666 10067 15694
rect 14587 15666 14592 15694
rect 14620 15666 14644 15694
rect 14672 15666 14696 15694
rect 14724 15666 14729 15694
rect 19249 15666 19254 15694
rect 19282 15666 19306 15694
rect 19334 15666 19358 15694
rect 19386 15666 19391 15694
rect 2932 15274 2937 15302
rect 2965 15274 2989 15302
rect 3017 15274 3041 15302
rect 3069 15274 3074 15302
rect 7594 15274 7599 15302
rect 7627 15274 7651 15302
rect 7679 15274 7703 15302
rect 7731 15274 7736 15302
rect 12256 15274 12261 15302
rect 12289 15274 12313 15302
rect 12341 15274 12365 15302
rect 12393 15274 12398 15302
rect 16918 15274 16923 15302
rect 16951 15274 16975 15302
rect 17003 15274 17027 15302
rect 17055 15274 17060 15302
rect 8297 15078 8302 15106
rect 8330 15078 8694 15106
rect 8722 15078 8727 15106
rect 8017 14966 8022 14994
rect 8050 14966 8414 14994
rect 8442 14966 8447 14994
rect 5263 14882 5268 14910
rect 5296 14882 5320 14910
rect 5348 14882 5372 14910
rect 5400 14882 5405 14910
rect 9925 14882 9930 14910
rect 9958 14882 9982 14910
rect 10010 14882 10034 14910
rect 10062 14882 10067 14910
rect 14587 14882 14592 14910
rect 14620 14882 14644 14910
rect 14672 14882 14696 14910
rect 14724 14882 14729 14910
rect 19249 14882 19254 14910
rect 19282 14882 19306 14910
rect 19334 14882 19358 14910
rect 19386 14882 19391 14910
rect 10369 14686 10374 14714
rect 10402 14686 10598 14714
rect 10626 14686 10631 14714
rect 2932 14490 2937 14518
rect 2965 14490 2989 14518
rect 3017 14490 3041 14518
rect 3069 14490 3074 14518
rect 7594 14490 7599 14518
rect 7627 14490 7651 14518
rect 7679 14490 7703 14518
rect 7731 14490 7736 14518
rect 12256 14490 12261 14518
rect 12289 14490 12313 14518
rect 12341 14490 12365 14518
rect 12393 14490 12398 14518
rect 16918 14490 16923 14518
rect 16951 14490 16975 14518
rect 17003 14490 17027 14518
rect 17055 14490 17060 14518
rect 5263 14098 5268 14126
rect 5296 14098 5320 14126
rect 5348 14098 5372 14126
rect 5400 14098 5405 14126
rect 9925 14098 9930 14126
rect 9958 14098 9982 14126
rect 10010 14098 10034 14126
rect 10062 14098 10067 14126
rect 14587 14098 14592 14126
rect 14620 14098 14644 14126
rect 14672 14098 14696 14126
rect 14724 14098 14729 14126
rect 19249 14098 19254 14126
rect 19282 14098 19306 14126
rect 19334 14098 19358 14126
rect 19386 14098 19391 14126
rect 2932 13706 2937 13734
rect 2965 13706 2989 13734
rect 3017 13706 3041 13734
rect 3069 13706 3074 13734
rect 7594 13706 7599 13734
rect 7627 13706 7651 13734
rect 7679 13706 7703 13734
rect 7731 13706 7736 13734
rect 12256 13706 12261 13734
rect 12289 13706 12313 13734
rect 12341 13706 12365 13734
rect 12393 13706 12398 13734
rect 16918 13706 16923 13734
rect 16951 13706 16975 13734
rect 17003 13706 17027 13734
rect 17055 13706 17060 13734
rect 5263 13314 5268 13342
rect 5296 13314 5320 13342
rect 5348 13314 5372 13342
rect 5400 13314 5405 13342
rect 9925 13314 9930 13342
rect 9958 13314 9982 13342
rect 10010 13314 10034 13342
rect 10062 13314 10067 13342
rect 14587 13314 14592 13342
rect 14620 13314 14644 13342
rect 14672 13314 14696 13342
rect 14724 13314 14729 13342
rect 19249 13314 19254 13342
rect 19282 13314 19306 13342
rect 19334 13314 19358 13342
rect 19386 13314 19391 13342
rect 2932 12922 2937 12950
rect 2965 12922 2989 12950
rect 3017 12922 3041 12950
rect 3069 12922 3074 12950
rect 7594 12922 7599 12950
rect 7627 12922 7651 12950
rect 7679 12922 7703 12950
rect 7731 12922 7736 12950
rect 12256 12922 12261 12950
rect 12289 12922 12313 12950
rect 12341 12922 12365 12950
rect 12393 12922 12398 12950
rect 16918 12922 16923 12950
rect 16951 12922 16975 12950
rect 17003 12922 17027 12950
rect 17055 12922 17060 12950
rect 0 12810 400 12824
rect 0 12782 966 12810
rect 994 12782 999 12810
rect 0 12768 400 12782
rect 5263 12530 5268 12558
rect 5296 12530 5320 12558
rect 5348 12530 5372 12558
rect 5400 12530 5405 12558
rect 9925 12530 9930 12558
rect 9958 12530 9982 12558
rect 10010 12530 10034 12558
rect 10062 12530 10067 12558
rect 14587 12530 14592 12558
rect 14620 12530 14644 12558
rect 14672 12530 14696 12558
rect 14724 12530 14729 12558
rect 19249 12530 19254 12558
rect 19282 12530 19306 12558
rect 19334 12530 19358 12558
rect 19386 12530 19391 12558
rect 0 12474 400 12488
rect 0 12446 854 12474
rect 882 12446 1246 12474
rect 1274 12446 1279 12474
rect 0 12432 400 12446
rect 1017 12390 1022 12418
rect 1050 12390 8022 12418
rect 8050 12390 8055 12418
rect 11209 12334 11214 12362
rect 11242 12334 17822 12362
rect 17850 12334 17855 12362
rect 0 12138 400 12152
rect 2932 12138 2937 12166
rect 2965 12138 2989 12166
rect 3017 12138 3041 12166
rect 3069 12138 3074 12166
rect 7594 12138 7599 12166
rect 7627 12138 7651 12166
rect 7679 12138 7703 12166
rect 7731 12138 7736 12166
rect 12256 12138 12261 12166
rect 12289 12138 12313 12166
rect 12341 12138 12365 12166
rect 12393 12138 12398 12166
rect 16918 12138 16923 12166
rect 16951 12138 16975 12166
rect 17003 12138 17027 12166
rect 17055 12138 17060 12166
rect 19600 12138 20000 12152
rect 0 12110 854 12138
rect 882 12110 1246 12138
rect 1274 12110 1279 12138
rect 18993 12110 18998 12138
rect 19026 12110 20000 12138
rect 0 12096 400 12110
rect 19600 12096 20000 12110
rect 1017 11830 1022 11858
rect 1050 11830 8022 11858
rect 8050 11830 8055 11858
rect 8521 11830 8526 11858
rect 8554 11830 8806 11858
rect 8834 11830 8839 11858
rect 18825 11830 18830 11858
rect 18858 11830 19110 11858
rect 19138 11830 19474 11858
rect 0 11802 400 11816
rect 19446 11802 19474 11830
rect 19600 11802 20000 11816
rect 0 11774 854 11802
rect 882 11774 1246 11802
rect 1274 11774 1279 11802
rect 19446 11774 20000 11802
rect 0 11760 400 11774
rect 5263 11746 5268 11774
rect 5296 11746 5320 11774
rect 5348 11746 5372 11774
rect 5400 11746 5405 11774
rect 9925 11746 9930 11774
rect 9958 11746 9982 11774
rect 10010 11746 10034 11774
rect 10062 11746 10067 11774
rect 14587 11746 14592 11774
rect 14620 11746 14644 11774
rect 14672 11746 14696 11774
rect 14724 11746 14729 11774
rect 19249 11746 19254 11774
rect 19282 11746 19306 11774
rect 19334 11746 19358 11774
rect 19386 11746 19391 11774
rect 19600 11760 20000 11774
rect 12049 11606 12054 11634
rect 12082 11606 18942 11634
rect 18970 11606 18975 11634
rect 0 11466 400 11480
rect 19600 11466 20000 11480
rect 0 11438 854 11466
rect 882 11438 1246 11466
rect 1274 11438 1279 11466
rect 18825 11438 18830 11466
rect 18858 11438 19110 11466
rect 19138 11438 20000 11466
rect 0 11424 400 11438
rect 19600 11424 20000 11438
rect 2932 11354 2937 11382
rect 2965 11354 2989 11382
rect 3017 11354 3041 11382
rect 3069 11354 3074 11382
rect 7594 11354 7599 11382
rect 7627 11354 7651 11382
rect 7679 11354 7703 11382
rect 7731 11354 7736 11382
rect 12256 11354 12261 11382
rect 12289 11354 12313 11382
rect 12341 11354 12365 11382
rect 12393 11354 12398 11382
rect 16918 11354 16923 11382
rect 16951 11354 16975 11382
rect 17003 11354 17027 11382
rect 17055 11354 17060 11382
rect 1017 11158 1022 11186
rect 1050 11158 7854 11186
rect 7882 11158 7887 11186
rect 0 11130 400 11144
rect 19600 11130 20000 11144
rect 0 11102 854 11130
rect 882 11102 1246 11130
rect 1274 11102 1279 11130
rect 18825 11102 18830 11130
rect 18858 11102 19110 11130
rect 19138 11102 20000 11130
rect 0 11088 400 11102
rect 19600 11088 20000 11102
rect 1353 11046 1358 11074
rect 1386 11046 8862 11074
rect 8890 11046 8895 11074
rect 10873 11046 10878 11074
rect 10906 11046 17822 11074
rect 17850 11046 17855 11074
rect 5263 10962 5268 10990
rect 5296 10962 5320 10990
rect 5348 10962 5372 10990
rect 5400 10962 5405 10990
rect 9925 10962 9930 10990
rect 9958 10962 9982 10990
rect 10010 10962 10034 10990
rect 10062 10962 10067 10990
rect 14587 10962 14592 10990
rect 14620 10962 14644 10990
rect 14672 10962 14696 10990
rect 14724 10962 14729 10990
rect 19249 10962 19254 10990
rect 19282 10962 19306 10990
rect 19334 10962 19358 10990
rect 19386 10962 19391 10990
rect 10705 10878 10710 10906
rect 10738 10878 11214 10906
rect 11242 10878 11247 10906
rect 15946 10878 18942 10906
rect 18970 10878 18975 10906
rect 1017 10822 1022 10850
rect 1050 10822 8246 10850
rect 8274 10822 8279 10850
rect 0 10794 400 10808
rect 15946 10794 15974 10878
rect 19600 10794 20000 10808
rect 0 10766 1190 10794
rect 1218 10766 1582 10794
rect 1610 10766 1615 10794
rect 10929 10766 10934 10794
rect 10962 10766 11158 10794
rect 11186 10766 11191 10794
rect 11601 10766 11606 10794
rect 11634 10766 15974 10794
rect 18993 10766 18998 10794
rect 19026 10766 20000 10794
rect 0 10752 400 10766
rect 19600 10752 20000 10766
rect 849 10710 854 10738
rect 882 10710 1470 10738
rect 1498 10710 1503 10738
rect 2932 10570 2937 10598
rect 2965 10570 2989 10598
rect 3017 10570 3041 10598
rect 3069 10570 3074 10598
rect 7594 10570 7599 10598
rect 7627 10570 7651 10598
rect 7679 10570 7703 10598
rect 7731 10570 7736 10598
rect 12256 10570 12261 10598
rect 12289 10570 12313 10598
rect 12341 10570 12365 10598
rect 12393 10570 12398 10598
rect 16918 10570 16923 10598
rect 16951 10570 16975 10598
rect 17003 10570 17027 10598
rect 17055 10570 17060 10598
rect 0 10458 400 10472
rect 19600 10458 20000 10472
rect 0 10430 854 10458
rect 882 10430 887 10458
rect 18265 10430 18270 10458
rect 18298 10430 19110 10458
rect 19138 10430 20000 10458
rect 0 10416 400 10430
rect 19600 10416 20000 10430
rect 11713 10374 11718 10402
rect 11746 10374 18886 10402
rect 18914 10374 18919 10402
rect 1073 10318 1078 10346
rect 1106 10318 7742 10346
rect 7770 10318 9422 10346
rect 9450 10318 9455 10346
rect 12217 10318 12222 10346
rect 12250 10318 18942 10346
rect 18970 10318 18975 10346
rect 1017 10262 1022 10290
rect 1050 10262 8862 10290
rect 8890 10262 8895 10290
rect 5263 10178 5268 10206
rect 5296 10178 5320 10206
rect 5348 10178 5372 10206
rect 5400 10178 5405 10206
rect 9925 10178 9930 10206
rect 9958 10178 9982 10206
rect 10010 10178 10034 10206
rect 10062 10178 10067 10206
rect 14587 10178 14592 10206
rect 14620 10178 14644 10206
rect 14672 10178 14696 10206
rect 14724 10178 14729 10206
rect 19249 10178 19254 10206
rect 19282 10178 19306 10206
rect 19334 10178 19358 10206
rect 19386 10178 19391 10206
rect 0 10122 400 10136
rect 19600 10122 20000 10136
rect 0 10094 854 10122
rect 882 10094 1246 10122
rect 1274 10094 1279 10122
rect 18825 10094 18830 10122
rect 18858 10094 20000 10122
rect 0 10080 400 10094
rect 19600 10080 20000 10094
rect 2417 10038 2422 10066
rect 2450 10038 8246 10066
rect 8274 10038 8279 10066
rect 8689 10038 8694 10066
rect 8722 10038 8727 10066
rect 8694 10010 8722 10038
rect 2137 9982 2142 10010
rect 2170 9982 8722 10010
rect 961 9870 966 9898
rect 994 9870 999 9898
rect 0 9786 400 9800
rect 966 9786 994 9870
rect 2932 9786 2937 9814
rect 2965 9786 2989 9814
rect 3017 9786 3041 9814
rect 3069 9786 3074 9814
rect 7594 9786 7599 9814
rect 7627 9786 7651 9814
rect 7679 9786 7703 9814
rect 7731 9786 7736 9814
rect 12256 9786 12261 9814
rect 12289 9786 12313 9814
rect 12341 9786 12365 9814
rect 12393 9786 12398 9814
rect 16918 9786 16923 9814
rect 16951 9786 16975 9814
rect 17003 9786 17027 9814
rect 17055 9786 17060 9814
rect 19600 9786 20000 9800
rect 0 9758 994 9786
rect 18601 9758 18606 9786
rect 18634 9758 19110 9786
rect 19138 9758 20000 9786
rect 0 9744 400 9758
rect 19600 9744 20000 9758
rect 9921 9646 9926 9674
rect 9954 9646 10822 9674
rect 10850 9646 10855 9674
rect 8241 9590 8246 9618
rect 8274 9590 8279 9618
rect 1129 9534 1134 9562
rect 1162 9534 7742 9562
rect 7770 9534 7775 9562
rect 8246 9506 8274 9590
rect 8353 9534 8358 9562
rect 8386 9534 8806 9562
rect 8834 9534 8839 9562
rect 18825 9534 18830 9562
rect 18858 9534 19138 9562
rect 19110 9506 19138 9534
rect 1017 9478 1022 9506
rect 1050 9478 8274 9506
rect 9305 9478 9310 9506
rect 9338 9478 10094 9506
rect 10122 9478 10127 9506
rect 10257 9478 10262 9506
rect 10290 9478 11270 9506
rect 11298 9478 11303 9506
rect 12161 9478 12166 9506
rect 12194 9478 18942 9506
rect 18970 9478 18975 9506
rect 19105 9478 19110 9506
rect 19138 9478 19474 9506
rect 0 9450 400 9464
rect 19446 9450 19474 9478
rect 19600 9450 20000 9464
rect 0 9422 854 9450
rect 882 9422 1246 9450
rect 1274 9422 1279 9450
rect 19446 9422 20000 9450
rect 0 9408 400 9422
rect 5263 9394 5268 9422
rect 5296 9394 5320 9422
rect 5348 9394 5372 9422
rect 5400 9394 5405 9422
rect 9925 9394 9930 9422
rect 9958 9394 9982 9422
rect 10010 9394 10034 9422
rect 10062 9394 10067 9422
rect 14587 9394 14592 9422
rect 14620 9394 14644 9422
rect 14672 9394 14696 9422
rect 14724 9394 14729 9422
rect 19249 9394 19254 9422
rect 19282 9394 19306 9422
rect 19334 9394 19358 9422
rect 19386 9394 19391 9422
rect 19600 9408 20000 9422
rect 11657 9310 11662 9338
rect 11690 9310 17822 9338
rect 17850 9310 17855 9338
rect 9193 9254 9198 9282
rect 9226 9254 9646 9282
rect 9674 9254 9679 9282
rect 1017 9198 1022 9226
rect 1050 9198 4214 9226
rect 8017 9198 8022 9226
rect 8050 9198 8694 9226
rect 8722 9198 8727 9226
rect 9361 9198 9366 9226
rect 9394 9198 9399 9226
rect 11713 9198 11718 9226
rect 11746 9198 18550 9226
rect 18578 9198 18583 9226
rect 4186 9170 4214 9198
rect 9366 9170 9394 9198
rect 4186 9142 9394 9170
rect 10593 9142 10598 9170
rect 10626 9142 12670 9170
rect 12698 9142 18886 9170
rect 18914 9142 18919 9170
rect 0 9114 400 9128
rect 19600 9114 20000 9128
rect 0 9086 854 9114
rect 882 9086 1246 9114
rect 1274 9086 1279 9114
rect 18825 9086 18830 9114
rect 18858 9086 19110 9114
rect 19138 9086 20000 9114
rect 0 9072 400 9086
rect 19600 9072 20000 9086
rect 2932 9002 2937 9030
rect 2965 9002 2989 9030
rect 3017 9002 3041 9030
rect 3069 9002 3074 9030
rect 7594 9002 7599 9030
rect 7627 9002 7651 9030
rect 7679 9002 7703 9030
rect 7731 9002 7736 9030
rect 12256 9002 12261 9030
rect 12289 9002 12313 9030
rect 12341 9002 12365 9030
rect 12393 9002 12398 9030
rect 16918 9002 16923 9030
rect 16951 9002 16975 9030
rect 17003 9002 17027 9030
rect 17055 9002 17060 9030
rect 11041 8918 11046 8946
rect 11074 8918 12950 8946
rect 12978 8918 18998 8946
rect 19026 8918 19031 8946
rect 12217 8862 12222 8890
rect 12250 8862 18606 8890
rect 18634 8862 18639 8890
rect 11713 8806 11718 8834
rect 11746 8806 18942 8834
rect 18970 8806 18975 8834
rect 0 8778 400 8792
rect 19600 8778 20000 8792
rect 0 8750 854 8778
rect 882 8750 1246 8778
rect 1274 8750 1279 8778
rect 10649 8750 10654 8778
rect 10682 8750 15974 8778
rect 18265 8750 18270 8778
rect 18298 8750 19110 8778
rect 19138 8750 20000 8778
rect 0 8736 400 8750
rect 15946 8722 15974 8750
rect 19600 8736 20000 8750
rect 15946 8694 18886 8722
rect 18914 8694 18919 8722
rect 5263 8610 5268 8638
rect 5296 8610 5320 8638
rect 5348 8610 5372 8638
rect 5400 8610 5405 8638
rect 9925 8610 9930 8638
rect 9958 8610 9982 8638
rect 10010 8610 10034 8638
rect 10062 8610 10067 8638
rect 14587 8610 14592 8638
rect 14620 8610 14644 8638
rect 14672 8610 14696 8638
rect 14724 8610 14729 8638
rect 19249 8610 19254 8638
rect 19282 8610 19306 8638
rect 19334 8610 19358 8638
rect 19386 8610 19391 8638
rect 0 8442 400 8456
rect 19600 8442 20000 8456
rect 0 8414 966 8442
rect 994 8414 999 8442
rect 18769 8414 18774 8442
rect 18802 8414 20000 8442
rect 0 8400 400 8414
rect 19600 8400 20000 8414
rect 1185 8358 1190 8386
rect 1218 8358 1582 8386
rect 1610 8358 1615 8386
rect 11097 8358 11102 8386
rect 11130 8358 18942 8386
rect 18970 8358 18975 8386
rect 1017 8302 1022 8330
rect 1050 8302 8638 8330
rect 8666 8302 8671 8330
rect 2932 8218 2937 8246
rect 2965 8218 2989 8246
rect 3017 8218 3041 8246
rect 3069 8218 3074 8246
rect 7594 8218 7599 8246
rect 7627 8218 7651 8246
rect 7679 8218 7703 8246
rect 7731 8218 7736 8246
rect 12256 8218 12261 8246
rect 12289 8218 12313 8246
rect 12341 8218 12365 8246
rect 12393 8218 12398 8246
rect 16918 8218 16923 8246
rect 16951 8218 16975 8246
rect 17003 8218 17027 8246
rect 17055 8218 17060 8246
rect 2137 8134 2142 8162
rect 2170 8134 7966 8162
rect 7994 8134 7999 8162
rect 0 8106 400 8120
rect 19600 8106 20000 8120
rect 0 8078 1190 8106
rect 1218 8078 1223 8106
rect 19161 8078 19166 8106
rect 19194 8078 20000 8106
rect 0 8064 400 8078
rect 19600 8064 20000 8078
rect 1353 8022 1358 8050
rect 1386 8022 7966 8050
rect 7994 8022 7999 8050
rect 4186 7966 7574 7994
rect 7602 7966 7607 7994
rect 7681 7966 7686 7994
rect 7714 7966 8302 7994
rect 8330 7966 9478 7994
rect 9506 7966 9511 7994
rect 4186 7938 4214 7966
rect 1017 7910 1022 7938
rect 1050 7910 4214 7938
rect 9249 7910 9254 7938
rect 9282 7910 10038 7938
rect 10066 7910 10071 7938
rect 10201 7910 10206 7938
rect 10234 7910 12614 7938
rect 12642 7910 12647 7938
rect 5263 7826 5268 7854
rect 5296 7826 5320 7854
rect 5348 7826 5372 7854
rect 5400 7826 5405 7854
rect 9925 7826 9930 7854
rect 9958 7826 9982 7854
rect 10010 7826 10034 7854
rect 10062 7826 10067 7854
rect 14587 7826 14592 7854
rect 14620 7826 14644 7854
rect 14672 7826 14696 7854
rect 14724 7826 14729 7854
rect 19249 7826 19254 7854
rect 19282 7826 19306 7854
rect 19334 7826 19358 7854
rect 19386 7826 19391 7854
rect 0 7770 400 7784
rect 19600 7770 20000 7784
rect 0 7742 910 7770
rect 938 7742 943 7770
rect 9865 7742 9870 7770
rect 9898 7742 12166 7770
rect 12194 7742 12199 7770
rect 18993 7742 18998 7770
rect 19026 7742 20000 7770
rect 0 7728 400 7742
rect 19600 7728 20000 7742
rect 7737 7686 7742 7714
rect 7770 7686 8246 7714
rect 8274 7686 8862 7714
rect 8890 7686 9310 7714
rect 9338 7686 9343 7714
rect 9473 7630 9478 7658
rect 9506 7630 9870 7658
rect 9898 7630 9903 7658
rect 2932 7434 2937 7462
rect 2965 7434 2989 7462
rect 3017 7434 3041 7462
rect 3069 7434 3074 7462
rect 7594 7434 7599 7462
rect 7627 7434 7651 7462
rect 7679 7434 7703 7462
rect 7731 7434 7736 7462
rect 12256 7434 12261 7462
rect 12289 7434 12313 7462
rect 12341 7434 12365 7462
rect 12393 7434 12398 7462
rect 16918 7434 16923 7462
rect 16951 7434 16975 7462
rect 17003 7434 17027 7462
rect 17055 7434 17060 7462
rect 19600 7434 20000 7448
rect 18825 7406 18830 7434
rect 18858 7406 19110 7434
rect 19138 7406 20000 7434
rect 19600 7392 20000 7406
rect 7345 7182 7350 7210
rect 7378 7182 8750 7210
rect 8778 7182 8783 7210
rect 19600 7098 20000 7112
rect 19446 7070 20000 7098
rect 5263 7042 5268 7070
rect 5296 7042 5320 7070
rect 5348 7042 5372 7070
rect 5400 7042 5405 7070
rect 9925 7042 9930 7070
rect 9958 7042 9982 7070
rect 10010 7042 10034 7070
rect 10062 7042 10067 7070
rect 14587 7042 14592 7070
rect 14620 7042 14644 7070
rect 14672 7042 14696 7070
rect 14724 7042 14729 7070
rect 19249 7042 19254 7070
rect 19282 7042 19306 7070
rect 19334 7042 19358 7070
rect 19386 7042 19391 7070
rect 19446 6986 19474 7070
rect 19600 7056 20000 7070
rect 18993 6958 18998 6986
rect 19026 6958 19474 6986
rect 11545 6790 11550 6818
rect 11578 6790 17654 6818
rect 17682 6790 17878 6818
rect 17906 6790 17911 6818
rect 2932 6650 2937 6678
rect 2965 6650 2989 6678
rect 3017 6650 3041 6678
rect 3069 6650 3074 6678
rect 7594 6650 7599 6678
rect 7627 6650 7651 6678
rect 7679 6650 7703 6678
rect 7731 6650 7736 6678
rect 12256 6650 12261 6678
rect 12289 6650 12313 6678
rect 12341 6650 12365 6678
rect 12393 6650 12398 6678
rect 16918 6650 16923 6678
rect 16951 6650 16975 6678
rect 17003 6650 17027 6678
rect 17055 6650 17060 6678
rect 5263 6258 5268 6286
rect 5296 6258 5320 6286
rect 5348 6258 5372 6286
rect 5400 6258 5405 6286
rect 9925 6258 9930 6286
rect 9958 6258 9982 6286
rect 10010 6258 10034 6286
rect 10062 6258 10067 6286
rect 14587 6258 14592 6286
rect 14620 6258 14644 6286
rect 14672 6258 14696 6286
rect 14724 6258 14729 6286
rect 19249 6258 19254 6286
rect 19282 6258 19306 6286
rect 19334 6258 19358 6286
rect 19386 6258 19391 6286
rect 7849 6006 7854 6034
rect 7882 6006 8414 6034
rect 8442 6006 8447 6034
rect 10313 5894 10318 5922
rect 10346 5894 11214 5922
rect 11242 5894 11247 5922
rect 2932 5866 2937 5894
rect 2965 5866 2989 5894
rect 3017 5866 3041 5894
rect 3069 5866 3074 5894
rect 7594 5866 7599 5894
rect 7627 5866 7651 5894
rect 7679 5866 7703 5894
rect 7731 5866 7736 5894
rect 12256 5866 12261 5894
rect 12289 5866 12313 5894
rect 12341 5866 12365 5894
rect 12393 5866 12398 5894
rect 16918 5866 16923 5894
rect 16951 5866 16975 5894
rect 17003 5866 17027 5894
rect 17055 5866 17060 5894
rect 5263 5474 5268 5502
rect 5296 5474 5320 5502
rect 5348 5474 5372 5502
rect 5400 5474 5405 5502
rect 9925 5474 9930 5502
rect 9958 5474 9982 5502
rect 10010 5474 10034 5502
rect 10062 5474 10067 5502
rect 14587 5474 14592 5502
rect 14620 5474 14644 5502
rect 14672 5474 14696 5502
rect 14724 5474 14729 5502
rect 19249 5474 19254 5502
rect 19282 5474 19306 5502
rect 19334 5474 19358 5502
rect 19386 5474 19391 5502
rect 2932 5082 2937 5110
rect 2965 5082 2989 5110
rect 3017 5082 3041 5110
rect 3069 5082 3074 5110
rect 7594 5082 7599 5110
rect 7627 5082 7651 5110
rect 7679 5082 7703 5110
rect 7731 5082 7736 5110
rect 12256 5082 12261 5110
rect 12289 5082 12313 5110
rect 12341 5082 12365 5110
rect 12393 5082 12398 5110
rect 16918 5082 16923 5110
rect 16951 5082 16975 5110
rect 17003 5082 17027 5110
rect 17055 5082 17060 5110
rect 5263 4690 5268 4718
rect 5296 4690 5320 4718
rect 5348 4690 5372 4718
rect 5400 4690 5405 4718
rect 9925 4690 9930 4718
rect 9958 4690 9982 4718
rect 10010 4690 10034 4718
rect 10062 4690 10067 4718
rect 14587 4690 14592 4718
rect 14620 4690 14644 4718
rect 14672 4690 14696 4718
rect 14724 4690 14729 4718
rect 19249 4690 19254 4718
rect 19282 4690 19306 4718
rect 19334 4690 19358 4718
rect 19386 4690 19391 4718
rect 2932 4298 2937 4326
rect 2965 4298 2989 4326
rect 3017 4298 3041 4326
rect 3069 4298 3074 4326
rect 7594 4298 7599 4326
rect 7627 4298 7651 4326
rect 7679 4298 7703 4326
rect 7731 4298 7736 4326
rect 12256 4298 12261 4326
rect 12289 4298 12313 4326
rect 12341 4298 12365 4326
rect 12393 4298 12398 4326
rect 16918 4298 16923 4326
rect 16951 4298 16975 4326
rect 17003 4298 17027 4326
rect 17055 4298 17060 4326
rect 5263 3906 5268 3934
rect 5296 3906 5320 3934
rect 5348 3906 5372 3934
rect 5400 3906 5405 3934
rect 9925 3906 9930 3934
rect 9958 3906 9982 3934
rect 10010 3906 10034 3934
rect 10062 3906 10067 3934
rect 14587 3906 14592 3934
rect 14620 3906 14644 3934
rect 14672 3906 14696 3934
rect 14724 3906 14729 3934
rect 19249 3906 19254 3934
rect 19282 3906 19306 3934
rect 19334 3906 19358 3934
rect 19386 3906 19391 3934
rect 2932 3514 2937 3542
rect 2965 3514 2989 3542
rect 3017 3514 3041 3542
rect 3069 3514 3074 3542
rect 7594 3514 7599 3542
rect 7627 3514 7651 3542
rect 7679 3514 7703 3542
rect 7731 3514 7736 3542
rect 12256 3514 12261 3542
rect 12289 3514 12313 3542
rect 12341 3514 12365 3542
rect 12393 3514 12398 3542
rect 16918 3514 16923 3542
rect 16951 3514 16975 3542
rect 17003 3514 17027 3542
rect 17055 3514 17060 3542
rect 5263 3122 5268 3150
rect 5296 3122 5320 3150
rect 5348 3122 5372 3150
rect 5400 3122 5405 3150
rect 9925 3122 9930 3150
rect 9958 3122 9982 3150
rect 10010 3122 10034 3150
rect 10062 3122 10067 3150
rect 14587 3122 14592 3150
rect 14620 3122 14644 3150
rect 14672 3122 14696 3150
rect 14724 3122 14729 3150
rect 19249 3122 19254 3150
rect 19282 3122 19306 3150
rect 19334 3122 19358 3150
rect 19386 3122 19391 3150
rect 2932 2730 2937 2758
rect 2965 2730 2989 2758
rect 3017 2730 3041 2758
rect 3069 2730 3074 2758
rect 7594 2730 7599 2758
rect 7627 2730 7651 2758
rect 7679 2730 7703 2758
rect 7731 2730 7736 2758
rect 12256 2730 12261 2758
rect 12289 2730 12313 2758
rect 12341 2730 12365 2758
rect 12393 2730 12398 2758
rect 16918 2730 16923 2758
rect 16951 2730 16975 2758
rect 17003 2730 17027 2758
rect 17055 2730 17060 2758
rect 9865 2478 9870 2506
rect 9898 2478 11382 2506
rect 11410 2478 11415 2506
rect 5263 2338 5268 2366
rect 5296 2338 5320 2366
rect 5348 2338 5372 2366
rect 5400 2338 5405 2366
rect 9925 2338 9930 2366
rect 9958 2338 9982 2366
rect 10010 2338 10034 2366
rect 10062 2338 10067 2366
rect 14587 2338 14592 2366
rect 14620 2338 14644 2366
rect 14672 2338 14696 2366
rect 14724 2338 14729 2366
rect 19249 2338 19254 2366
rect 19282 2338 19306 2366
rect 19334 2338 19358 2366
rect 19386 2338 19391 2366
rect 7289 2254 7294 2282
rect 7322 2254 8190 2282
rect 8218 2254 8223 2282
rect 9417 2254 9422 2282
rect 9450 2254 9926 2282
rect 9954 2254 9959 2282
rect 6505 2086 6510 2114
rect 6538 2086 6846 2114
rect 6874 2086 6879 2114
rect 12105 2030 12110 2058
rect 12138 2030 13118 2058
rect 13146 2030 13151 2058
rect 2932 1946 2937 1974
rect 2965 1946 2989 1974
rect 3017 1946 3041 1974
rect 3069 1946 3074 1974
rect 7594 1946 7599 1974
rect 7627 1946 7651 1974
rect 7679 1946 7703 1974
rect 7731 1946 7736 1974
rect 12256 1946 12261 1974
rect 12289 1946 12313 1974
rect 12341 1946 12365 1974
rect 12393 1946 12398 1974
rect 16918 1946 16923 1974
rect 16951 1946 16975 1974
rect 17003 1946 17027 1974
rect 17055 1946 17060 1974
rect 11769 1806 11774 1834
rect 11802 1806 12782 1834
rect 12810 1806 12815 1834
rect 7793 1750 7798 1778
rect 7826 1750 8134 1778
rect 8162 1750 8167 1778
rect 8017 1694 8022 1722
rect 8050 1694 8358 1722
rect 8386 1694 8391 1722
rect 10761 1694 10766 1722
rect 10794 1694 10990 1722
rect 11018 1694 11023 1722
rect 5263 1554 5268 1582
rect 5296 1554 5320 1582
rect 5348 1554 5372 1582
rect 5400 1554 5405 1582
rect 9925 1554 9930 1582
rect 9958 1554 9982 1582
rect 10010 1554 10034 1582
rect 10062 1554 10067 1582
rect 14587 1554 14592 1582
rect 14620 1554 14644 1582
rect 14672 1554 14696 1582
rect 14724 1554 14729 1582
rect 19249 1554 19254 1582
rect 19282 1554 19306 1582
rect 19334 1554 19358 1582
rect 19386 1554 19391 1582
<< via3 >>
rect 2937 18410 2965 18438
rect 2989 18410 3017 18438
rect 3041 18410 3069 18438
rect 7599 18410 7627 18438
rect 7651 18410 7679 18438
rect 7703 18410 7731 18438
rect 12261 18410 12289 18438
rect 12313 18410 12341 18438
rect 12365 18410 12393 18438
rect 16923 18410 16951 18438
rect 16975 18410 17003 18438
rect 17027 18410 17055 18438
rect 5268 18018 5296 18046
rect 5320 18018 5348 18046
rect 5372 18018 5400 18046
rect 9930 18018 9958 18046
rect 9982 18018 10010 18046
rect 10034 18018 10062 18046
rect 14592 18018 14620 18046
rect 14644 18018 14672 18046
rect 14696 18018 14724 18046
rect 19254 18018 19282 18046
rect 19306 18018 19334 18046
rect 19358 18018 19386 18046
rect 2937 17626 2965 17654
rect 2989 17626 3017 17654
rect 3041 17626 3069 17654
rect 7599 17626 7627 17654
rect 7651 17626 7679 17654
rect 7703 17626 7731 17654
rect 12261 17626 12289 17654
rect 12313 17626 12341 17654
rect 12365 17626 12393 17654
rect 16923 17626 16951 17654
rect 16975 17626 17003 17654
rect 17027 17626 17055 17654
rect 5268 17234 5296 17262
rect 5320 17234 5348 17262
rect 5372 17234 5400 17262
rect 9930 17234 9958 17262
rect 9982 17234 10010 17262
rect 10034 17234 10062 17262
rect 14592 17234 14620 17262
rect 14644 17234 14672 17262
rect 14696 17234 14724 17262
rect 19254 17234 19282 17262
rect 19306 17234 19334 17262
rect 19358 17234 19386 17262
rect 2937 16842 2965 16870
rect 2989 16842 3017 16870
rect 3041 16842 3069 16870
rect 7599 16842 7627 16870
rect 7651 16842 7679 16870
rect 7703 16842 7731 16870
rect 12261 16842 12289 16870
rect 12313 16842 12341 16870
rect 12365 16842 12393 16870
rect 16923 16842 16951 16870
rect 16975 16842 17003 16870
rect 17027 16842 17055 16870
rect 5268 16450 5296 16478
rect 5320 16450 5348 16478
rect 5372 16450 5400 16478
rect 9930 16450 9958 16478
rect 9982 16450 10010 16478
rect 10034 16450 10062 16478
rect 14592 16450 14620 16478
rect 14644 16450 14672 16478
rect 14696 16450 14724 16478
rect 19254 16450 19282 16478
rect 19306 16450 19334 16478
rect 19358 16450 19386 16478
rect 2937 16058 2965 16086
rect 2989 16058 3017 16086
rect 3041 16058 3069 16086
rect 7599 16058 7627 16086
rect 7651 16058 7679 16086
rect 7703 16058 7731 16086
rect 12261 16058 12289 16086
rect 12313 16058 12341 16086
rect 12365 16058 12393 16086
rect 16923 16058 16951 16086
rect 16975 16058 17003 16086
rect 17027 16058 17055 16086
rect 5268 15666 5296 15694
rect 5320 15666 5348 15694
rect 5372 15666 5400 15694
rect 9930 15666 9958 15694
rect 9982 15666 10010 15694
rect 10034 15666 10062 15694
rect 14592 15666 14620 15694
rect 14644 15666 14672 15694
rect 14696 15666 14724 15694
rect 19254 15666 19282 15694
rect 19306 15666 19334 15694
rect 19358 15666 19386 15694
rect 2937 15274 2965 15302
rect 2989 15274 3017 15302
rect 3041 15274 3069 15302
rect 7599 15274 7627 15302
rect 7651 15274 7679 15302
rect 7703 15274 7731 15302
rect 12261 15274 12289 15302
rect 12313 15274 12341 15302
rect 12365 15274 12393 15302
rect 16923 15274 16951 15302
rect 16975 15274 17003 15302
rect 17027 15274 17055 15302
rect 5268 14882 5296 14910
rect 5320 14882 5348 14910
rect 5372 14882 5400 14910
rect 9930 14882 9958 14910
rect 9982 14882 10010 14910
rect 10034 14882 10062 14910
rect 14592 14882 14620 14910
rect 14644 14882 14672 14910
rect 14696 14882 14724 14910
rect 19254 14882 19282 14910
rect 19306 14882 19334 14910
rect 19358 14882 19386 14910
rect 2937 14490 2965 14518
rect 2989 14490 3017 14518
rect 3041 14490 3069 14518
rect 7599 14490 7627 14518
rect 7651 14490 7679 14518
rect 7703 14490 7731 14518
rect 12261 14490 12289 14518
rect 12313 14490 12341 14518
rect 12365 14490 12393 14518
rect 16923 14490 16951 14518
rect 16975 14490 17003 14518
rect 17027 14490 17055 14518
rect 5268 14098 5296 14126
rect 5320 14098 5348 14126
rect 5372 14098 5400 14126
rect 9930 14098 9958 14126
rect 9982 14098 10010 14126
rect 10034 14098 10062 14126
rect 14592 14098 14620 14126
rect 14644 14098 14672 14126
rect 14696 14098 14724 14126
rect 19254 14098 19282 14126
rect 19306 14098 19334 14126
rect 19358 14098 19386 14126
rect 2937 13706 2965 13734
rect 2989 13706 3017 13734
rect 3041 13706 3069 13734
rect 7599 13706 7627 13734
rect 7651 13706 7679 13734
rect 7703 13706 7731 13734
rect 12261 13706 12289 13734
rect 12313 13706 12341 13734
rect 12365 13706 12393 13734
rect 16923 13706 16951 13734
rect 16975 13706 17003 13734
rect 17027 13706 17055 13734
rect 5268 13314 5296 13342
rect 5320 13314 5348 13342
rect 5372 13314 5400 13342
rect 9930 13314 9958 13342
rect 9982 13314 10010 13342
rect 10034 13314 10062 13342
rect 14592 13314 14620 13342
rect 14644 13314 14672 13342
rect 14696 13314 14724 13342
rect 19254 13314 19282 13342
rect 19306 13314 19334 13342
rect 19358 13314 19386 13342
rect 2937 12922 2965 12950
rect 2989 12922 3017 12950
rect 3041 12922 3069 12950
rect 7599 12922 7627 12950
rect 7651 12922 7679 12950
rect 7703 12922 7731 12950
rect 12261 12922 12289 12950
rect 12313 12922 12341 12950
rect 12365 12922 12393 12950
rect 16923 12922 16951 12950
rect 16975 12922 17003 12950
rect 17027 12922 17055 12950
rect 5268 12530 5296 12558
rect 5320 12530 5348 12558
rect 5372 12530 5400 12558
rect 9930 12530 9958 12558
rect 9982 12530 10010 12558
rect 10034 12530 10062 12558
rect 14592 12530 14620 12558
rect 14644 12530 14672 12558
rect 14696 12530 14724 12558
rect 19254 12530 19282 12558
rect 19306 12530 19334 12558
rect 19358 12530 19386 12558
rect 2937 12138 2965 12166
rect 2989 12138 3017 12166
rect 3041 12138 3069 12166
rect 7599 12138 7627 12166
rect 7651 12138 7679 12166
rect 7703 12138 7731 12166
rect 12261 12138 12289 12166
rect 12313 12138 12341 12166
rect 12365 12138 12393 12166
rect 16923 12138 16951 12166
rect 16975 12138 17003 12166
rect 17027 12138 17055 12166
rect 5268 11746 5296 11774
rect 5320 11746 5348 11774
rect 5372 11746 5400 11774
rect 9930 11746 9958 11774
rect 9982 11746 10010 11774
rect 10034 11746 10062 11774
rect 14592 11746 14620 11774
rect 14644 11746 14672 11774
rect 14696 11746 14724 11774
rect 19254 11746 19282 11774
rect 19306 11746 19334 11774
rect 19358 11746 19386 11774
rect 2937 11354 2965 11382
rect 2989 11354 3017 11382
rect 3041 11354 3069 11382
rect 7599 11354 7627 11382
rect 7651 11354 7679 11382
rect 7703 11354 7731 11382
rect 12261 11354 12289 11382
rect 12313 11354 12341 11382
rect 12365 11354 12393 11382
rect 16923 11354 16951 11382
rect 16975 11354 17003 11382
rect 17027 11354 17055 11382
rect 5268 10962 5296 10990
rect 5320 10962 5348 10990
rect 5372 10962 5400 10990
rect 9930 10962 9958 10990
rect 9982 10962 10010 10990
rect 10034 10962 10062 10990
rect 14592 10962 14620 10990
rect 14644 10962 14672 10990
rect 14696 10962 14724 10990
rect 19254 10962 19282 10990
rect 19306 10962 19334 10990
rect 19358 10962 19386 10990
rect 2937 10570 2965 10598
rect 2989 10570 3017 10598
rect 3041 10570 3069 10598
rect 7599 10570 7627 10598
rect 7651 10570 7679 10598
rect 7703 10570 7731 10598
rect 12261 10570 12289 10598
rect 12313 10570 12341 10598
rect 12365 10570 12393 10598
rect 16923 10570 16951 10598
rect 16975 10570 17003 10598
rect 17027 10570 17055 10598
rect 5268 10178 5296 10206
rect 5320 10178 5348 10206
rect 5372 10178 5400 10206
rect 9930 10178 9958 10206
rect 9982 10178 10010 10206
rect 10034 10178 10062 10206
rect 14592 10178 14620 10206
rect 14644 10178 14672 10206
rect 14696 10178 14724 10206
rect 19254 10178 19282 10206
rect 19306 10178 19334 10206
rect 19358 10178 19386 10206
rect 2937 9786 2965 9814
rect 2989 9786 3017 9814
rect 3041 9786 3069 9814
rect 7599 9786 7627 9814
rect 7651 9786 7679 9814
rect 7703 9786 7731 9814
rect 12261 9786 12289 9814
rect 12313 9786 12341 9814
rect 12365 9786 12393 9814
rect 16923 9786 16951 9814
rect 16975 9786 17003 9814
rect 17027 9786 17055 9814
rect 5268 9394 5296 9422
rect 5320 9394 5348 9422
rect 5372 9394 5400 9422
rect 9930 9394 9958 9422
rect 9982 9394 10010 9422
rect 10034 9394 10062 9422
rect 14592 9394 14620 9422
rect 14644 9394 14672 9422
rect 14696 9394 14724 9422
rect 19254 9394 19282 9422
rect 19306 9394 19334 9422
rect 19358 9394 19386 9422
rect 2937 9002 2965 9030
rect 2989 9002 3017 9030
rect 3041 9002 3069 9030
rect 7599 9002 7627 9030
rect 7651 9002 7679 9030
rect 7703 9002 7731 9030
rect 12261 9002 12289 9030
rect 12313 9002 12341 9030
rect 12365 9002 12393 9030
rect 16923 9002 16951 9030
rect 16975 9002 17003 9030
rect 17027 9002 17055 9030
rect 5268 8610 5296 8638
rect 5320 8610 5348 8638
rect 5372 8610 5400 8638
rect 9930 8610 9958 8638
rect 9982 8610 10010 8638
rect 10034 8610 10062 8638
rect 14592 8610 14620 8638
rect 14644 8610 14672 8638
rect 14696 8610 14724 8638
rect 19254 8610 19282 8638
rect 19306 8610 19334 8638
rect 19358 8610 19386 8638
rect 2937 8218 2965 8246
rect 2989 8218 3017 8246
rect 3041 8218 3069 8246
rect 7599 8218 7627 8246
rect 7651 8218 7679 8246
rect 7703 8218 7731 8246
rect 12261 8218 12289 8246
rect 12313 8218 12341 8246
rect 12365 8218 12393 8246
rect 16923 8218 16951 8246
rect 16975 8218 17003 8246
rect 17027 8218 17055 8246
rect 5268 7826 5296 7854
rect 5320 7826 5348 7854
rect 5372 7826 5400 7854
rect 9930 7826 9958 7854
rect 9982 7826 10010 7854
rect 10034 7826 10062 7854
rect 14592 7826 14620 7854
rect 14644 7826 14672 7854
rect 14696 7826 14724 7854
rect 19254 7826 19282 7854
rect 19306 7826 19334 7854
rect 19358 7826 19386 7854
rect 2937 7434 2965 7462
rect 2989 7434 3017 7462
rect 3041 7434 3069 7462
rect 7599 7434 7627 7462
rect 7651 7434 7679 7462
rect 7703 7434 7731 7462
rect 12261 7434 12289 7462
rect 12313 7434 12341 7462
rect 12365 7434 12393 7462
rect 16923 7434 16951 7462
rect 16975 7434 17003 7462
rect 17027 7434 17055 7462
rect 5268 7042 5296 7070
rect 5320 7042 5348 7070
rect 5372 7042 5400 7070
rect 9930 7042 9958 7070
rect 9982 7042 10010 7070
rect 10034 7042 10062 7070
rect 14592 7042 14620 7070
rect 14644 7042 14672 7070
rect 14696 7042 14724 7070
rect 19254 7042 19282 7070
rect 19306 7042 19334 7070
rect 19358 7042 19386 7070
rect 2937 6650 2965 6678
rect 2989 6650 3017 6678
rect 3041 6650 3069 6678
rect 7599 6650 7627 6678
rect 7651 6650 7679 6678
rect 7703 6650 7731 6678
rect 12261 6650 12289 6678
rect 12313 6650 12341 6678
rect 12365 6650 12393 6678
rect 16923 6650 16951 6678
rect 16975 6650 17003 6678
rect 17027 6650 17055 6678
rect 5268 6258 5296 6286
rect 5320 6258 5348 6286
rect 5372 6258 5400 6286
rect 9930 6258 9958 6286
rect 9982 6258 10010 6286
rect 10034 6258 10062 6286
rect 14592 6258 14620 6286
rect 14644 6258 14672 6286
rect 14696 6258 14724 6286
rect 19254 6258 19282 6286
rect 19306 6258 19334 6286
rect 19358 6258 19386 6286
rect 2937 5866 2965 5894
rect 2989 5866 3017 5894
rect 3041 5866 3069 5894
rect 7599 5866 7627 5894
rect 7651 5866 7679 5894
rect 7703 5866 7731 5894
rect 12261 5866 12289 5894
rect 12313 5866 12341 5894
rect 12365 5866 12393 5894
rect 16923 5866 16951 5894
rect 16975 5866 17003 5894
rect 17027 5866 17055 5894
rect 5268 5474 5296 5502
rect 5320 5474 5348 5502
rect 5372 5474 5400 5502
rect 9930 5474 9958 5502
rect 9982 5474 10010 5502
rect 10034 5474 10062 5502
rect 14592 5474 14620 5502
rect 14644 5474 14672 5502
rect 14696 5474 14724 5502
rect 19254 5474 19282 5502
rect 19306 5474 19334 5502
rect 19358 5474 19386 5502
rect 2937 5082 2965 5110
rect 2989 5082 3017 5110
rect 3041 5082 3069 5110
rect 7599 5082 7627 5110
rect 7651 5082 7679 5110
rect 7703 5082 7731 5110
rect 12261 5082 12289 5110
rect 12313 5082 12341 5110
rect 12365 5082 12393 5110
rect 16923 5082 16951 5110
rect 16975 5082 17003 5110
rect 17027 5082 17055 5110
rect 5268 4690 5296 4718
rect 5320 4690 5348 4718
rect 5372 4690 5400 4718
rect 9930 4690 9958 4718
rect 9982 4690 10010 4718
rect 10034 4690 10062 4718
rect 14592 4690 14620 4718
rect 14644 4690 14672 4718
rect 14696 4690 14724 4718
rect 19254 4690 19282 4718
rect 19306 4690 19334 4718
rect 19358 4690 19386 4718
rect 2937 4298 2965 4326
rect 2989 4298 3017 4326
rect 3041 4298 3069 4326
rect 7599 4298 7627 4326
rect 7651 4298 7679 4326
rect 7703 4298 7731 4326
rect 12261 4298 12289 4326
rect 12313 4298 12341 4326
rect 12365 4298 12393 4326
rect 16923 4298 16951 4326
rect 16975 4298 17003 4326
rect 17027 4298 17055 4326
rect 5268 3906 5296 3934
rect 5320 3906 5348 3934
rect 5372 3906 5400 3934
rect 9930 3906 9958 3934
rect 9982 3906 10010 3934
rect 10034 3906 10062 3934
rect 14592 3906 14620 3934
rect 14644 3906 14672 3934
rect 14696 3906 14724 3934
rect 19254 3906 19282 3934
rect 19306 3906 19334 3934
rect 19358 3906 19386 3934
rect 2937 3514 2965 3542
rect 2989 3514 3017 3542
rect 3041 3514 3069 3542
rect 7599 3514 7627 3542
rect 7651 3514 7679 3542
rect 7703 3514 7731 3542
rect 12261 3514 12289 3542
rect 12313 3514 12341 3542
rect 12365 3514 12393 3542
rect 16923 3514 16951 3542
rect 16975 3514 17003 3542
rect 17027 3514 17055 3542
rect 5268 3122 5296 3150
rect 5320 3122 5348 3150
rect 5372 3122 5400 3150
rect 9930 3122 9958 3150
rect 9982 3122 10010 3150
rect 10034 3122 10062 3150
rect 14592 3122 14620 3150
rect 14644 3122 14672 3150
rect 14696 3122 14724 3150
rect 19254 3122 19282 3150
rect 19306 3122 19334 3150
rect 19358 3122 19386 3150
rect 2937 2730 2965 2758
rect 2989 2730 3017 2758
rect 3041 2730 3069 2758
rect 7599 2730 7627 2758
rect 7651 2730 7679 2758
rect 7703 2730 7731 2758
rect 12261 2730 12289 2758
rect 12313 2730 12341 2758
rect 12365 2730 12393 2758
rect 16923 2730 16951 2758
rect 16975 2730 17003 2758
rect 17027 2730 17055 2758
rect 5268 2338 5296 2366
rect 5320 2338 5348 2366
rect 5372 2338 5400 2366
rect 9930 2338 9958 2366
rect 9982 2338 10010 2366
rect 10034 2338 10062 2366
rect 14592 2338 14620 2366
rect 14644 2338 14672 2366
rect 14696 2338 14724 2366
rect 19254 2338 19282 2366
rect 19306 2338 19334 2366
rect 19358 2338 19386 2366
rect 2937 1946 2965 1974
rect 2989 1946 3017 1974
rect 3041 1946 3069 1974
rect 7599 1946 7627 1974
rect 7651 1946 7679 1974
rect 7703 1946 7731 1974
rect 12261 1946 12289 1974
rect 12313 1946 12341 1974
rect 12365 1946 12393 1974
rect 16923 1946 16951 1974
rect 16975 1946 17003 1974
rect 17027 1946 17055 1974
rect 5268 1554 5296 1582
rect 5320 1554 5348 1582
rect 5372 1554 5400 1582
rect 9930 1554 9958 1582
rect 9982 1554 10010 1582
rect 10034 1554 10062 1582
rect 14592 1554 14620 1582
rect 14644 1554 14672 1582
rect 14696 1554 14724 1582
rect 19254 1554 19282 1582
rect 19306 1554 19334 1582
rect 19358 1554 19386 1582
<< metal4 >>
rect 2923 18438 3083 18454
rect 2923 18410 2937 18438
rect 2965 18410 2989 18438
rect 3017 18410 3041 18438
rect 3069 18410 3083 18438
rect 2923 17654 3083 18410
rect 2923 17626 2937 17654
rect 2965 17626 2989 17654
rect 3017 17626 3041 17654
rect 3069 17626 3083 17654
rect 2923 16870 3083 17626
rect 2923 16842 2937 16870
rect 2965 16842 2989 16870
rect 3017 16842 3041 16870
rect 3069 16842 3083 16870
rect 2923 16086 3083 16842
rect 2923 16058 2937 16086
rect 2965 16058 2989 16086
rect 3017 16058 3041 16086
rect 3069 16058 3083 16086
rect 2923 15302 3083 16058
rect 2923 15274 2937 15302
rect 2965 15274 2989 15302
rect 3017 15274 3041 15302
rect 3069 15274 3083 15302
rect 2923 14518 3083 15274
rect 2923 14490 2937 14518
rect 2965 14490 2989 14518
rect 3017 14490 3041 14518
rect 3069 14490 3083 14518
rect 2923 13734 3083 14490
rect 2923 13706 2937 13734
rect 2965 13706 2989 13734
rect 3017 13706 3041 13734
rect 3069 13706 3083 13734
rect 2923 12950 3083 13706
rect 2923 12922 2937 12950
rect 2965 12922 2989 12950
rect 3017 12922 3041 12950
rect 3069 12922 3083 12950
rect 2923 12166 3083 12922
rect 2923 12138 2937 12166
rect 2965 12138 2989 12166
rect 3017 12138 3041 12166
rect 3069 12138 3083 12166
rect 2923 11382 3083 12138
rect 2923 11354 2937 11382
rect 2965 11354 2989 11382
rect 3017 11354 3041 11382
rect 3069 11354 3083 11382
rect 2923 10598 3083 11354
rect 2923 10570 2937 10598
rect 2965 10570 2989 10598
rect 3017 10570 3041 10598
rect 3069 10570 3083 10598
rect 2923 9814 3083 10570
rect 2923 9786 2937 9814
rect 2965 9786 2989 9814
rect 3017 9786 3041 9814
rect 3069 9786 3083 9814
rect 2923 9030 3083 9786
rect 2923 9002 2937 9030
rect 2965 9002 2989 9030
rect 3017 9002 3041 9030
rect 3069 9002 3083 9030
rect 2923 8246 3083 9002
rect 2923 8218 2937 8246
rect 2965 8218 2989 8246
rect 3017 8218 3041 8246
rect 3069 8218 3083 8246
rect 2923 7462 3083 8218
rect 2923 7434 2937 7462
rect 2965 7434 2989 7462
rect 3017 7434 3041 7462
rect 3069 7434 3083 7462
rect 2923 6678 3083 7434
rect 2923 6650 2937 6678
rect 2965 6650 2989 6678
rect 3017 6650 3041 6678
rect 3069 6650 3083 6678
rect 2923 5894 3083 6650
rect 2923 5866 2937 5894
rect 2965 5866 2989 5894
rect 3017 5866 3041 5894
rect 3069 5866 3083 5894
rect 2923 5110 3083 5866
rect 2923 5082 2937 5110
rect 2965 5082 2989 5110
rect 3017 5082 3041 5110
rect 3069 5082 3083 5110
rect 2923 4326 3083 5082
rect 2923 4298 2937 4326
rect 2965 4298 2989 4326
rect 3017 4298 3041 4326
rect 3069 4298 3083 4326
rect 2923 3542 3083 4298
rect 2923 3514 2937 3542
rect 2965 3514 2989 3542
rect 3017 3514 3041 3542
rect 3069 3514 3083 3542
rect 2923 2758 3083 3514
rect 2923 2730 2937 2758
rect 2965 2730 2989 2758
rect 3017 2730 3041 2758
rect 3069 2730 3083 2758
rect 2923 1974 3083 2730
rect 2923 1946 2937 1974
rect 2965 1946 2989 1974
rect 3017 1946 3041 1974
rect 3069 1946 3083 1974
rect 2923 1538 3083 1946
rect 5254 18046 5414 18454
rect 5254 18018 5268 18046
rect 5296 18018 5320 18046
rect 5348 18018 5372 18046
rect 5400 18018 5414 18046
rect 5254 17262 5414 18018
rect 5254 17234 5268 17262
rect 5296 17234 5320 17262
rect 5348 17234 5372 17262
rect 5400 17234 5414 17262
rect 5254 16478 5414 17234
rect 5254 16450 5268 16478
rect 5296 16450 5320 16478
rect 5348 16450 5372 16478
rect 5400 16450 5414 16478
rect 5254 15694 5414 16450
rect 5254 15666 5268 15694
rect 5296 15666 5320 15694
rect 5348 15666 5372 15694
rect 5400 15666 5414 15694
rect 5254 14910 5414 15666
rect 5254 14882 5268 14910
rect 5296 14882 5320 14910
rect 5348 14882 5372 14910
rect 5400 14882 5414 14910
rect 5254 14126 5414 14882
rect 5254 14098 5268 14126
rect 5296 14098 5320 14126
rect 5348 14098 5372 14126
rect 5400 14098 5414 14126
rect 5254 13342 5414 14098
rect 5254 13314 5268 13342
rect 5296 13314 5320 13342
rect 5348 13314 5372 13342
rect 5400 13314 5414 13342
rect 5254 12558 5414 13314
rect 5254 12530 5268 12558
rect 5296 12530 5320 12558
rect 5348 12530 5372 12558
rect 5400 12530 5414 12558
rect 5254 11774 5414 12530
rect 5254 11746 5268 11774
rect 5296 11746 5320 11774
rect 5348 11746 5372 11774
rect 5400 11746 5414 11774
rect 5254 10990 5414 11746
rect 5254 10962 5268 10990
rect 5296 10962 5320 10990
rect 5348 10962 5372 10990
rect 5400 10962 5414 10990
rect 5254 10206 5414 10962
rect 5254 10178 5268 10206
rect 5296 10178 5320 10206
rect 5348 10178 5372 10206
rect 5400 10178 5414 10206
rect 5254 9422 5414 10178
rect 5254 9394 5268 9422
rect 5296 9394 5320 9422
rect 5348 9394 5372 9422
rect 5400 9394 5414 9422
rect 5254 8638 5414 9394
rect 5254 8610 5268 8638
rect 5296 8610 5320 8638
rect 5348 8610 5372 8638
rect 5400 8610 5414 8638
rect 5254 7854 5414 8610
rect 5254 7826 5268 7854
rect 5296 7826 5320 7854
rect 5348 7826 5372 7854
rect 5400 7826 5414 7854
rect 5254 7070 5414 7826
rect 5254 7042 5268 7070
rect 5296 7042 5320 7070
rect 5348 7042 5372 7070
rect 5400 7042 5414 7070
rect 5254 6286 5414 7042
rect 5254 6258 5268 6286
rect 5296 6258 5320 6286
rect 5348 6258 5372 6286
rect 5400 6258 5414 6286
rect 5254 5502 5414 6258
rect 5254 5474 5268 5502
rect 5296 5474 5320 5502
rect 5348 5474 5372 5502
rect 5400 5474 5414 5502
rect 5254 4718 5414 5474
rect 5254 4690 5268 4718
rect 5296 4690 5320 4718
rect 5348 4690 5372 4718
rect 5400 4690 5414 4718
rect 5254 3934 5414 4690
rect 5254 3906 5268 3934
rect 5296 3906 5320 3934
rect 5348 3906 5372 3934
rect 5400 3906 5414 3934
rect 5254 3150 5414 3906
rect 5254 3122 5268 3150
rect 5296 3122 5320 3150
rect 5348 3122 5372 3150
rect 5400 3122 5414 3150
rect 5254 2366 5414 3122
rect 5254 2338 5268 2366
rect 5296 2338 5320 2366
rect 5348 2338 5372 2366
rect 5400 2338 5414 2366
rect 5254 1582 5414 2338
rect 5254 1554 5268 1582
rect 5296 1554 5320 1582
rect 5348 1554 5372 1582
rect 5400 1554 5414 1582
rect 5254 1538 5414 1554
rect 7585 18438 7745 18454
rect 7585 18410 7599 18438
rect 7627 18410 7651 18438
rect 7679 18410 7703 18438
rect 7731 18410 7745 18438
rect 7585 17654 7745 18410
rect 7585 17626 7599 17654
rect 7627 17626 7651 17654
rect 7679 17626 7703 17654
rect 7731 17626 7745 17654
rect 7585 16870 7745 17626
rect 7585 16842 7599 16870
rect 7627 16842 7651 16870
rect 7679 16842 7703 16870
rect 7731 16842 7745 16870
rect 7585 16086 7745 16842
rect 7585 16058 7599 16086
rect 7627 16058 7651 16086
rect 7679 16058 7703 16086
rect 7731 16058 7745 16086
rect 7585 15302 7745 16058
rect 7585 15274 7599 15302
rect 7627 15274 7651 15302
rect 7679 15274 7703 15302
rect 7731 15274 7745 15302
rect 7585 14518 7745 15274
rect 7585 14490 7599 14518
rect 7627 14490 7651 14518
rect 7679 14490 7703 14518
rect 7731 14490 7745 14518
rect 7585 13734 7745 14490
rect 7585 13706 7599 13734
rect 7627 13706 7651 13734
rect 7679 13706 7703 13734
rect 7731 13706 7745 13734
rect 7585 12950 7745 13706
rect 7585 12922 7599 12950
rect 7627 12922 7651 12950
rect 7679 12922 7703 12950
rect 7731 12922 7745 12950
rect 7585 12166 7745 12922
rect 7585 12138 7599 12166
rect 7627 12138 7651 12166
rect 7679 12138 7703 12166
rect 7731 12138 7745 12166
rect 7585 11382 7745 12138
rect 7585 11354 7599 11382
rect 7627 11354 7651 11382
rect 7679 11354 7703 11382
rect 7731 11354 7745 11382
rect 7585 10598 7745 11354
rect 7585 10570 7599 10598
rect 7627 10570 7651 10598
rect 7679 10570 7703 10598
rect 7731 10570 7745 10598
rect 7585 9814 7745 10570
rect 7585 9786 7599 9814
rect 7627 9786 7651 9814
rect 7679 9786 7703 9814
rect 7731 9786 7745 9814
rect 7585 9030 7745 9786
rect 7585 9002 7599 9030
rect 7627 9002 7651 9030
rect 7679 9002 7703 9030
rect 7731 9002 7745 9030
rect 7585 8246 7745 9002
rect 7585 8218 7599 8246
rect 7627 8218 7651 8246
rect 7679 8218 7703 8246
rect 7731 8218 7745 8246
rect 7585 7462 7745 8218
rect 7585 7434 7599 7462
rect 7627 7434 7651 7462
rect 7679 7434 7703 7462
rect 7731 7434 7745 7462
rect 7585 6678 7745 7434
rect 7585 6650 7599 6678
rect 7627 6650 7651 6678
rect 7679 6650 7703 6678
rect 7731 6650 7745 6678
rect 7585 5894 7745 6650
rect 7585 5866 7599 5894
rect 7627 5866 7651 5894
rect 7679 5866 7703 5894
rect 7731 5866 7745 5894
rect 7585 5110 7745 5866
rect 7585 5082 7599 5110
rect 7627 5082 7651 5110
rect 7679 5082 7703 5110
rect 7731 5082 7745 5110
rect 7585 4326 7745 5082
rect 7585 4298 7599 4326
rect 7627 4298 7651 4326
rect 7679 4298 7703 4326
rect 7731 4298 7745 4326
rect 7585 3542 7745 4298
rect 7585 3514 7599 3542
rect 7627 3514 7651 3542
rect 7679 3514 7703 3542
rect 7731 3514 7745 3542
rect 7585 2758 7745 3514
rect 7585 2730 7599 2758
rect 7627 2730 7651 2758
rect 7679 2730 7703 2758
rect 7731 2730 7745 2758
rect 7585 1974 7745 2730
rect 7585 1946 7599 1974
rect 7627 1946 7651 1974
rect 7679 1946 7703 1974
rect 7731 1946 7745 1974
rect 7585 1538 7745 1946
rect 9916 18046 10076 18454
rect 9916 18018 9930 18046
rect 9958 18018 9982 18046
rect 10010 18018 10034 18046
rect 10062 18018 10076 18046
rect 9916 17262 10076 18018
rect 9916 17234 9930 17262
rect 9958 17234 9982 17262
rect 10010 17234 10034 17262
rect 10062 17234 10076 17262
rect 9916 16478 10076 17234
rect 9916 16450 9930 16478
rect 9958 16450 9982 16478
rect 10010 16450 10034 16478
rect 10062 16450 10076 16478
rect 9916 15694 10076 16450
rect 9916 15666 9930 15694
rect 9958 15666 9982 15694
rect 10010 15666 10034 15694
rect 10062 15666 10076 15694
rect 9916 14910 10076 15666
rect 9916 14882 9930 14910
rect 9958 14882 9982 14910
rect 10010 14882 10034 14910
rect 10062 14882 10076 14910
rect 9916 14126 10076 14882
rect 9916 14098 9930 14126
rect 9958 14098 9982 14126
rect 10010 14098 10034 14126
rect 10062 14098 10076 14126
rect 9916 13342 10076 14098
rect 9916 13314 9930 13342
rect 9958 13314 9982 13342
rect 10010 13314 10034 13342
rect 10062 13314 10076 13342
rect 9916 12558 10076 13314
rect 9916 12530 9930 12558
rect 9958 12530 9982 12558
rect 10010 12530 10034 12558
rect 10062 12530 10076 12558
rect 9916 11774 10076 12530
rect 9916 11746 9930 11774
rect 9958 11746 9982 11774
rect 10010 11746 10034 11774
rect 10062 11746 10076 11774
rect 9916 10990 10076 11746
rect 9916 10962 9930 10990
rect 9958 10962 9982 10990
rect 10010 10962 10034 10990
rect 10062 10962 10076 10990
rect 9916 10206 10076 10962
rect 9916 10178 9930 10206
rect 9958 10178 9982 10206
rect 10010 10178 10034 10206
rect 10062 10178 10076 10206
rect 9916 9422 10076 10178
rect 9916 9394 9930 9422
rect 9958 9394 9982 9422
rect 10010 9394 10034 9422
rect 10062 9394 10076 9422
rect 9916 8638 10076 9394
rect 9916 8610 9930 8638
rect 9958 8610 9982 8638
rect 10010 8610 10034 8638
rect 10062 8610 10076 8638
rect 9916 7854 10076 8610
rect 9916 7826 9930 7854
rect 9958 7826 9982 7854
rect 10010 7826 10034 7854
rect 10062 7826 10076 7854
rect 9916 7070 10076 7826
rect 9916 7042 9930 7070
rect 9958 7042 9982 7070
rect 10010 7042 10034 7070
rect 10062 7042 10076 7070
rect 9916 6286 10076 7042
rect 9916 6258 9930 6286
rect 9958 6258 9982 6286
rect 10010 6258 10034 6286
rect 10062 6258 10076 6286
rect 9916 5502 10076 6258
rect 9916 5474 9930 5502
rect 9958 5474 9982 5502
rect 10010 5474 10034 5502
rect 10062 5474 10076 5502
rect 9916 4718 10076 5474
rect 9916 4690 9930 4718
rect 9958 4690 9982 4718
rect 10010 4690 10034 4718
rect 10062 4690 10076 4718
rect 9916 3934 10076 4690
rect 9916 3906 9930 3934
rect 9958 3906 9982 3934
rect 10010 3906 10034 3934
rect 10062 3906 10076 3934
rect 9916 3150 10076 3906
rect 9916 3122 9930 3150
rect 9958 3122 9982 3150
rect 10010 3122 10034 3150
rect 10062 3122 10076 3150
rect 9916 2366 10076 3122
rect 9916 2338 9930 2366
rect 9958 2338 9982 2366
rect 10010 2338 10034 2366
rect 10062 2338 10076 2366
rect 9916 1582 10076 2338
rect 9916 1554 9930 1582
rect 9958 1554 9982 1582
rect 10010 1554 10034 1582
rect 10062 1554 10076 1582
rect 9916 1538 10076 1554
rect 12247 18438 12407 18454
rect 12247 18410 12261 18438
rect 12289 18410 12313 18438
rect 12341 18410 12365 18438
rect 12393 18410 12407 18438
rect 12247 17654 12407 18410
rect 12247 17626 12261 17654
rect 12289 17626 12313 17654
rect 12341 17626 12365 17654
rect 12393 17626 12407 17654
rect 12247 16870 12407 17626
rect 12247 16842 12261 16870
rect 12289 16842 12313 16870
rect 12341 16842 12365 16870
rect 12393 16842 12407 16870
rect 12247 16086 12407 16842
rect 12247 16058 12261 16086
rect 12289 16058 12313 16086
rect 12341 16058 12365 16086
rect 12393 16058 12407 16086
rect 12247 15302 12407 16058
rect 12247 15274 12261 15302
rect 12289 15274 12313 15302
rect 12341 15274 12365 15302
rect 12393 15274 12407 15302
rect 12247 14518 12407 15274
rect 12247 14490 12261 14518
rect 12289 14490 12313 14518
rect 12341 14490 12365 14518
rect 12393 14490 12407 14518
rect 12247 13734 12407 14490
rect 12247 13706 12261 13734
rect 12289 13706 12313 13734
rect 12341 13706 12365 13734
rect 12393 13706 12407 13734
rect 12247 12950 12407 13706
rect 12247 12922 12261 12950
rect 12289 12922 12313 12950
rect 12341 12922 12365 12950
rect 12393 12922 12407 12950
rect 12247 12166 12407 12922
rect 12247 12138 12261 12166
rect 12289 12138 12313 12166
rect 12341 12138 12365 12166
rect 12393 12138 12407 12166
rect 12247 11382 12407 12138
rect 12247 11354 12261 11382
rect 12289 11354 12313 11382
rect 12341 11354 12365 11382
rect 12393 11354 12407 11382
rect 12247 10598 12407 11354
rect 12247 10570 12261 10598
rect 12289 10570 12313 10598
rect 12341 10570 12365 10598
rect 12393 10570 12407 10598
rect 12247 9814 12407 10570
rect 12247 9786 12261 9814
rect 12289 9786 12313 9814
rect 12341 9786 12365 9814
rect 12393 9786 12407 9814
rect 12247 9030 12407 9786
rect 12247 9002 12261 9030
rect 12289 9002 12313 9030
rect 12341 9002 12365 9030
rect 12393 9002 12407 9030
rect 12247 8246 12407 9002
rect 12247 8218 12261 8246
rect 12289 8218 12313 8246
rect 12341 8218 12365 8246
rect 12393 8218 12407 8246
rect 12247 7462 12407 8218
rect 12247 7434 12261 7462
rect 12289 7434 12313 7462
rect 12341 7434 12365 7462
rect 12393 7434 12407 7462
rect 12247 6678 12407 7434
rect 12247 6650 12261 6678
rect 12289 6650 12313 6678
rect 12341 6650 12365 6678
rect 12393 6650 12407 6678
rect 12247 5894 12407 6650
rect 12247 5866 12261 5894
rect 12289 5866 12313 5894
rect 12341 5866 12365 5894
rect 12393 5866 12407 5894
rect 12247 5110 12407 5866
rect 12247 5082 12261 5110
rect 12289 5082 12313 5110
rect 12341 5082 12365 5110
rect 12393 5082 12407 5110
rect 12247 4326 12407 5082
rect 12247 4298 12261 4326
rect 12289 4298 12313 4326
rect 12341 4298 12365 4326
rect 12393 4298 12407 4326
rect 12247 3542 12407 4298
rect 12247 3514 12261 3542
rect 12289 3514 12313 3542
rect 12341 3514 12365 3542
rect 12393 3514 12407 3542
rect 12247 2758 12407 3514
rect 12247 2730 12261 2758
rect 12289 2730 12313 2758
rect 12341 2730 12365 2758
rect 12393 2730 12407 2758
rect 12247 1974 12407 2730
rect 12247 1946 12261 1974
rect 12289 1946 12313 1974
rect 12341 1946 12365 1974
rect 12393 1946 12407 1974
rect 12247 1538 12407 1946
rect 14578 18046 14738 18454
rect 14578 18018 14592 18046
rect 14620 18018 14644 18046
rect 14672 18018 14696 18046
rect 14724 18018 14738 18046
rect 14578 17262 14738 18018
rect 14578 17234 14592 17262
rect 14620 17234 14644 17262
rect 14672 17234 14696 17262
rect 14724 17234 14738 17262
rect 14578 16478 14738 17234
rect 14578 16450 14592 16478
rect 14620 16450 14644 16478
rect 14672 16450 14696 16478
rect 14724 16450 14738 16478
rect 14578 15694 14738 16450
rect 14578 15666 14592 15694
rect 14620 15666 14644 15694
rect 14672 15666 14696 15694
rect 14724 15666 14738 15694
rect 14578 14910 14738 15666
rect 14578 14882 14592 14910
rect 14620 14882 14644 14910
rect 14672 14882 14696 14910
rect 14724 14882 14738 14910
rect 14578 14126 14738 14882
rect 14578 14098 14592 14126
rect 14620 14098 14644 14126
rect 14672 14098 14696 14126
rect 14724 14098 14738 14126
rect 14578 13342 14738 14098
rect 14578 13314 14592 13342
rect 14620 13314 14644 13342
rect 14672 13314 14696 13342
rect 14724 13314 14738 13342
rect 14578 12558 14738 13314
rect 14578 12530 14592 12558
rect 14620 12530 14644 12558
rect 14672 12530 14696 12558
rect 14724 12530 14738 12558
rect 14578 11774 14738 12530
rect 14578 11746 14592 11774
rect 14620 11746 14644 11774
rect 14672 11746 14696 11774
rect 14724 11746 14738 11774
rect 14578 10990 14738 11746
rect 14578 10962 14592 10990
rect 14620 10962 14644 10990
rect 14672 10962 14696 10990
rect 14724 10962 14738 10990
rect 14578 10206 14738 10962
rect 14578 10178 14592 10206
rect 14620 10178 14644 10206
rect 14672 10178 14696 10206
rect 14724 10178 14738 10206
rect 14578 9422 14738 10178
rect 14578 9394 14592 9422
rect 14620 9394 14644 9422
rect 14672 9394 14696 9422
rect 14724 9394 14738 9422
rect 14578 8638 14738 9394
rect 14578 8610 14592 8638
rect 14620 8610 14644 8638
rect 14672 8610 14696 8638
rect 14724 8610 14738 8638
rect 14578 7854 14738 8610
rect 14578 7826 14592 7854
rect 14620 7826 14644 7854
rect 14672 7826 14696 7854
rect 14724 7826 14738 7854
rect 14578 7070 14738 7826
rect 14578 7042 14592 7070
rect 14620 7042 14644 7070
rect 14672 7042 14696 7070
rect 14724 7042 14738 7070
rect 14578 6286 14738 7042
rect 14578 6258 14592 6286
rect 14620 6258 14644 6286
rect 14672 6258 14696 6286
rect 14724 6258 14738 6286
rect 14578 5502 14738 6258
rect 14578 5474 14592 5502
rect 14620 5474 14644 5502
rect 14672 5474 14696 5502
rect 14724 5474 14738 5502
rect 14578 4718 14738 5474
rect 14578 4690 14592 4718
rect 14620 4690 14644 4718
rect 14672 4690 14696 4718
rect 14724 4690 14738 4718
rect 14578 3934 14738 4690
rect 14578 3906 14592 3934
rect 14620 3906 14644 3934
rect 14672 3906 14696 3934
rect 14724 3906 14738 3934
rect 14578 3150 14738 3906
rect 14578 3122 14592 3150
rect 14620 3122 14644 3150
rect 14672 3122 14696 3150
rect 14724 3122 14738 3150
rect 14578 2366 14738 3122
rect 14578 2338 14592 2366
rect 14620 2338 14644 2366
rect 14672 2338 14696 2366
rect 14724 2338 14738 2366
rect 14578 1582 14738 2338
rect 14578 1554 14592 1582
rect 14620 1554 14644 1582
rect 14672 1554 14696 1582
rect 14724 1554 14738 1582
rect 14578 1538 14738 1554
rect 16909 18438 17069 18454
rect 16909 18410 16923 18438
rect 16951 18410 16975 18438
rect 17003 18410 17027 18438
rect 17055 18410 17069 18438
rect 16909 17654 17069 18410
rect 16909 17626 16923 17654
rect 16951 17626 16975 17654
rect 17003 17626 17027 17654
rect 17055 17626 17069 17654
rect 16909 16870 17069 17626
rect 16909 16842 16923 16870
rect 16951 16842 16975 16870
rect 17003 16842 17027 16870
rect 17055 16842 17069 16870
rect 16909 16086 17069 16842
rect 16909 16058 16923 16086
rect 16951 16058 16975 16086
rect 17003 16058 17027 16086
rect 17055 16058 17069 16086
rect 16909 15302 17069 16058
rect 16909 15274 16923 15302
rect 16951 15274 16975 15302
rect 17003 15274 17027 15302
rect 17055 15274 17069 15302
rect 16909 14518 17069 15274
rect 16909 14490 16923 14518
rect 16951 14490 16975 14518
rect 17003 14490 17027 14518
rect 17055 14490 17069 14518
rect 16909 13734 17069 14490
rect 16909 13706 16923 13734
rect 16951 13706 16975 13734
rect 17003 13706 17027 13734
rect 17055 13706 17069 13734
rect 16909 12950 17069 13706
rect 16909 12922 16923 12950
rect 16951 12922 16975 12950
rect 17003 12922 17027 12950
rect 17055 12922 17069 12950
rect 16909 12166 17069 12922
rect 16909 12138 16923 12166
rect 16951 12138 16975 12166
rect 17003 12138 17027 12166
rect 17055 12138 17069 12166
rect 16909 11382 17069 12138
rect 16909 11354 16923 11382
rect 16951 11354 16975 11382
rect 17003 11354 17027 11382
rect 17055 11354 17069 11382
rect 16909 10598 17069 11354
rect 16909 10570 16923 10598
rect 16951 10570 16975 10598
rect 17003 10570 17027 10598
rect 17055 10570 17069 10598
rect 16909 9814 17069 10570
rect 16909 9786 16923 9814
rect 16951 9786 16975 9814
rect 17003 9786 17027 9814
rect 17055 9786 17069 9814
rect 16909 9030 17069 9786
rect 16909 9002 16923 9030
rect 16951 9002 16975 9030
rect 17003 9002 17027 9030
rect 17055 9002 17069 9030
rect 16909 8246 17069 9002
rect 16909 8218 16923 8246
rect 16951 8218 16975 8246
rect 17003 8218 17027 8246
rect 17055 8218 17069 8246
rect 16909 7462 17069 8218
rect 16909 7434 16923 7462
rect 16951 7434 16975 7462
rect 17003 7434 17027 7462
rect 17055 7434 17069 7462
rect 16909 6678 17069 7434
rect 16909 6650 16923 6678
rect 16951 6650 16975 6678
rect 17003 6650 17027 6678
rect 17055 6650 17069 6678
rect 16909 5894 17069 6650
rect 16909 5866 16923 5894
rect 16951 5866 16975 5894
rect 17003 5866 17027 5894
rect 17055 5866 17069 5894
rect 16909 5110 17069 5866
rect 16909 5082 16923 5110
rect 16951 5082 16975 5110
rect 17003 5082 17027 5110
rect 17055 5082 17069 5110
rect 16909 4326 17069 5082
rect 16909 4298 16923 4326
rect 16951 4298 16975 4326
rect 17003 4298 17027 4326
rect 17055 4298 17069 4326
rect 16909 3542 17069 4298
rect 16909 3514 16923 3542
rect 16951 3514 16975 3542
rect 17003 3514 17027 3542
rect 17055 3514 17069 3542
rect 16909 2758 17069 3514
rect 16909 2730 16923 2758
rect 16951 2730 16975 2758
rect 17003 2730 17027 2758
rect 17055 2730 17069 2758
rect 16909 1974 17069 2730
rect 16909 1946 16923 1974
rect 16951 1946 16975 1974
rect 17003 1946 17027 1974
rect 17055 1946 17069 1974
rect 16909 1538 17069 1946
rect 19240 18046 19400 18454
rect 19240 18018 19254 18046
rect 19282 18018 19306 18046
rect 19334 18018 19358 18046
rect 19386 18018 19400 18046
rect 19240 17262 19400 18018
rect 19240 17234 19254 17262
rect 19282 17234 19306 17262
rect 19334 17234 19358 17262
rect 19386 17234 19400 17262
rect 19240 16478 19400 17234
rect 19240 16450 19254 16478
rect 19282 16450 19306 16478
rect 19334 16450 19358 16478
rect 19386 16450 19400 16478
rect 19240 15694 19400 16450
rect 19240 15666 19254 15694
rect 19282 15666 19306 15694
rect 19334 15666 19358 15694
rect 19386 15666 19400 15694
rect 19240 14910 19400 15666
rect 19240 14882 19254 14910
rect 19282 14882 19306 14910
rect 19334 14882 19358 14910
rect 19386 14882 19400 14910
rect 19240 14126 19400 14882
rect 19240 14098 19254 14126
rect 19282 14098 19306 14126
rect 19334 14098 19358 14126
rect 19386 14098 19400 14126
rect 19240 13342 19400 14098
rect 19240 13314 19254 13342
rect 19282 13314 19306 13342
rect 19334 13314 19358 13342
rect 19386 13314 19400 13342
rect 19240 12558 19400 13314
rect 19240 12530 19254 12558
rect 19282 12530 19306 12558
rect 19334 12530 19358 12558
rect 19386 12530 19400 12558
rect 19240 11774 19400 12530
rect 19240 11746 19254 11774
rect 19282 11746 19306 11774
rect 19334 11746 19358 11774
rect 19386 11746 19400 11774
rect 19240 10990 19400 11746
rect 19240 10962 19254 10990
rect 19282 10962 19306 10990
rect 19334 10962 19358 10990
rect 19386 10962 19400 10990
rect 19240 10206 19400 10962
rect 19240 10178 19254 10206
rect 19282 10178 19306 10206
rect 19334 10178 19358 10206
rect 19386 10178 19400 10206
rect 19240 9422 19400 10178
rect 19240 9394 19254 9422
rect 19282 9394 19306 9422
rect 19334 9394 19358 9422
rect 19386 9394 19400 9422
rect 19240 8638 19400 9394
rect 19240 8610 19254 8638
rect 19282 8610 19306 8638
rect 19334 8610 19358 8638
rect 19386 8610 19400 8638
rect 19240 7854 19400 8610
rect 19240 7826 19254 7854
rect 19282 7826 19306 7854
rect 19334 7826 19358 7854
rect 19386 7826 19400 7854
rect 19240 7070 19400 7826
rect 19240 7042 19254 7070
rect 19282 7042 19306 7070
rect 19334 7042 19358 7070
rect 19386 7042 19400 7070
rect 19240 6286 19400 7042
rect 19240 6258 19254 6286
rect 19282 6258 19306 6286
rect 19334 6258 19358 6286
rect 19386 6258 19400 6286
rect 19240 5502 19400 6258
rect 19240 5474 19254 5502
rect 19282 5474 19306 5502
rect 19334 5474 19358 5502
rect 19386 5474 19400 5502
rect 19240 4718 19400 5474
rect 19240 4690 19254 4718
rect 19282 4690 19306 4718
rect 19334 4690 19358 4718
rect 19386 4690 19400 4718
rect 19240 3934 19400 4690
rect 19240 3906 19254 3934
rect 19282 3906 19306 3934
rect 19334 3906 19358 3934
rect 19386 3906 19400 3934
rect 19240 3150 19400 3906
rect 19240 3122 19254 3150
rect 19282 3122 19306 3150
rect 19334 3122 19358 3150
rect 19386 3122 19400 3150
rect 19240 2366 19400 3122
rect 19240 2338 19254 2366
rect 19282 2338 19306 2366
rect 19334 2338 19358 2366
rect 19386 2338 19400 2366
rect 19240 1582 19400 2338
rect 19240 1554 19254 1582
rect 19282 1554 19306 1582
rect 19334 1554 19358 1582
rect 19386 1554 19400 1582
rect 19240 1538 19400 1554
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _18_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9576 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _19_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10024 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _20_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10528 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _21_
timestamp 1698431365
transform 1 0 11088 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _22_
timestamp 1698431365
transform 1 0 10584 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _23_
timestamp 1698431365
transform 1 0 11424 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _24_
timestamp 1698431365
transform 1 0 10416 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _25_
timestamp 1698431365
transform 1 0 10976 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _26_
timestamp 1698431365
transform 1 0 10584 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _27_
timestamp 1698431365
transform 1 0 10640 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _28_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _29_
timestamp 1698431365
transform -1 0 9744 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _30_
timestamp 1698431365
transform 1 0 7504 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _31_
timestamp 1698431365
transform -1 0 8232 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _32_
timestamp 1698431365
transform 1 0 8680 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _33_
timestamp 1698431365
transform 1 0 9968 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _34_
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _35_
timestamp 1698431365
transform 1 0 9632 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _36_
timestamp 1698431365
transform -1 0 8512 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _37_
timestamp 1698431365
transform -1 0 8344 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _38_
timestamp 1698431365
transform -1 0 9072 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _39_
timestamp 1698431365
transform -1 0 9408 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _40_
timestamp 1698431365
transform 1 0 7784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _41_
timestamp 1698431365
transform -1 0 8512 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _42_
timestamp 1698431365
transform 1 0 7952 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _43_
timestamp 1698431365
transform -1 0 8960 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _44_
timestamp 1698431365
transform 1 0 7784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _45_
timestamp 1698431365
transform -1 0 8960 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _46_
timestamp 1698431365
transform 1 0 7952 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _47_
timestamp 1698431365
transform -1 0 8960 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__18__I test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9576 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__20__I2
timestamp 1698431365
transform 1 0 12656 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__20__I3
timestamp 1698431365
transform -1 0 12992 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__28__I
timestamp 1698431365
transform 1 0 8624 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__38__I
timestamp 1698431365
transform 1 0 8400 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__40__I0
timestamp 1698431365
transform -1 0 7784 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__44__I2
timestamp 1698431365
transform -1 0 7784 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 18872 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 1232 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 9464 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 18872 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 18872 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 18872 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 8400 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 11480 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 10472 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 8120 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 18760 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 9128 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 1232 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 8792 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 18648 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 18872 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 10192 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 10136 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 896 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 6776 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform -1 0 18872 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 9184 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 7448 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 1232 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 1232 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform 1 0 1232 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 1232 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 18872 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 19208 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 11144 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 10808 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 1568 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform 1 0 9520 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform 1 0 9856 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 7784 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform 1 0 1456 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform -1 0 7560 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform 1 0 1232 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform -1 0 7784 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform 1 0 8848 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform -1 0 11144 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform -1 0 10808 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform -1 0 6552 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform 1 0 1232 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform -1 0 9800 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698431365
transform 1 0 1232 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698431365
transform 1 0 10136 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output51_I
timestamp 1698431365
transform 1 0 17640 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output61_I
timestamp 1698431365
transform -1 0 2464 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8400 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 10304 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10416 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_199 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11816 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 12040 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698431365
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698431365
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_308 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17920 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_324
timestamp 1698431365
transform 1 0 18816 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_328
timestamp 1698431365
transform 1 0 19040 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_330
timestamp 1698431365
transform 1 0 19152 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_72
timestamp 1698431365
transform 1 0 4704 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_88 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5600 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_96
timestamp 1698431365
transform 1 0 6048 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_100
timestamp 1698431365
transform 1 0 6272 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_102
timestamp 1698431365
transform 1 0 6384 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_105
timestamp 1698431365
transform 1 0 6552 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 8456 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_142
timestamp 1698431365
transform 1 0 8624 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_148
timestamp 1698431365
transform 1 0 8960 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_154
timestamp 1698431365
transform 1 0 9296 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_160
timestamp 1698431365
transform 1 0 9632 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_166
timestamp 1698431365
transform 1 0 9968 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_168
timestamp 1698431365
transform 1 0 10080 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_171
timestamp 1698431365
transform 1 0 10248 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_175
timestamp 1698431365
transform 1 0 10472 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_181
timestamp 1698431365
transform 1 0 10808 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_187
timestamp 1698431365
transform 1 0 11144 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_193
timestamp 1698431365
transform 1 0 11480 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698431365
transform 1 0 14000 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698431365
transform 1 0 15792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698431365
transform 1 0 16240 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_282
timestamp 1698431365
transform 1 0 16464 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_314
timestamp 1698431365
transform 1 0 18256 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_330
timestamp 1698431365
transform 1 0 19152 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_107
timestamp 1698431365
transform 1 0 6664 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_115
timestamp 1698431365
transform 1 0 7112 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_121
timestamp 1698431365
transform 1 0 7448 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_127
timestamp 1698431365
transform 1 0 7784 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_133
timestamp 1698431365
transform 1 0 8120 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_135
timestamp 1698431365
transform 1 0 8232 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_138
timestamp 1698431365
transform 1 0 8400 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_170
timestamp 1698431365
transform 1 0 10192 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 10416 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_317
timestamp 1698431365
transform 1 0 18424 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_325
timestamp 1698431365
transform 1 0 18872 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_329
timestamp 1698431365
transform 1 0 19096 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_282
timestamp 1698431365
transform 1 0 16464 0 -1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_314
timestamp 1698431365
transform 1 0 18256 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_330
timestamp 1698431365
transform 1 0 19152 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_317
timestamp 1698431365
transform 1 0 18424 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_325
timestamp 1698431365
transform 1 0 18872 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_329
timestamp 1698431365
transform 1 0 19096 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_282
timestamp 1698431365
transform 1 0 16464 0 -1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_314
timestamp 1698431365
transform 1 0 18256 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_330
timestamp 1698431365
transform 1 0 19152 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698431365
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_317
timestamp 1698431365
transform 1 0 18424 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_325
timestamp 1698431365
transform 1 0 18872 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_329
timestamp 1698431365
transform 1 0 19096 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698431365
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_282
timestamp 1698431365
transform 1 0 16464 0 -1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_314
timestamp 1698431365
transform 1 0 18256 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_330
timestamp 1698431365
transform 1 0 19152 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698431365
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698431365
transform 1 0 18424 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_325
timestamp 1698431365
transform 1 0 18872 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_329
timestamp 1698431365
transform 1 0 19096 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698431365
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_282
timestamp 1698431365
transform 1 0 16464 0 -1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_314
timestamp 1698431365
transform 1 0 18256 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_330
timestamp 1698431365
transform 1 0 19152 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698431365
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698431365
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_317
timestamp 1698431365
transform 1 0 18424 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_325
timestamp 1698431365
transform 1 0 18872 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_329
timestamp 1698431365
transform 1 0 19096 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698431365
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698431365
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_282
timestamp 1698431365
transform 1 0 16464 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_314
timestamp 1698431365
transform 1 0 18256 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_330
timestamp 1698431365
transform 1 0 19152 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698431365
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698431365
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698431365
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_317
timestamp 1698431365
transform 1 0 18424 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_325
timestamp 1698431365
transform 1 0 18872 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_329
timestamp 1698431365
transform 1 0 19096 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698431365
transform 1 0 8624 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 12208 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698431365
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698431365
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_282
timestamp 1698431365
transform 1 0 16464 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_298
timestamp 1698431365
transform 1 0 17360 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_302
timestamp 1698431365
transform 1 0 17584 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698431365
transform 1 0 6664 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698431365
transform 1 0 7560 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_137
timestamp 1698431365
transform 1 0 8344 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_141
timestamp 1698431365
transform 1 0 8568 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698431365
transform 1 0 10584 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698431365
transform 1 0 14168 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698431365
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_317
timestamp 1698431365
transform 1 0 18424 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_321
timestamp 1698431365
transform 1 0 18648 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_2
timestamp 1698431365
transform 1 0 784 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_6
timestamp 1698431365
transform 1 0 1008 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698431365
transform 1 0 4704 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_104
timestamp 1698431365
transform 1 0 6496 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698431365
transform 1 0 8624 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_182
timestamp 1698431365
transform 1 0 10864 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_198
timestamp 1698431365
transform 1 0 11760 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698431365
transform 1 0 12208 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698431365
transform 1 0 12544 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698431365
transform 1 0 16128 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_282
timestamp 1698431365
transform 1 0 16464 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_298
timestamp 1698431365
transform 1 0 17360 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_302
timestamp 1698431365
transform 1 0 17584 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_304
timestamp 1698431365
transform 1 0 17696 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_8
timestamp 1698431365
transform 1 0 1120 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_12
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698431365
transform 1 0 2240 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698431365
transform 1 0 2464 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698431365
transform 1 0 6664 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_115
timestamp 1698431365
transform 1 0 7112 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_119
timestamp 1698431365
transform 1 0 7336 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_121
timestamp 1698431365
transform 1 0 7448 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_154
timestamp 1698431365
transform 1 0 9296 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_158
timestamp 1698431365
transform 1 0 9520 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 10304 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 10416 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698431365
transform 1 0 10584 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698431365
transform 1 0 14168 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698431365
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698431365
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698431365
transform 1 0 18424 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_325
timestamp 1698431365
transform 1 0 18872 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_14
timestamp 1698431365
transform 1 0 1456 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_18
timestamp 1698431365
transform 1 0 1680 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_50
timestamp 1698431365
transform 1 0 3472 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698431365
transform 1 0 4704 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_104
timestamp 1698431365
transform 1 0 6496 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_120
timestamp 1698431365
transform 1 0 7392 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_128
timestamp 1698431365
transform 1 0 7840 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_135
timestamp 1698431365
transform 1 0 8232 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698431365
transform 1 0 8456 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_142
timestamp 1698431365
transform 1 0 8624 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698431365
transform 1 0 12208 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698431365
transform 1 0 12544 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698431365
transform 1 0 16128 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698431365
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698431365
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698431365
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698431365
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698431365
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698431365
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_107
timestamp 1698431365
transform 1 0 6664 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_139
timestamp 1698431365
transform 1 0 8456 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_141
timestamp 1698431365
transform 1 0 8568 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_152
timestamp 1698431365
transform 1 0 9184 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_162
timestamp 1698431365
transform 1 0 9744 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_170
timestamp 1698431365
transform 1 0 10192 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 10416 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_209
timestamp 1698431365
transform 1 0 12376 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698431365
transform 1 0 14168 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698431365
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_311
timestamp 1698431365
transform 1 0 18088 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 18424 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_8
timestamp 1698431365
transform 1 0 1120 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_12
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_44
timestamp 1698431365
transform 1 0 3136 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698431365
transform 1 0 4032 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698431365
transform 1 0 4480 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698431365
transform 1 0 4704 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_136
timestamp 1698431365
transform 1 0 8288 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_156
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_172
timestamp 1698431365
transform 1 0 10304 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698431365
transform 1 0 12320 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 12544 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_216
timestamp 1698431365
transform 1 0 12768 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_220
timestamp 1698431365
transform 1 0 12992 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_252
timestamp 1698431365
transform 1 0 14784 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_268
timestamp 1698431365
transform 1 0 15680 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 16128 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698431365
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698431365
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698431365
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_8
timestamp 1698431365
transform 1 0 1120 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_12
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698431365
transform 1 0 2240 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698431365
transform 1 0 2464 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_107
timestamp 1698431365
transform 1 0 6664 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_123
timestamp 1698431365
transform 1 0 7560 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698431365
transform 1 0 10360 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_177
timestamp 1698431365
transform 1 0 10584 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_185
timestamp 1698431365
transform 1 0 11032 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_198
timestamp 1698431365
transform 1 0 11760 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_230
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_238
timestamp 1698431365
transform 1 0 14000 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698431365
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698431365
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698431365
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698431365
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698431365
transform 1 0 2240 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698431365
transform 1 0 4032 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698431365
transform 1 0 4480 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698431365
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_104
timestamp 1698431365
transform 1 0 6496 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_120
timestamp 1698431365
transform 1 0 7392 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_128
timestamp 1698431365
transform 1 0 7840 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_132
timestamp 1698431365
transform 1 0 8064 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_148
timestamp 1698431365
transform 1 0 8960 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_156
timestamp 1698431365
transform 1 0 9408 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_159
timestamp 1698431365
transform 1 0 9576 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_191
timestamp 1698431365
transform 1 0 11368 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698431365
transform 1 0 12264 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698431365
transform 1 0 12544 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698431365
transform 1 0 16128 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698431365
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_314
timestamp 1698431365
transform 1 0 18256 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_318
timestamp 1698431365
transform 1 0 18480 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_321
timestamp 1698431365
transform 1 0 18648 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_8
timestamp 1698431365
transform 1 0 1120 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_12
timestamp 1698431365
transform 1 0 1344 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698431365
transform 1 0 2240 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698431365
transform 1 0 2464 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_107
timestamp 1698431365
transform 1 0 6664 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_123
timestamp 1698431365
transform 1 0 7560 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_159
timestamp 1698431365
transform 1 0 9576 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_209
timestamp 1698431365
transform 1 0 12376 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698431365
transform 1 0 14168 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698431365
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_311
timestamp 1698431365
transform 1 0 18088 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698431365
transform 1 0 18424 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_8
timestamp 1698431365
transform 1 0 1120 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_12
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_16
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_48
timestamp 1698431365
transform 1 0 3360 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_64
timestamp 1698431365
transform 1 0 4256 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 4480 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698431365
transform 1 0 4704 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 8288 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_142
timestamp 1698431365
transform 1 0 8624 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698431365
transform 1 0 12208 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698431365
transform 1 0 12544 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 16128 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_282
timestamp 1698431365
transform 1 0 16464 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_298
timestamp 1698431365
transform 1 0 17360 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_302
timestamp 1698431365
transform 1 0 17584 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_304
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_14
timestamp 1698431365
transform 1 0 1456 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_18
timestamp 1698431365
transform 1 0 1680 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698431365
transform 1 0 6664 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_123
timestamp 1698431365
transform 1 0 7560 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_127
timestamp 1698431365
transform 1 0 7784 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_129
timestamp 1698431365
transform 1 0 7896 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_162
timestamp 1698431365
transform 1 0 9744 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_170
timestamp 1698431365
transform 1 0 10192 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698431365
transform 1 0 10416 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698431365
transform 1 0 10584 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_190
timestamp 1698431365
transform 1 0 11312 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_222
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_238
timestamp 1698431365
transform 1 0 14000 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698431365
transform 1 0 14224 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 14336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698431365
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698431365
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698431365
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698431365
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_8
timestamp 1698431365
transform 1 0 1120 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_12
timestamp 1698431365
transform 1 0 1344 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_44
timestamp 1698431365
transform 1 0 3136 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698431365
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698431365
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698431365
transform 1 0 4704 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 8288 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_148
timestamp 1698431365
transform 1 0 8960 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_180
timestamp 1698431365
transform 1 0 10752 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_196
timestamp 1698431365
transform 1 0 11648 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_204
timestamp 1698431365
transform 1 0 12096 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_208
timestamp 1698431365
transform 1 0 12320 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698431365
transform 1 0 12544 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698431365
transform 1 0 16128 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698431365
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698431365
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698431365
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_8
timestamp 1698431365
transform 1 0 1120 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_12
timestamp 1698431365
transform 1 0 1344 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698431365
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698431365
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698431365
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698431365
transform 1 0 6664 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_123
timestamp 1698431365
transform 1 0 7560 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_127
timestamp 1698431365
transform 1 0 7784 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_129
timestamp 1698431365
transform 1 0 7896 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_162
timestamp 1698431365
transform 1 0 9744 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_170
timestamp 1698431365
transform 1 0 10192 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 10416 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_177
timestamp 1698431365
transform 1 0 10584 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698431365
transform 1 0 14168 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698431365
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698431365
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698431365
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_8
timestamp 1698431365
transform 1 0 1120 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_12
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_44
timestamp 1698431365
transform 1 0 3136 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698431365
transform 1 0 4032 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698431365
transform 1 0 4480 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698431365
transform 1 0 4704 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 8288 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_148
timestamp 1698431365
transform 1 0 8960 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_180
timestamp 1698431365
transform 1 0 10752 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_196
timestamp 1698431365
transform 1 0 11648 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_204
timestamp 1698431365
transform 1 0 12096 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698431365
transform 1 0 12320 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698431365
transform 1 0 12544 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698431365
transform 1 0 16128 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_282
timestamp 1698431365
transform 1 0 16464 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_298
timestamp 1698431365
transform 1 0 17360 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_302
timestamp 1698431365
transform 1 0 17584 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_304
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_8
timestamp 1698431365
transform 1 0 1120 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_12
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698431365
transform 1 0 2240 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698431365
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698431365
transform 1 0 6664 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 10248 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698431365
transform 1 0 10584 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698431365
transform 1 0 14168 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698431365
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698431365
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_317
timestamp 1698431365
transform 1 0 18424 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_325
timestamp 1698431365
transform 1 0 18872 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_329
timestamp 1698431365
transform 1 0 19096 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_28
timestamp 1698431365
transform 1 0 2240 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_32
timestamp 1698431365
transform 1 0 2464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_64
timestamp 1698431365
transform 1 0 4256 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 4480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 4704 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 8288 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_142
timestamp 1698431365
transform 1 0 8624 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 12208 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698431365
transform 1 0 12544 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 16128 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698431365
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_314
timestamp 1698431365
transform 1 0 18256 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_330
timestamp 1698431365
transform 1 0 19152 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698431365
transform 1 0 6664 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 10248 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698431365
transform 1 0 10584 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698431365
transform 1 0 14168 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698431365
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_317
timestamp 1698431365
transform 1 0 18424 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_325
timestamp 1698431365
transform 1 0 18872 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_329
timestamp 1698431365
transform 1 0 19096 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698431365
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698431365
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698431365
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698431365
transform 1 0 8624 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 12208 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698431365
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698431365
transform 1 0 16464 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_314
timestamp 1698431365
transform 1 0 18256 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_330
timestamp 1698431365
transform 1 0 19152 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698431365
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698431365
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698431365
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698431365
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_317
timestamp 1698431365
transform 1 0 18424 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_325
timestamp 1698431365
transform 1 0 18872 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_329
timestamp 1698431365
transform 1 0 19096 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698431365
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698431365
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698431365
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_282
timestamp 1698431365
transform 1 0 16464 0 -1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_314
timestamp 1698431365
transform 1 0 18256 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_330
timestamp 1698431365
transform 1 0 19152 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698431365
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698431365
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_317
timestamp 1698431365
transform 1 0 18424 0 1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_325
timestamp 1698431365
transform 1 0 18872 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_329
timestamp 1698431365
transform 1 0 19096 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_282
timestamp 1698431365
transform 1 0 16464 0 -1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_314
timestamp 1698431365
transform 1 0 18256 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_330
timestamp 1698431365
transform 1 0 19152 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_317
timestamp 1698431365
transform 1 0 18424 0 1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_325
timestamp 1698431365
transform 1 0 18872 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_329
timestamp 1698431365
transform 1 0 19096 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_282
timestamp 1698431365
transform 1 0 16464 0 -1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_314
timestamp 1698431365
transform 1 0 18256 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_330
timestamp 1698431365
transform 1 0 19152 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_317
timestamp 1698431365
transform 1 0 18424 0 1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_325
timestamp 1698431365
transform 1 0 18872 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_329
timestamp 1698431365
transform 1 0 19096 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_282
timestamp 1698431365
transform 1 0 16464 0 -1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_314
timestamp 1698431365
transform 1 0 18256 0 -1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_330
timestamp 1698431365
transform 1 0 19152 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_107
timestamp 1698431365
transform 1 0 6664 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_139
timestamp 1698431365
transform 1 0 8456 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_145
timestamp 1698431365
transform 1 0 8792 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_151
timestamp 1698431365
transform 1 0 9128 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_157
timestamp 1698431365
transform 1 0 9464 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_163
timestamp 1698431365
transform 1 0 9800 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_169
timestamp 1698431365
transform 1 0 10136 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 10360 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_317
timestamp 1698431365
transform 1 0 18424 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_325
timestamp 1698431365
transform 1 0 18872 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_329
timestamp 1698431365
transform 1 0 19096 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_72
timestamp 1698431365
transform 1 0 4704 0 -1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_104
timestamp 1698431365
transform 1 0 6496 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_120
timestamp 1698431365
transform 1 0 7392 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_123
timestamp 1698431365
transform 1 0 7560 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 8456 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_142
timestamp 1698431365
transform 1 0 8624 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_144
timestamp 1698431365
transform 1 0 8736 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_175
timestamp 1698431365
transform 1 0 10472 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_181
timestamp 1698431365
transform 1 0 10808 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_187
timestamp 1698431365
transform 1 0 11144 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_203
timestamp 1698431365
transform 1 0 12040 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_207
timestamp 1698431365
transform 1 0 12264 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_209
timestamp 1698431365
transform 1 0 12376 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_282
timestamp 1698431365
transform 1 0 16464 0 -1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_314
timestamp 1698431365
transform 1 0 18256 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_330
timestamp 1698431365
transform 1 0 19152 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_36
timestamp 1698431365
transform 1 0 2688 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_70
timestamp 1698431365
transform 1 0 4592 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_104
timestamp 1698431365
transform 1 0 6496 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_108
timestamp 1698431365
transform 1 0 6720 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_138
timestamp 1698431365
transform 1 0 8400 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_165
timestamp 1698431365
transform 1 0 9912 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_167
timestamp 1698431365
transform 1 0 10024 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_172
timestamp 1698431365
transform 1 0 10304 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 10416 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_193
timestamp 1698431365
transform 1 0 11480 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_201
timestamp 1698431365
transform 1 0 11928 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_203
timestamp 1698431365
transform 1 0 12040 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_206
timestamp 1698431365
transform 1 0 12208 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_240
timestamp 1698431365
transform 1 0 14112 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_274
timestamp 1698431365
transform 1 0 16016 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_308
timestamp 1698431365
transform 1 0 17920 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_324
timestamp 1698431365
transform 1 0 18816 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_328
timestamp 1698431365
transform 1 0 19040 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_330
timestamp 1698431365
transform 1 0 19152 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19208 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 784 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 9800 0 -1 18032
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 18872 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 19208 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 19208 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 19208 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 7952 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 11816 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 10808 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform -1 0 8456 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 18872 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 1120 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 9464 0 -1 18032
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 784 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 8792 0 -1 18032
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 19208 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform -1 0 19208 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 10808 0 1 18032
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 10136 0 -1 18032
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform 1 0 784 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 7112 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform -1 0 19208 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform 1 0 8848 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform 1 0 7448 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform 1 0 784 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 784 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 784 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 784 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 19208 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 19208 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform -1 0 11480 0 1 18032
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 10808 0 1 18032
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform -1 0 19208 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 1120 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform -1 0 9520 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform -1 0 9856 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform 1 0 7784 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 784 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform 1 0 7784 0 -1 18032
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform 1 0 784 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform 1 0 8120 0 -1 18032
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698431365
transform 1 0 8512 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698431365
transform -1 0 11480 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1698431365
transform -1 0 11144 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698431365
transform 1 0 6776 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698431365
transform 1 0 784 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698431365
transform -1 0 10136 0 -1 18032
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input49
timestamp 1698431365
transform 1 0 784 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1698431365
transform -1 0 10192 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output51 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17752 0 -1 7056
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output52
timestamp 1698431365
transform -1 0 2240 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output53
timestamp 1698431365
transform -1 0 8288 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output54
timestamp 1698431365
transform 1 0 17752 0 -1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output55
timestamp 1698431365
transform 1 0 17752 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output56
timestamp 1698431365
transform 1 0 17752 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output57
timestamp 1698431365
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output58
timestamp 1698431365
transform 1 0 12544 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output59
timestamp 1698431365
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output60
timestamp 1698431365
transform -1 0 7952 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output61
timestamp 1698431365
transform -1 0 2240 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output62
timestamp 1698431365
transform 1 0 8456 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_43 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 19320 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_44
timestamp 1698431365
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 19320 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_45
timestamp 1698431365
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 19320 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_46
timestamp 1698431365
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 19320 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_47
timestamp 1698431365
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 19320 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_48
timestamp 1698431365
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 19320 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_49
timestamp 1698431365
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 19320 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_50
timestamp 1698431365
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 19320 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_51
timestamp 1698431365
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 19320 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_52
timestamp 1698431365
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 19320 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_53
timestamp 1698431365
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 19320 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_54
timestamp 1698431365
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 19320 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_55
timestamp 1698431365
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 19320 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_56
timestamp 1698431365
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 19320 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_57
timestamp 1698431365
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 19320 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_58
timestamp 1698431365
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 19320 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_59
timestamp 1698431365
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 19320 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_60
timestamp 1698431365
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 19320 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_61
timestamp 1698431365
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 19320 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_62
timestamp 1698431365
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 19320 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_63
timestamp 1698431365
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 19320 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_64
timestamp 1698431365
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 19320 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_65
timestamp 1698431365
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 19320 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_66
timestamp 1698431365
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 19320 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_67
timestamp 1698431365
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 19320 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_68
timestamp 1698431365
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 19320 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_69
timestamp 1698431365
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 19320 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_70
timestamp 1698431365
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 19320 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_71
timestamp 1698431365
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 19320 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_72
timestamp 1698431365
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 19320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_73
timestamp 1698431365
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 19320 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_74
timestamp 1698431365
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 19320 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_75
timestamp 1698431365
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 19320 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_76
timestamp 1698431365
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 19320 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_77
timestamp 1698431365
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 19320 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_78
timestamp 1698431365
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 19320 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_79
timestamp 1698431365
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 19320 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_80
timestamp 1698431365
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 19320 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_81
timestamp 1698431365
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 19320 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_82
timestamp 1698431365
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 19320 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_83
timestamp 1698431365
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 19320 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_84
timestamp 1698431365
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 19320 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_85
timestamp 1698431365
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 19320 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_86 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_87
timestamp 1698431365
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_88
timestamp 1698431365
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_89
timestamp 1698431365
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90
timestamp 1698431365
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698431365
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698431365
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698431365
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698431365
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_95
timestamp 1698431365
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_96
timestamp 1698431365
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_97
timestamp 1698431365
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_98
timestamp 1698431365
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_99
timestamp 1698431365
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_100
timestamp 1698431365
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_101
timestamp 1698431365
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_102
timestamp 1698431365
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_103
timestamp 1698431365
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_104
timestamp 1698431365
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_105
timestamp 1698431365
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_106
timestamp 1698431365
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_107
timestamp 1698431365
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_108
timestamp 1698431365
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_109
timestamp 1698431365
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_110
timestamp 1698431365
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_111
timestamp 1698431365
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_112
timestamp 1698431365
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_113
timestamp 1698431365
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_114
timestamp 1698431365
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_115
timestamp 1698431365
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_116
timestamp 1698431365
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_117
timestamp 1698431365
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_118
timestamp 1698431365
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_119
timestamp 1698431365
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_120
timestamp 1698431365
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_121
timestamp 1698431365
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_122
timestamp 1698431365
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_123
timestamp 1698431365
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_124
timestamp 1698431365
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_125
timestamp 1698431365
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_126
timestamp 1698431365
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_127
timestamp 1698431365
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_128
timestamp 1698431365
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_129
timestamp 1698431365
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_130
timestamp 1698431365
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_131
timestamp 1698431365
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_132
timestamp 1698431365
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_133
timestamp 1698431365
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_134
timestamp 1698431365
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_135
timestamp 1698431365
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_136
timestamp 1698431365
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_137
timestamp 1698431365
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_138
timestamp 1698431365
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_139
timestamp 1698431365
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_140
timestamp 1698431365
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_141
timestamp 1698431365
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_142
timestamp 1698431365
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_143
timestamp 1698431365
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_144
timestamp 1698431365
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_145
timestamp 1698431365
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_146
timestamp 1698431365
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_147
timestamp 1698431365
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_148
timestamp 1698431365
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_149
timestamp 1698431365
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_150
timestamp 1698431365
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_151
timestamp 1698431365
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_152
timestamp 1698431365
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_153
timestamp 1698431365
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_154
timestamp 1698431365
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_155
timestamp 1698431365
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_156
timestamp 1698431365
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_157
timestamp 1698431365
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_158
timestamp 1698431365
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_159
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_160
timestamp 1698431365
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_161
timestamp 1698431365
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_162
timestamp 1698431365
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_163
timestamp 1698431365
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_164
timestamp 1698431365
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_165
timestamp 1698431365
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_166
timestamp 1698431365
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_167
timestamp 1698431365
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_168
timestamp 1698431365
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_169
timestamp 1698431365
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_170
timestamp 1698431365
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_171
timestamp 1698431365
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_172
timestamp 1698431365
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_173
timestamp 1698431365
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_174
timestamp 1698431365
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_175
timestamp 1698431365
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_176
timestamp 1698431365
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_177
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_178
timestamp 1698431365
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_179
timestamp 1698431365
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_180
timestamp 1698431365
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_181
timestamp 1698431365
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_182
timestamp 1698431365
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_183
timestamp 1698431365
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_184
timestamp 1698431365
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_185
timestamp 1698431365
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_186
timestamp 1698431365
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_187
timestamp 1698431365
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_188
timestamp 1698431365
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_189
timestamp 1698431365
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_190
timestamp 1698431365
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_191
timestamp 1698431365
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_192
timestamp 1698431365
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_193
timestamp 1698431365
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_194
timestamp 1698431365
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_195
timestamp 1698431365
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_196
timestamp 1698431365
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_197
timestamp 1698431365
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_198
timestamp 1698431365
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_199
timestamp 1698431365
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_200
timestamp 1698431365
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_201
timestamp 1698431365
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_202
timestamp 1698431365
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_203
timestamp 1698431365
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_204
timestamp 1698431365
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_205
timestamp 1698431365
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_206
timestamp 1698431365
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_207
timestamp 1698431365
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_208
timestamp 1698431365
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_209
timestamp 1698431365
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_210
timestamp 1698431365
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_211
timestamp 1698431365
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_212
timestamp 1698431365
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_213
timestamp 1698431365
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_214
timestamp 1698431365
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_215
timestamp 1698431365
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_216
timestamp 1698431365
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_217
timestamp 1698431365
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_218
timestamp 1698431365
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_219
timestamp 1698431365
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_220
timestamp 1698431365
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_221
timestamp 1698431365
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_222
timestamp 1698431365
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_223
timestamp 1698431365
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_224
timestamp 1698431365
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_225
timestamp 1698431365
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_226
timestamp 1698431365
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_227
timestamp 1698431365
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_228
timestamp 1698431365
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_229
timestamp 1698431365
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_230
timestamp 1698431365
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_231
timestamp 1698431365
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_232
timestamp 1698431365
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_233
timestamp 1698431365
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_234
timestamp 1698431365
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_235
timestamp 1698431365
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_236
timestamp 1698431365
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_237
timestamp 1698431365
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_238
timestamp 1698431365
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_239
timestamp 1698431365
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_240
timestamp 1698431365
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_241
timestamp 1698431365
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_242
timestamp 1698431365
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_243
timestamp 1698431365
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_244
timestamp 1698431365
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_245
timestamp 1698431365
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_246
timestamp 1698431365
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_247
timestamp 1698431365
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_248
timestamp 1698431365
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_249
timestamp 1698431365
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_250
timestamp 1698431365
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_251
timestamp 1698431365
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_252
timestamp 1698431365
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_253
timestamp 1698431365
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_254
timestamp 1698431365
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_255
timestamp 1698431365
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_256
timestamp 1698431365
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_257
timestamp 1698431365
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_258
timestamp 1698431365
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_259
timestamp 1698431365
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_260
timestamp 1698431365
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_261
timestamp 1698431365
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_262
timestamp 1698431365
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_263
timestamp 1698431365
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_264
timestamp 1698431365
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_265
timestamp 1698431365
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_266
timestamp 1698431365
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_267
timestamp 1698431365
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_268
timestamp 1698431365
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_269
timestamp 1698431365
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_270
timestamp 1698431365
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_271
timestamp 1698431365
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_272
timestamp 1698431365
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_273
timestamp 1698431365
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_274
timestamp 1698431365
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_275
timestamp 1698431365
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_276
timestamp 1698431365
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_277
timestamp 1698431365
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_278
timestamp 1698431365
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_279
timestamp 1698431365
transform 1 0 2576 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_280
timestamp 1698431365
transform 1 0 4480 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_281
timestamp 1698431365
transform 1 0 6384 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_282
timestamp 1698431365
transform 1 0 8288 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_283
timestamp 1698431365
transform 1 0 10192 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698431365
transform 1 0 12096 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698431365
transform 1 0 14000 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698431365
transform 1 0 15904 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698431365
transform 1 0 17808 0 1 18032
box -43 -43 155 435
<< labels >>
flabel metal3 s 19600 7056 20000 7112 0 FreeSans 224 0 0 0 out[0]
port 0 nsew signal tristate
flabel metal3 s 0 9744 400 9800 0 FreeSans 224 0 0 0 out[10]
port 1 nsew signal tristate
flabel metal2 s 7392 19600 7448 20000 0 FreeSans 224 90 0 0 out[11]
port 2 nsew signal tristate
flabel metal3 s 19600 7728 20000 7784 0 FreeSans 224 0 0 0 out[1]
port 3 nsew signal tristate
flabel metal3 s 19600 12096 20000 12152 0 FreeSans 224 0 0 0 out[2]
port 4 nsew signal tristate
flabel metal3 s 19600 10752 20000 10808 0 FreeSans 224 0 0 0 out[3]
port 5 nsew signal tristate
flabel metal3 s 0 8400 400 8456 0 FreeSans 224 0 0 0 out[4]
port 6 nsew signal tristate
flabel metal2 s 12096 0 12152 400 0 FreeSans 224 90 0 0 out[5]
port 7 nsew signal tristate
flabel metal2 s 11760 0 11816 400 0 FreeSans 224 90 0 0 out[6]
port 8 nsew signal tristate
flabel metal2 s 6384 0 6440 400 0 FreeSans 224 90 0 0 out[7]
port 9 nsew signal tristate
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 out[8]
port 10 nsew signal tristate
flabel metal2 s 8400 19600 8456 20000 0 FreeSans 224 90 0 0 out[9]
port 11 nsew signal tristate
flabel metal3 s 19600 9408 20000 9464 0 FreeSans 224 0 0 0 proj_out[0]
port 12 nsew signal input
flabel metal3 s 0 9072 400 9128 0 FreeSans 224 0 0 0 proj_out[10]
port 13 nsew signal input
flabel metal2 s 9408 19600 9464 20000 0 FreeSans 224 90 0 0 proj_out[11]
port 14 nsew signal input
flabel metal3 s 19600 10080 20000 10136 0 FreeSans 224 0 0 0 proj_out[12]
port 15 nsew signal input
flabel metal3 s 19600 8736 20000 8792 0 FreeSans 224 0 0 0 proj_out[13]
port 16 nsew signal input
flabel metal3 s 19600 11088 20000 11144 0 FreeSans 224 0 0 0 proj_out[14]
port 17 nsew signal input
flabel metal3 s 19600 11760 20000 11816 0 FreeSans 224 0 0 0 proj_out[15]
port 18 nsew signal input
flabel metal2 s 8400 0 8456 400 0 FreeSans 224 90 0 0 proj_out[16]
port 19 nsew signal input
flabel metal2 s 11424 0 11480 400 0 FreeSans 224 90 0 0 proj_out[17]
port 20 nsew signal input
flabel metal2 s 10416 0 10472 400 0 FreeSans 224 90 0 0 proj_out[18]
port 21 nsew signal input
flabel metal2 s 8064 0 8120 400 0 FreeSans 224 90 0 0 proj_out[19]
port 22 nsew signal input
flabel metal3 s 19600 8400 20000 8456 0 FreeSans 224 0 0 0 proj_out[1]
port 23 nsew signal input
flabel metal3 s 0 10752 400 10808 0 FreeSans 224 0 0 0 proj_out[20]
port 24 nsew signal input
flabel metal2 s 9072 19600 9128 20000 0 FreeSans 224 90 0 0 proj_out[21]
port 25 nsew signal input
flabel metal3 s 0 10080 400 10136 0 FreeSans 224 0 0 0 proj_out[22]
port 26 nsew signal input
flabel metal2 s 8736 19600 8792 20000 0 FreeSans 224 90 0 0 proj_out[23]
port 27 nsew signal input
flabel metal3 s 19600 9744 20000 9800 0 FreeSans 224 0 0 0 proj_out[24]
port 28 nsew signal input
flabel metal3 s 19600 9072 20000 9128 0 FreeSans 224 0 0 0 proj_out[25]
port 29 nsew signal input
flabel metal2 s 10416 19600 10472 20000 0 FreeSans 224 90 0 0 proj_out[26]
port 30 nsew signal input
flabel metal2 s 10080 19600 10136 20000 0 FreeSans 224 90 0 0 proj_out[27]
port 31 nsew signal input
flabel metal3 s 0 7728 400 7784 0 FreeSans 224 0 0 0 proj_out[28]
port 32 nsew signal input
flabel metal2 s 7056 0 7112 400 0 FreeSans 224 90 0 0 proj_out[29]
port 33 nsew signal input
flabel metal3 s 19600 11424 20000 11480 0 FreeSans 224 0 0 0 proj_out[2]
port 34 nsew signal input
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 proj_out[30]
port 35 nsew signal input
flabel metal2 s 7392 0 7448 400 0 FreeSans 224 90 0 0 proj_out[31]
port 36 nsew signal input
flabel metal3 s 0 11088 400 11144 0 FreeSans 224 0 0 0 proj_out[32]
port 37 nsew signal input
flabel metal3 s 0 12096 400 12152 0 FreeSans 224 0 0 0 proj_out[33]
port 38 nsew signal input
flabel metal3 s 0 12432 400 12488 0 FreeSans 224 0 0 0 proj_out[34]
port 39 nsew signal input
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 proj_out[35]
port 40 nsew signal input
flabel metal3 s 19600 7392 20000 7448 0 FreeSans 224 0 0 0 proj_out[36]
port 41 nsew signal input
flabel metal3 s 19600 8064 20000 8120 0 FreeSans 224 0 0 0 proj_out[37]
port 42 nsew signal input
flabel metal2 s 11088 19600 11144 20000 0 FreeSans 224 90 0 0 proj_out[38]
port 43 nsew signal input
flabel metal2 s 10752 19600 10808 20000 0 FreeSans 224 90 0 0 proj_out[39]
port 44 nsew signal input
flabel metal3 s 19600 10416 20000 10472 0 FreeSans 224 0 0 0 proj_out[3]
port 45 nsew signal input
flabel metal3 s 0 8064 400 8120 0 FreeSans 224 0 0 0 proj_out[40]
port 46 nsew signal input
flabel metal2 s 9408 0 9464 400 0 FreeSans 224 90 0 0 proj_out[41]
port 47 nsew signal input
flabel metal2 s 9744 0 9800 400 0 FreeSans 224 90 0 0 proj_out[42]
port 48 nsew signal input
flabel metal2 s 7728 0 7784 400 0 FreeSans 224 90 0 0 proj_out[43]
port 49 nsew signal input
flabel metal3 s 0 10416 400 10472 0 FreeSans 224 0 0 0 proj_out[44]
port 50 nsew signal input
flabel metal2 s 7728 19600 7784 20000 0 FreeSans 224 90 0 0 proj_out[45]
port 51 nsew signal input
flabel metal3 s 0 9408 400 9464 0 FreeSans 224 0 0 0 proj_out[46]
port 52 nsew signal input
flabel metal2 s 8064 19600 8120 20000 0 FreeSans 224 90 0 0 proj_out[47]
port 53 nsew signal input
flabel metal2 s 8736 0 8792 400 0 FreeSans 224 90 0 0 proj_out[4]
port 54 nsew signal input
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 proj_out[5]
port 55 nsew signal input
flabel metal2 s 10752 0 10808 400 0 FreeSans 224 90 0 0 proj_out[6]
port 56 nsew signal input
flabel metal2 s 6720 0 6776 400 0 FreeSans 224 90 0 0 proj_out[7]
port 57 nsew signal input
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 proj_out[8]
port 58 nsew signal input
flabel metal2 s 9744 19600 9800 20000 0 FreeSans 224 90 0 0 proj_out[9]
port 59 nsew signal input
flabel metal3 s 0 8736 400 8792 0 FreeSans 224 0 0 0 sel[0]
port 60 nsew signal input
flabel metal2 s 10080 0 10136 400 0 FreeSans 224 90 0 0 sel[1]
port 61 nsew signal input
flabel metal4 s 2923 1538 3083 18454 0 FreeSans 640 90 0 0 vdd
port 62 nsew power bidirectional
flabel metal4 s 7585 1538 7745 18454 0 FreeSans 640 90 0 0 vdd
port 62 nsew power bidirectional
flabel metal4 s 12247 1538 12407 18454 0 FreeSans 640 90 0 0 vdd
port 62 nsew power bidirectional
flabel metal4 s 16909 1538 17069 18454 0 FreeSans 640 90 0 0 vdd
port 62 nsew power bidirectional
flabel metal4 s 5254 1538 5414 18454 0 FreeSans 640 90 0 0 vss
port 63 nsew ground bidirectional
flabel metal4 s 9916 1538 10076 18454 0 FreeSans 640 90 0 0 vss
port 63 nsew ground bidirectional
flabel metal4 s 14578 1538 14738 18454 0 FreeSans 640 90 0 0 vss
port 63 nsew ground bidirectional
flabel metal4 s 19240 1538 19400 18454 0 FreeSans 640 90 0 0 vss
port 63 nsew ground bidirectional
rlabel metal1 9996 18424 9996 18424 0 vdd
rlabel via1 10036 18032 10036 18032 0 vss
rlabel metal2 10836 10584 10836 10584 0 _00_
rlabel metal2 11368 10388 11368 10388 0 _01_
rlabel metal2 11116 9408 11116 9408 0 _02_
rlabel metal2 11340 8708 11340 8708 0 _03_
rlabel metal2 11004 10976 11004 10976 0 _04_
rlabel metal2 11200 10332 11200 10332 0 _05_
rlabel metal2 9324 7672 9324 7672 0 _06_
rlabel metal3 8008 7980 8008 7980 0 _07_
rlabel metal2 8092 8204 8092 8204 0 _08_
rlabel metal3 9660 7924 9660 7924 0 _09_
rlabel metal2 9688 7756 9688 7756 0 _10_
rlabel metal2 8036 7756 8036 7756 0 _11_
rlabel metal2 8204 11564 8204 11564 0 _12_
rlabel metal2 8876 11564 8876 11564 0 _13_
rlabel metal2 8372 10136 8372 10136 0 _14_
rlabel metal2 8820 11704 8820 11704 0 _15_
rlabel metal3 8596 9548 8596 9548 0 _16_
rlabel metal2 8540 11312 8540 11312 0 _17_
rlabel metal2 12180 9352 12180 9352 0 net1
rlabel metal2 10304 7644 10304 7644 0 net10
rlabel metal2 7308 4956 7308 4956 0 net11
rlabel metal2 12236 8848 12236 8848 0 net12
rlabel metal2 8876 10724 8876 10724 0 net13
rlabel metal2 9212 17766 9212 17766 0 net14
rlabel metal3 4956 10276 4956 10276 0 net15
rlabel metal2 9156 11466 9156 11466 0 net16
rlabel metal3 11648 9156 11648 9156 0 net17
rlabel metal3 13314 8764 13314 8764 0 net18
rlabel metal2 10500 11298 10500 11298 0 net19
rlabel metal2 1036 9240 1036 9240 0 net2
rlabel metal2 10640 10444 10640 10444 0 net20
rlabel metal3 2618 7924 2618 7924 0 net21
rlabel metal2 7364 4732 7364 4732 0 net22
rlabel metal2 12068 11200 12068 11200 0 net23
rlabel metal2 9128 7588 9128 7588 0 net24
rlabel metal2 7700 2464 7700 2464 0 net25
rlabel metal2 1036 11144 1036 11144 0 net26
rlabel metal2 8036 12208 8036 12208 0 net27
rlabel metal2 1092 12628 1092 12628 0 net28
rlabel metal2 8036 11536 8036 11536 0 net29
rlabel metal2 9576 13524 9576 13524 0 net3
rlabel metal2 12964 9044 12964 9044 0 net30
rlabel metal2 11116 8596 11116 8596 0 net31
rlabel metal3 11060 10780 11060 10780 0 net32
rlabel metal2 11088 10388 11088 10388 0 net33
rlabel metal2 12236 10360 12236 10360 0 net34
rlabel metal2 1372 8260 1372 8260 0 net35
rlabel metal2 9212 6580 9212 6580 0 net36
rlabel metal2 9604 4676 9604 4676 0 net37
rlabel metal2 8036 4956 8036 4956 0 net38
rlabel metal2 8260 10612 8260 10612 0 net39
rlabel metal2 18620 10178 18620 10178 0 net4
rlabel metal3 8232 14980 8232 14980 0 net40
rlabel metal3 8260 9548 8260 9548 0 net41
rlabel metal2 8456 11172 8456 11172 0 net42
rlabel metal2 9044 8036 9044 8036 0 net43
rlabel metal2 11228 3808 11228 3808 0 net44
rlabel metal2 10724 7602 10724 7602 0 net45
rlabel metal2 7028 3234 7028 3234 0 net46
rlabel metal2 1092 10976 1092 10976 0 net47
rlabel metal2 9520 13468 9520 13468 0 net48
rlabel metal2 1036 8400 1036 8400 0 net49
rlabel metal2 18956 8792 18956 8792 0 net5
rlabel metal2 9520 8820 9520 8820 0 net50
rlabel metal2 11452 9604 11452 9604 0 net51
rlabel metal3 8708 10024 8708 10024 0 net52
rlabel metal2 8260 18228 8260 18228 0 net53
rlabel metal2 11676 9408 11676 9408 0 net54
rlabel metal2 11228 11732 11228 11732 0 net55
rlabel metal2 17836 10920 17836 10920 0 net56
rlabel metal2 2156 8484 2156 8484 0 net57
rlabel metal3 11424 7924 11424 7924 0 net58
rlabel metal2 9884 7840 9884 7840 0 net59
rlabel metal3 13790 10780 13790 10780 0 net6
rlabel metal3 7980 1764 7980 1764 0 net60
rlabel metal2 2156 13104 2156 13104 0 net61
rlabel metal2 8708 11956 8708 11956 0 net62
rlabel metal2 18900 11116 18900 11116 0 net7
rlabel metal2 8540 8036 8540 8036 0 net8
rlabel metal2 11564 1666 11564 1666 0 net9
rlabel metal2 19012 6888 19012 6888 0 out[0]
rlabel metal3 679 9772 679 9772 0 out[10]
rlabel metal2 7420 18949 7420 18949 0 out[11]
rlabel metal2 19012 7672 19012 7672 0 out[1]
rlabel metal2 19012 12180 19012 12180 0 out[2]
rlabel metal2 19012 10752 19012 10752 0 out[3]
rlabel metal3 679 8428 679 8428 0 out[4]
rlabel metal3 12628 2044 12628 2044 0 out[5]
rlabel metal3 12292 1820 12292 1820 0 out[6]
rlabel metal2 6412 1099 6412 1099 0 out[7]
rlabel metal3 679 12796 679 12796 0 out[8]
rlabel metal2 8428 18977 8428 18977 0 out[9]
rlabel metal2 19124 9520 19124 9520 0 proj_out[0]
rlabel metal2 868 9156 868 9156 0 proj_out[10]
rlabel metal2 9660 18060 9660 18060 0 proj_out[11]
rlabel metal3 19229 10108 19229 10108 0 proj_out[12]
rlabel metal3 19369 8764 19369 8764 0 proj_out[13]
rlabel metal3 19369 11116 19369 11116 0 proj_out[14]
rlabel metal2 19124 11872 19124 11872 0 proj_out[15]
rlabel metal2 8428 1029 8428 1029 0 proj_out[16]
rlabel metal2 11564 1260 11564 1260 0 proj_out[17]
rlabel metal2 10556 1260 10556 1260 0 proj_out[18]
rlabel metal2 8204 1540 8204 1540 0 proj_out[19]
rlabel metal3 19201 8428 19201 8428 0 proj_out[1]
rlabel metal2 1204 10948 1204 10948 0 proj_out[20]
rlabel metal2 9324 18060 9324 18060 0 proj_out[21]
rlabel metal2 868 10220 868 10220 0 proj_out[22]
rlabel metal2 8820 17892 8820 17892 0 proj_out[23]
rlabel metal2 19124 9884 19124 9884 0 proj_out[24]
rlabel metal2 19124 9156 19124 9156 0 proj_out[25]
rlabel metal2 10164 18480 10164 18480 0 proj_out[26]
rlabel metal2 10164 17892 10164 17892 0 proj_out[27]
rlabel metal3 651 7756 651 7756 0 proj_out[28]
rlabel metal2 7196 1960 7196 1960 0 proj_out[29]
rlabel metal2 19124 11508 19124 11508 0 proj_out[2]
rlabel metal2 9044 1260 9044 1260 0 proj_out[30]
rlabel metal2 7532 1848 7532 1848 0 proj_out[31]
rlabel metal3 623 11116 623 11116 0 proj_out[32]
rlabel metal2 868 12236 868 12236 0 proj_out[33]
rlabel metal2 868 12572 868 12572 0 proj_out[34]
rlabel metal2 868 11844 868 11844 0 proj_out[35]
rlabel metal2 19124 7336 19124 7336 0 proj_out[36]
rlabel metal3 19397 8092 19397 8092 0 proj_out[37]
rlabel metal2 11228 18228 11228 18228 0 proj_out[38]
rlabel metal2 10836 18228 10836 18228 0 proj_out[39]
rlabel metal2 19124 10416 19124 10416 0 proj_out[3]
rlabel metal2 1204 8260 1204 8260 0 proj_out[40]
rlabel metal2 9492 2100 9492 2100 0 proj_out[41]
rlabel metal2 9828 2100 9828 2100 0 proj_out[42]
rlabel metal2 7756 1029 7756 1029 0 proj_out[43]
rlabel metal2 868 10612 868 10612 0 proj_out[44]
rlabel metal2 7868 18200 7868 18200 0 proj_out[45]
rlabel metal2 868 9492 868 9492 0 proj_out[46]
rlabel metal2 8148 17892 8148 17892 0 proj_out[47]
rlabel metal2 8708 1260 8708 1260 0 proj_out[4]
rlabel metal2 11228 1260 11228 1260 0 proj_out[5]
rlabel metal2 11004 1932 11004 1932 0 proj_out[6]
rlabel metal2 6860 1792 6860 1792 0 proj_out[7]
rlabel metal2 868 11508 868 11508 0 proj_out[8]
rlabel metal2 9996 17808 9996 17808 0 proj_out[9]
rlabel metal2 868 8652 868 8652 0 sel[0]
rlabel metal2 10136 2100 10136 2100 0 sel[1]
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
