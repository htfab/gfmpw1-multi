magic
tech gf180mcuD
magscale 1 10
timestamp 1702441479
<< metal1 >>
rect 1344 36874 38640 36908
rect 1344 36822 5876 36874
rect 5928 36822 5980 36874
rect 6032 36822 6084 36874
rect 6136 36822 15200 36874
rect 15252 36822 15304 36874
rect 15356 36822 15408 36874
rect 15460 36822 24524 36874
rect 24576 36822 24628 36874
rect 24680 36822 24732 36874
rect 24784 36822 33848 36874
rect 33900 36822 33952 36874
rect 34004 36822 34056 36874
rect 34108 36822 38640 36874
rect 1344 36788 38640 36822
rect 17166 36706 17218 36718
rect 17166 36642 17218 36654
rect 22094 36706 22146 36718
rect 22094 36642 22146 36654
rect 10222 36594 10274 36606
rect 10222 36530 10274 36542
rect 28478 36594 28530 36606
rect 28478 36530 28530 36542
rect 19854 36482 19906 36494
rect 26238 36482 26290 36494
rect 10994 36430 11006 36482
rect 11058 36430 11070 36482
rect 11666 36430 11678 36482
rect 11730 36430 11742 36482
rect 12338 36430 12350 36482
rect 12402 36430 12414 36482
rect 13458 36430 13470 36482
rect 13522 36430 13534 36482
rect 14130 36430 14142 36482
rect 14194 36430 14206 36482
rect 14802 36430 14814 36482
rect 14866 36430 14878 36482
rect 15474 36430 15486 36482
rect 15538 36430 15550 36482
rect 16146 36430 16158 36482
rect 16210 36430 16222 36482
rect 19170 36430 19182 36482
rect 19234 36430 19246 36482
rect 21074 36430 21086 36482
rect 21138 36430 21150 36482
rect 24770 36430 24782 36482
rect 24834 36430 24846 36482
rect 25442 36430 25454 36482
rect 25506 36430 25518 36482
rect 26786 36430 26798 36482
rect 26850 36430 26862 36482
rect 27458 36430 27470 36482
rect 27522 36430 27534 36482
rect 19854 36418 19906 36430
rect 26238 36418 26290 36430
rect 10670 36370 10722 36382
rect 10670 36306 10722 36318
rect 12574 36258 12626 36270
rect 14366 36258 14418 36270
rect 11218 36206 11230 36258
rect 11282 36206 11294 36258
rect 11890 36206 11902 36258
rect 11954 36206 11966 36258
rect 13682 36206 13694 36258
rect 13746 36206 13758 36258
rect 12574 36194 12626 36206
rect 14366 36194 14418 36206
rect 15038 36258 15090 36270
rect 15038 36194 15090 36206
rect 15710 36258 15762 36270
rect 20190 36258 20242 36270
rect 16370 36206 16382 36258
rect 16434 36206 16446 36258
rect 15710 36194 15762 36206
rect 20190 36194 20242 36206
rect 24558 36258 24610 36270
rect 24558 36194 24610 36206
rect 25230 36258 25282 36270
rect 25230 36194 25282 36206
rect 25902 36258 25954 36270
rect 25902 36194 25954 36206
rect 26574 36258 26626 36270
rect 26574 36194 26626 36206
rect 27246 36258 27298 36270
rect 27246 36194 27298 36206
rect 1344 36090 38800 36124
rect 1344 36038 10538 36090
rect 10590 36038 10642 36090
rect 10694 36038 10746 36090
rect 10798 36038 19862 36090
rect 19914 36038 19966 36090
rect 20018 36038 20070 36090
rect 20122 36038 29186 36090
rect 29238 36038 29290 36090
rect 29342 36038 29394 36090
rect 29446 36038 38510 36090
rect 38562 36038 38614 36090
rect 38666 36038 38718 36090
rect 38770 36038 38800 36090
rect 1344 36004 38800 36038
rect 14030 35922 14082 35934
rect 14030 35858 14082 35870
rect 14590 35922 14642 35934
rect 14590 35858 14642 35870
rect 15262 35922 15314 35934
rect 15262 35858 15314 35870
rect 15934 35922 15986 35934
rect 15934 35858 15986 35870
rect 16494 35922 16546 35934
rect 16494 35858 16546 35870
rect 16942 35922 16994 35934
rect 16942 35858 16994 35870
rect 19854 35922 19906 35934
rect 19854 35858 19906 35870
rect 21422 35922 21474 35934
rect 21422 35858 21474 35870
rect 25454 35922 25506 35934
rect 25454 35858 25506 35870
rect 25902 35922 25954 35934
rect 25902 35858 25954 35870
rect 26350 35922 26402 35934
rect 26350 35858 26402 35870
rect 26910 35922 26962 35934
rect 26910 35858 26962 35870
rect 17726 35810 17778 35822
rect 17726 35746 17778 35758
rect 18062 35810 18114 35822
rect 18062 35746 18114 35758
rect 18398 35810 18450 35822
rect 18398 35746 18450 35758
rect 18734 35810 18786 35822
rect 18734 35746 18786 35758
rect 19070 35810 19122 35822
rect 19070 35746 19122 35758
rect 19406 35810 19458 35822
rect 19406 35746 19458 35758
rect 23326 35810 23378 35822
rect 23326 35746 23378 35758
rect 23998 35810 24050 35822
rect 23998 35746 24050 35758
rect 27134 35810 27186 35822
rect 27134 35746 27186 35758
rect 13346 35646 13358 35698
rect 13410 35646 13422 35698
rect 20514 35646 20526 35698
rect 20578 35646 20590 35698
rect 23538 35646 23550 35698
rect 23602 35646 23614 35698
rect 24210 35646 24222 35698
rect 24274 35646 24286 35698
rect 27346 35646 27358 35698
rect 27410 35646 27422 35698
rect 11442 35534 11454 35586
rect 11506 35534 11518 35586
rect 1344 35306 38640 35340
rect 1344 35254 5876 35306
rect 5928 35254 5980 35306
rect 6032 35254 6084 35306
rect 6136 35254 15200 35306
rect 15252 35254 15304 35306
rect 15356 35254 15408 35306
rect 15460 35254 24524 35306
rect 24576 35254 24628 35306
rect 24680 35254 24732 35306
rect 24784 35254 33848 35306
rect 33900 35254 33952 35306
rect 34004 35254 34056 35306
rect 34108 35254 38640 35306
rect 1344 35220 38640 35254
rect 12798 35026 12850 35038
rect 12798 34962 12850 34974
rect 18174 35026 18226 35038
rect 18174 34962 18226 34974
rect 18846 35026 18898 35038
rect 18846 34962 18898 34974
rect 21534 35026 21586 35038
rect 21534 34962 21586 34974
rect 23102 35026 23154 35038
rect 23102 34962 23154 34974
rect 23774 35026 23826 35038
rect 23774 34962 23826 34974
rect 21758 34914 21810 34926
rect 21758 34850 21810 34862
rect 22094 34690 22146 34702
rect 22094 34626 22146 34638
rect 24334 34690 24386 34702
rect 24334 34626 24386 34638
rect 1344 34522 38800 34556
rect 1344 34470 10538 34522
rect 10590 34470 10642 34522
rect 10694 34470 10746 34522
rect 10798 34470 19862 34522
rect 19914 34470 19966 34522
rect 20018 34470 20070 34522
rect 20122 34470 29186 34522
rect 29238 34470 29290 34522
rect 29342 34470 29394 34522
rect 29446 34470 38510 34522
rect 38562 34470 38614 34522
rect 38666 34470 38718 34522
rect 38770 34470 38800 34522
rect 1344 34436 38800 34470
rect 1344 33738 38640 33772
rect 1344 33686 5876 33738
rect 5928 33686 5980 33738
rect 6032 33686 6084 33738
rect 6136 33686 15200 33738
rect 15252 33686 15304 33738
rect 15356 33686 15408 33738
rect 15460 33686 24524 33738
rect 24576 33686 24628 33738
rect 24680 33686 24732 33738
rect 24784 33686 33848 33738
rect 33900 33686 33952 33738
rect 34004 33686 34056 33738
rect 34108 33686 38640 33738
rect 1344 33652 38640 33686
rect 1344 32954 38800 32988
rect 1344 32902 10538 32954
rect 10590 32902 10642 32954
rect 10694 32902 10746 32954
rect 10798 32902 19862 32954
rect 19914 32902 19966 32954
rect 20018 32902 20070 32954
rect 20122 32902 29186 32954
rect 29238 32902 29290 32954
rect 29342 32902 29394 32954
rect 29446 32902 38510 32954
rect 38562 32902 38614 32954
rect 38666 32902 38718 32954
rect 38770 32902 38800 32954
rect 1344 32868 38800 32902
rect 1344 32170 38640 32204
rect 1344 32118 5876 32170
rect 5928 32118 5980 32170
rect 6032 32118 6084 32170
rect 6136 32118 15200 32170
rect 15252 32118 15304 32170
rect 15356 32118 15408 32170
rect 15460 32118 24524 32170
rect 24576 32118 24628 32170
rect 24680 32118 24732 32170
rect 24784 32118 33848 32170
rect 33900 32118 33952 32170
rect 34004 32118 34056 32170
rect 34108 32118 38640 32170
rect 1344 32084 38640 32118
rect 1344 31386 38800 31420
rect 1344 31334 10538 31386
rect 10590 31334 10642 31386
rect 10694 31334 10746 31386
rect 10798 31334 19862 31386
rect 19914 31334 19966 31386
rect 20018 31334 20070 31386
rect 20122 31334 29186 31386
rect 29238 31334 29290 31386
rect 29342 31334 29394 31386
rect 29446 31334 38510 31386
rect 38562 31334 38614 31386
rect 38666 31334 38718 31386
rect 38770 31334 38800 31386
rect 1344 31300 38800 31334
rect 37886 31106 37938 31118
rect 37886 31042 37938 31054
rect 38222 30994 38274 31006
rect 38222 30930 38274 30942
rect 37662 30882 37714 30894
rect 37662 30818 37714 30830
rect 1344 30602 38640 30636
rect 1344 30550 5876 30602
rect 5928 30550 5980 30602
rect 6032 30550 6084 30602
rect 6136 30550 15200 30602
rect 15252 30550 15304 30602
rect 15356 30550 15408 30602
rect 15460 30550 24524 30602
rect 24576 30550 24628 30602
rect 24680 30550 24732 30602
rect 24784 30550 33848 30602
rect 33900 30550 33952 30602
rect 34004 30550 34056 30602
rect 34108 30550 38640 30602
rect 1344 30516 38640 30550
rect 37662 30098 37714 30110
rect 37662 30034 37714 30046
rect 38222 30098 38274 30110
rect 38222 30034 38274 30046
rect 37886 29986 37938 29998
rect 37886 29922 37938 29934
rect 1344 29818 38800 29852
rect 1344 29766 10538 29818
rect 10590 29766 10642 29818
rect 10694 29766 10746 29818
rect 10798 29766 19862 29818
rect 19914 29766 19966 29818
rect 20018 29766 20070 29818
rect 20122 29766 29186 29818
rect 29238 29766 29290 29818
rect 29342 29766 29394 29818
rect 29446 29766 38510 29818
rect 38562 29766 38614 29818
rect 38666 29766 38718 29818
rect 38770 29766 38800 29818
rect 1344 29732 38800 29766
rect 37886 29538 37938 29550
rect 37886 29474 37938 29486
rect 38222 29426 38274 29438
rect 4274 29374 4286 29426
rect 4338 29374 4350 29426
rect 38222 29362 38274 29374
rect 37662 29314 37714 29326
rect 37662 29250 37714 29262
rect 1934 29202 1986 29214
rect 1934 29138 1986 29150
rect 1344 29034 38640 29068
rect 1344 28982 5876 29034
rect 5928 28982 5980 29034
rect 6032 28982 6084 29034
rect 6136 28982 15200 29034
rect 15252 28982 15304 29034
rect 15356 28982 15408 29034
rect 15460 28982 24524 29034
rect 24576 28982 24628 29034
rect 24680 28982 24732 29034
rect 24784 28982 33848 29034
rect 33900 28982 33952 29034
rect 34004 28982 34056 29034
rect 34108 28982 38640 29034
rect 1344 28948 38640 28982
rect 1710 28642 1762 28654
rect 1710 28578 1762 28590
rect 2494 28642 2546 28654
rect 2494 28578 2546 28590
rect 37662 28642 37714 28654
rect 38098 28590 38110 28642
rect 38162 28590 38174 28642
rect 37662 28578 37714 28590
rect 37886 28530 37938 28542
rect 37886 28466 37938 28478
rect 2034 28366 2046 28418
rect 2098 28366 2110 28418
rect 1344 28250 38800 28284
rect 1344 28198 10538 28250
rect 10590 28198 10642 28250
rect 10694 28198 10746 28250
rect 10798 28198 19862 28250
rect 19914 28198 19966 28250
rect 20018 28198 20070 28250
rect 20122 28198 29186 28250
rect 29238 28198 29290 28250
rect 29342 28198 29394 28250
rect 29446 28198 38510 28250
rect 38562 28198 38614 28250
rect 38666 28198 38718 28250
rect 38770 28198 38800 28250
rect 1344 28164 38800 28198
rect 20514 28030 20526 28082
rect 20578 28030 20590 28082
rect 37886 27970 37938 27982
rect 2034 27918 2046 27970
rect 2098 27918 2110 27970
rect 19842 27918 19854 27970
rect 19906 27918 19918 27970
rect 20290 27918 20302 27970
rect 20354 27918 20366 27970
rect 37886 27906 37938 27918
rect 1710 27858 1762 27870
rect 38222 27858 38274 27870
rect 19506 27806 19518 27858
rect 19570 27806 19582 27858
rect 1710 27794 1762 27806
rect 38222 27794 38274 27806
rect 2494 27746 2546 27758
rect 2494 27682 2546 27694
rect 2942 27746 2994 27758
rect 2942 27682 2994 27694
rect 37214 27746 37266 27758
rect 37214 27682 37266 27694
rect 37662 27746 37714 27758
rect 37662 27682 37714 27694
rect 1344 27466 38640 27500
rect 1344 27414 5876 27466
rect 5928 27414 5980 27466
rect 6032 27414 6084 27466
rect 6136 27414 15200 27466
rect 15252 27414 15304 27466
rect 15356 27414 15408 27466
rect 15460 27414 24524 27466
rect 24576 27414 24628 27466
rect 24680 27414 24732 27466
rect 24784 27414 33848 27466
rect 33900 27414 33952 27466
rect 34004 27414 34056 27466
rect 34108 27414 38640 27466
rect 1344 27380 38640 27414
rect 19842 27246 19854 27298
rect 19906 27246 19918 27298
rect 17490 27134 17502 27186
rect 17554 27134 17566 27186
rect 16270 27074 16322 27086
rect 20638 27074 20690 27086
rect 1810 27022 1822 27074
rect 1874 27022 1886 27074
rect 16482 27022 16494 27074
rect 16546 27022 16558 27074
rect 17602 27022 17614 27074
rect 17666 27022 17678 27074
rect 18722 27022 18734 27074
rect 18786 27022 18798 27074
rect 19730 27022 19742 27074
rect 19794 27022 19806 27074
rect 20178 27022 20190 27074
rect 20242 27022 20254 27074
rect 16270 27010 16322 27022
rect 20638 27010 20690 27022
rect 37662 27074 37714 27086
rect 38098 27022 38110 27074
rect 38162 27022 38174 27074
rect 37662 27010 37714 27022
rect 2046 26962 2098 26974
rect 2046 26898 2098 26910
rect 2382 26962 2434 26974
rect 2382 26898 2434 26910
rect 3166 26962 3218 26974
rect 3166 26898 3218 26910
rect 17054 26962 17106 26974
rect 17054 26898 17106 26910
rect 18174 26962 18226 26974
rect 21310 26962 21362 26974
rect 18498 26910 18510 26962
rect 18562 26910 18574 26962
rect 18174 26898 18226 26910
rect 21310 26898 21362 26910
rect 21646 26962 21698 26974
rect 21646 26898 21698 26910
rect 37326 26962 37378 26974
rect 37326 26898 37378 26910
rect 2718 26850 2770 26862
rect 2718 26786 2770 26798
rect 21534 26850 21586 26862
rect 21534 26786 21586 26798
rect 36990 26850 37042 26862
rect 36990 26786 37042 26798
rect 1344 26682 38800 26716
rect 1344 26630 10538 26682
rect 10590 26630 10642 26682
rect 10694 26630 10746 26682
rect 10798 26630 19862 26682
rect 19914 26630 19966 26682
rect 20018 26630 20070 26682
rect 20122 26630 29186 26682
rect 29238 26630 29290 26682
rect 29342 26630 29394 26682
rect 29446 26630 38510 26682
rect 38562 26630 38614 26682
rect 38666 26630 38718 26682
rect 38770 26630 38800 26682
rect 1344 26596 38800 26630
rect 15038 26514 15090 26526
rect 15038 26450 15090 26462
rect 17726 26514 17778 26526
rect 17726 26450 17778 26462
rect 37662 26514 37714 26526
rect 37662 26450 37714 26462
rect 2046 26402 2098 26414
rect 2046 26338 2098 26350
rect 14814 26402 14866 26414
rect 14814 26338 14866 26350
rect 37886 26402 37938 26414
rect 37886 26338 37938 26350
rect 1710 26290 1762 26302
rect 1710 26226 1762 26238
rect 14702 26290 14754 26302
rect 38222 26290 38274 26302
rect 15586 26238 15598 26290
rect 15650 26238 15662 26290
rect 16594 26238 16606 26290
rect 16658 26238 16670 26290
rect 18498 26238 18510 26290
rect 18562 26238 18574 26290
rect 19506 26238 19518 26290
rect 19570 26238 19582 26290
rect 20290 26238 20302 26290
rect 20354 26238 20366 26290
rect 20962 26238 20974 26290
rect 21026 26238 21038 26290
rect 14702 26226 14754 26238
rect 38222 26226 38274 26238
rect 2494 26178 2546 26190
rect 37214 26178 37266 26190
rect 15810 26126 15822 26178
rect 15874 26126 15886 26178
rect 16370 26126 16382 26178
rect 16434 26126 16446 26178
rect 21410 26126 21422 26178
rect 21474 26126 21486 26178
rect 2494 26114 2546 26126
rect 37214 26114 37266 26126
rect 19618 26014 19630 26066
rect 19682 26014 19694 26066
rect 1344 25898 38640 25932
rect 1344 25846 5876 25898
rect 5928 25846 5980 25898
rect 6032 25846 6084 25898
rect 6136 25846 15200 25898
rect 15252 25846 15304 25898
rect 15356 25846 15408 25898
rect 15460 25846 24524 25898
rect 24576 25846 24628 25898
rect 24680 25846 24732 25898
rect 24784 25846 33848 25898
rect 33900 25846 33952 25898
rect 34004 25846 34056 25898
rect 34108 25846 38640 25898
rect 1344 25812 38640 25846
rect 14366 25730 14418 25742
rect 14366 25666 14418 25678
rect 14702 25730 14754 25742
rect 14702 25666 14754 25678
rect 19182 25618 19234 25630
rect 15698 25566 15710 25618
rect 15762 25566 15774 25618
rect 16482 25566 16494 25618
rect 16546 25566 16558 25618
rect 19182 25554 19234 25566
rect 21870 25618 21922 25630
rect 21870 25554 21922 25566
rect 13682 25454 13694 25506
rect 13746 25454 13758 25506
rect 15586 25454 15598 25506
rect 15650 25454 15662 25506
rect 16594 25454 16606 25506
rect 16658 25454 16670 25506
rect 17378 25454 17390 25506
rect 17442 25454 17454 25506
rect 18610 25454 18622 25506
rect 18674 25454 18686 25506
rect 19618 25454 19630 25506
rect 19682 25454 19694 25506
rect 22194 25454 22206 25506
rect 22258 25454 22270 25506
rect 22642 25454 22654 25506
rect 22706 25454 22718 25506
rect 23426 25454 23438 25506
rect 23490 25454 23502 25506
rect 23986 25454 23998 25506
rect 24050 25454 24062 25506
rect 24882 25454 24894 25506
rect 24946 25454 24958 25506
rect 1710 25394 1762 25406
rect 21422 25394 21474 25406
rect 13570 25342 13582 25394
rect 13634 25342 13646 25394
rect 20066 25342 20078 25394
rect 20130 25342 20142 25394
rect 1710 25330 1762 25342
rect 21422 25330 21474 25342
rect 21534 25394 21586 25406
rect 37662 25394 37714 25406
rect 22866 25342 22878 25394
rect 22930 25342 22942 25394
rect 21534 25330 21586 25342
rect 37662 25330 37714 25342
rect 38222 25394 38274 25406
rect 38222 25330 38274 25342
rect 2046 25282 2098 25294
rect 2046 25218 2098 25230
rect 2494 25282 2546 25294
rect 2494 25218 2546 25230
rect 21198 25282 21250 25294
rect 21198 25218 21250 25230
rect 37886 25282 37938 25294
rect 37886 25218 37938 25230
rect 1344 25114 38800 25148
rect 1344 25062 10538 25114
rect 10590 25062 10642 25114
rect 10694 25062 10746 25114
rect 10798 25062 19862 25114
rect 19914 25062 19966 25114
rect 20018 25062 20070 25114
rect 20122 25062 29186 25114
rect 29238 25062 29290 25114
rect 29342 25062 29394 25114
rect 29446 25062 38510 25114
rect 38562 25062 38614 25114
rect 38666 25062 38718 25114
rect 38770 25062 38800 25114
rect 1344 25028 38800 25062
rect 22878 24946 22930 24958
rect 22878 24882 22930 24894
rect 22654 24834 22706 24846
rect 2034 24782 2046 24834
rect 2098 24782 2110 24834
rect 16258 24782 16270 24834
rect 16322 24782 16334 24834
rect 22654 24770 22706 24782
rect 22990 24834 23042 24846
rect 37886 24834 37938 24846
rect 26562 24782 26574 24834
rect 26626 24782 26638 24834
rect 22990 24770 23042 24782
rect 37886 24770 37938 24782
rect 1710 24722 1762 24734
rect 1710 24658 1762 24670
rect 12350 24722 12402 24734
rect 13134 24722 13186 24734
rect 27022 24722 27074 24734
rect 38222 24722 38274 24734
rect 12562 24670 12574 24722
rect 12626 24670 12638 24722
rect 14690 24670 14702 24722
rect 14754 24670 14766 24722
rect 15698 24670 15710 24722
rect 15762 24670 15774 24722
rect 17938 24670 17950 24722
rect 18002 24670 18014 24722
rect 18722 24670 18734 24722
rect 18786 24670 18798 24722
rect 20290 24670 20302 24722
rect 20354 24670 20366 24722
rect 20962 24670 20974 24722
rect 21026 24670 21038 24722
rect 25890 24670 25902 24722
rect 25954 24670 25966 24722
rect 26450 24670 26462 24722
rect 26514 24670 26526 24722
rect 27794 24670 27806 24722
rect 27858 24670 27870 24722
rect 28690 24670 28702 24722
rect 28754 24670 28766 24722
rect 12350 24658 12402 24670
rect 13134 24658 13186 24670
rect 27022 24658 27074 24670
rect 38222 24658 38274 24670
rect 2494 24610 2546 24622
rect 25566 24610 25618 24622
rect 14578 24558 14590 24610
rect 14642 24558 14654 24610
rect 21746 24558 21758 24610
rect 21810 24558 21822 24610
rect 2494 24546 2546 24558
rect 25566 24546 25618 24558
rect 37662 24610 37714 24622
rect 37662 24546 37714 24558
rect 15810 24446 15822 24498
rect 15874 24446 15886 24498
rect 19618 24446 19630 24498
rect 19682 24446 19694 24498
rect 1344 24330 38640 24364
rect 1344 24278 5876 24330
rect 5928 24278 5980 24330
rect 6032 24278 6084 24330
rect 6136 24278 15200 24330
rect 15252 24278 15304 24330
rect 15356 24278 15408 24330
rect 15460 24278 24524 24330
rect 24576 24278 24628 24330
rect 24680 24278 24732 24330
rect 24784 24278 33848 24330
rect 33900 24278 33952 24330
rect 34004 24278 34056 24330
rect 34108 24278 38640 24330
rect 1344 24244 38640 24278
rect 14578 24110 14590 24162
rect 14642 24110 14654 24162
rect 17826 24110 17838 24162
rect 17890 24110 17902 24162
rect 21870 24050 21922 24062
rect 12450 23998 12462 24050
rect 12514 23998 12526 24050
rect 16706 23998 16718 24050
rect 16770 23998 16782 24050
rect 21870 23986 21922 23998
rect 21198 23938 21250 23950
rect 14354 23886 14366 23938
rect 14418 23886 14430 23938
rect 14690 23886 14702 23938
rect 14754 23886 14766 23938
rect 15586 23886 15598 23938
rect 15650 23886 15662 23938
rect 17490 23886 17502 23938
rect 17554 23886 17566 23938
rect 18610 23886 18622 23938
rect 18674 23886 18686 23938
rect 19618 23886 19630 23938
rect 19682 23886 19694 23938
rect 22194 23886 22206 23938
rect 22258 23886 22270 23938
rect 22754 23886 22766 23938
rect 22818 23886 22830 23938
rect 23426 23886 23438 23938
rect 23490 23886 23502 23938
rect 24098 23886 24110 23938
rect 24162 23886 24174 23938
rect 24994 23886 25006 23938
rect 25058 23886 25070 23938
rect 21198 23874 21250 23886
rect 21422 23826 21474 23838
rect 20066 23774 20078 23826
rect 20130 23774 20142 23826
rect 21422 23762 21474 23774
rect 21534 23826 21586 23838
rect 21534 23762 21586 23774
rect 38222 23826 38274 23838
rect 38222 23762 38274 23774
rect 1710 23714 1762 23726
rect 2494 23714 2546 23726
rect 2034 23662 2046 23714
rect 2098 23662 2110 23714
rect 1710 23650 1762 23662
rect 2494 23650 2546 23662
rect 12910 23714 12962 23726
rect 12910 23650 12962 23662
rect 13918 23714 13970 23726
rect 13918 23650 13970 23662
rect 16270 23714 16322 23726
rect 37662 23714 37714 23726
rect 22866 23662 22878 23714
rect 22930 23662 22942 23714
rect 16270 23650 16322 23662
rect 37662 23650 37714 23662
rect 37886 23714 37938 23726
rect 37886 23650 37938 23662
rect 1344 23546 38800 23580
rect 1344 23494 10538 23546
rect 10590 23494 10642 23546
rect 10694 23494 10746 23546
rect 10798 23494 19862 23546
rect 19914 23494 19966 23546
rect 20018 23494 20070 23546
rect 20122 23494 29186 23546
rect 29238 23494 29290 23546
rect 29342 23494 29394 23546
rect 29446 23494 38510 23546
rect 38562 23494 38614 23546
rect 38666 23494 38718 23546
rect 38770 23494 38800 23546
rect 1344 23460 38800 23494
rect 21410 23326 21422 23378
rect 21474 23326 21486 23378
rect 26450 23326 26462 23378
rect 26514 23326 26526 23378
rect 2034 23214 2046 23266
rect 2098 23214 2110 23266
rect 16706 23214 16718 23266
rect 16770 23214 16782 23266
rect 18610 23214 18622 23266
rect 18674 23214 18686 23266
rect 23538 23214 23550 23266
rect 23602 23214 23614 23266
rect 37874 23214 37886 23266
rect 37938 23214 37950 23266
rect 1710 23154 1762 23166
rect 1710 23090 1762 23102
rect 13582 23154 13634 23166
rect 17390 23154 17442 23166
rect 20078 23154 20130 23166
rect 21086 23154 21138 23166
rect 38222 23154 38274 23166
rect 15026 23102 15038 23154
rect 15090 23102 15102 23154
rect 15586 23102 15598 23154
rect 15650 23102 15662 23154
rect 17826 23102 17838 23154
rect 17890 23102 17902 23154
rect 19170 23102 19182 23154
rect 19234 23102 19246 23154
rect 19730 23102 19742 23154
rect 19794 23102 19806 23154
rect 20402 23102 20414 23154
rect 20466 23102 20478 23154
rect 23314 23102 23326 23154
rect 23378 23102 23390 23154
rect 25778 23102 25790 23154
rect 25842 23102 25854 23154
rect 26338 23102 26350 23154
rect 26402 23102 26414 23154
rect 27010 23102 27022 23154
rect 27074 23102 27086 23154
rect 27682 23102 27694 23154
rect 27746 23102 27758 23154
rect 28466 23102 28478 23154
rect 28530 23102 28542 23154
rect 13582 23090 13634 23102
rect 17390 23090 17442 23102
rect 20078 23090 20130 23102
rect 21086 23090 21138 23102
rect 38222 23090 38274 23102
rect 2494 23042 2546 23054
rect 25454 23042 25506 23054
rect 13122 22990 13134 23042
rect 13186 22990 13198 23042
rect 14466 22990 14478 23042
rect 14530 22990 14542 23042
rect 2494 22978 2546 22990
rect 25454 22978 25506 22990
rect 37662 23042 37714 23054
rect 37662 22978 37714 22990
rect 20178 22878 20190 22930
rect 20242 22878 20254 22930
rect 1344 22762 38640 22796
rect 1344 22710 5876 22762
rect 5928 22710 5980 22762
rect 6032 22710 6084 22762
rect 6136 22710 15200 22762
rect 15252 22710 15304 22762
rect 15356 22710 15408 22762
rect 15460 22710 24524 22762
rect 24576 22710 24628 22762
rect 24680 22710 24732 22762
rect 24784 22710 33848 22762
rect 33900 22710 33952 22762
rect 34004 22710 34056 22762
rect 34108 22710 38640 22762
rect 1344 22676 38640 22710
rect 20402 22542 20414 22594
rect 20466 22591 20478 22594
rect 20850 22591 20862 22594
rect 20466 22545 20862 22591
rect 20466 22542 20478 22545
rect 20850 22542 20862 22545
rect 20914 22542 20926 22594
rect 15586 22430 15598 22482
rect 15650 22430 15662 22482
rect 17714 22430 17726 22482
rect 17778 22430 17790 22482
rect 20066 22430 20078 22482
rect 20130 22430 20142 22482
rect 19630 22370 19682 22382
rect 13794 22318 13806 22370
rect 13858 22318 13870 22370
rect 15922 22318 15934 22370
rect 15986 22318 15998 22370
rect 16818 22318 16830 22370
rect 16882 22318 16894 22370
rect 17602 22318 17614 22370
rect 17666 22318 17678 22370
rect 18498 22318 18510 22370
rect 18562 22318 18574 22370
rect 19630 22306 19682 22318
rect 1710 22258 1762 22270
rect 21534 22258 21586 22270
rect 2034 22206 2046 22258
rect 2098 22206 2110 22258
rect 1710 22194 1762 22206
rect 21534 22194 21586 22206
rect 21870 22258 21922 22270
rect 21870 22194 21922 22206
rect 21982 22258 22034 22270
rect 21982 22194 22034 22206
rect 36542 22258 36594 22270
rect 36542 22194 36594 22206
rect 37550 22258 37602 22270
rect 37550 22194 37602 22206
rect 38222 22258 38274 22270
rect 38222 22194 38274 22206
rect 2382 22146 2434 22158
rect 3166 22146 3218 22158
rect 2706 22094 2718 22146
rect 2770 22094 2782 22146
rect 2382 22082 2434 22094
rect 3166 22082 3218 22094
rect 14478 22146 14530 22158
rect 14478 22082 14530 22094
rect 20638 22146 20690 22158
rect 20638 22082 20690 22094
rect 21198 22146 21250 22158
rect 21198 22082 21250 22094
rect 21422 22146 21474 22158
rect 21422 22082 21474 22094
rect 22206 22146 22258 22158
rect 22206 22082 22258 22094
rect 23438 22146 23490 22158
rect 23438 22082 23490 22094
rect 24222 22146 24274 22158
rect 24222 22082 24274 22094
rect 37214 22146 37266 22158
rect 37214 22082 37266 22094
rect 37886 22146 37938 22158
rect 37886 22082 37938 22094
rect 1344 21978 38800 22012
rect 1344 21926 10538 21978
rect 10590 21926 10642 21978
rect 10694 21926 10746 21978
rect 10798 21926 19862 21978
rect 19914 21926 19966 21978
rect 20018 21926 20070 21978
rect 20122 21926 29186 21978
rect 29238 21926 29290 21978
rect 29342 21926 29394 21978
rect 29446 21926 38510 21978
rect 38562 21926 38614 21978
rect 38666 21926 38718 21978
rect 38770 21926 38800 21978
rect 1344 21892 38800 21926
rect 2494 21810 2546 21822
rect 2494 21746 2546 21758
rect 17390 21810 17442 21822
rect 17390 21746 17442 21758
rect 37886 21698 37938 21710
rect 2034 21646 2046 21698
rect 2098 21646 2110 21698
rect 19730 21646 19742 21698
rect 19794 21646 19806 21698
rect 20402 21646 20414 21698
rect 20466 21646 20478 21698
rect 21074 21646 21086 21698
rect 21138 21646 21150 21698
rect 23986 21646 23998 21698
rect 24050 21646 24062 21698
rect 37886 21634 37938 21646
rect 1710 21586 1762 21598
rect 25230 21586 25282 21598
rect 12338 21534 12350 21586
rect 12402 21534 12414 21586
rect 13570 21534 13582 21586
rect 13634 21534 13646 21586
rect 14914 21534 14926 21586
rect 14978 21534 14990 21586
rect 15362 21534 15374 21586
rect 15426 21534 15438 21586
rect 19506 21534 19518 21586
rect 19570 21534 19582 21586
rect 20514 21534 20526 21586
rect 20578 21534 20590 21586
rect 21410 21534 21422 21586
rect 21474 21534 21486 21586
rect 22082 21534 22094 21586
rect 22146 21534 22158 21586
rect 23762 21534 23774 21586
rect 23826 21534 23838 21586
rect 1710 21522 1762 21534
rect 25230 21522 25282 21534
rect 25790 21586 25842 21598
rect 25790 21522 25842 21534
rect 37550 21586 37602 21598
rect 37550 21522 37602 21534
rect 38222 21586 38274 21598
rect 38222 21522 38274 21534
rect 2942 21474 2994 21486
rect 2942 21410 2994 21422
rect 12126 21474 12178 21486
rect 17950 21474 18002 21486
rect 23214 21474 23266 21486
rect 15810 21422 15822 21474
rect 15874 21422 15886 21474
rect 18498 21422 18510 21474
rect 18562 21422 18574 21474
rect 20290 21422 20302 21474
rect 20354 21422 20366 21474
rect 22866 21422 22878 21474
rect 22930 21422 22942 21474
rect 12126 21410 12178 21422
rect 17950 21410 18002 21422
rect 23214 21410 23266 21422
rect 24446 21474 24498 21486
rect 24446 21410 24498 21422
rect 37214 21474 37266 21486
rect 37214 21410 37266 21422
rect 24334 21362 24386 21374
rect 15698 21310 15710 21362
rect 15762 21310 15774 21362
rect 24334 21298 24386 21310
rect 1344 21194 38640 21228
rect 1344 21142 5876 21194
rect 5928 21142 5980 21194
rect 6032 21142 6084 21194
rect 6136 21142 15200 21194
rect 15252 21142 15304 21194
rect 15356 21142 15408 21194
rect 15460 21142 24524 21194
rect 24576 21142 24628 21194
rect 24680 21142 24732 21194
rect 24784 21142 33848 21194
rect 33900 21142 33952 21194
rect 34004 21142 34056 21194
rect 34108 21142 38640 21194
rect 1344 21108 38640 21142
rect 20638 21026 20690 21038
rect 17378 20974 17390 21026
rect 17442 20974 17454 21026
rect 20638 20962 20690 20974
rect 28254 20914 28306 20926
rect 12450 20862 12462 20914
rect 12514 20862 12526 20914
rect 16930 20862 16942 20914
rect 16994 20862 17006 20914
rect 28254 20850 28306 20862
rect 11342 20802 11394 20814
rect 11342 20738 11394 20750
rect 12910 20802 12962 20814
rect 18958 20802 19010 20814
rect 13458 20750 13470 20802
rect 13522 20750 13534 20802
rect 13794 20750 13806 20802
rect 13858 20750 13870 20802
rect 15362 20750 15374 20802
rect 15426 20750 15438 20802
rect 16818 20750 16830 20802
rect 16882 20750 16894 20802
rect 12910 20738 12962 20750
rect 18958 20738 19010 20750
rect 20078 20802 20130 20814
rect 20078 20738 20130 20750
rect 20190 20802 20242 20814
rect 20190 20738 20242 20750
rect 20526 20802 20578 20814
rect 21298 20750 21310 20802
rect 21362 20750 21374 20802
rect 22306 20750 22318 20802
rect 22370 20750 22382 20802
rect 23426 20750 23438 20802
rect 23490 20750 23502 20802
rect 24322 20750 24334 20802
rect 24386 20750 24398 20802
rect 24882 20750 24894 20802
rect 24946 20750 24958 20802
rect 25554 20750 25566 20802
rect 25618 20750 25630 20802
rect 26226 20750 26238 20802
rect 26290 20750 26302 20802
rect 27122 20750 27134 20802
rect 27186 20750 27198 20802
rect 20526 20738 20578 20750
rect 11790 20690 11842 20702
rect 11790 20626 11842 20638
rect 18286 20690 18338 20702
rect 23998 20690 24050 20702
rect 22530 20638 22542 20690
rect 22594 20638 22606 20690
rect 23090 20638 23102 20690
rect 23154 20638 23166 20690
rect 18286 20626 18338 20638
rect 23998 20626 24050 20638
rect 27806 20690 27858 20702
rect 27806 20626 27858 20638
rect 38222 20690 38274 20702
rect 38222 20626 38274 20638
rect 1710 20578 1762 20590
rect 2494 20578 2546 20590
rect 21198 20578 21250 20590
rect 37662 20578 37714 20590
rect 2034 20526 2046 20578
rect 2098 20526 2110 20578
rect 18610 20526 18622 20578
rect 18674 20526 18686 20578
rect 24994 20526 25006 20578
rect 25058 20526 25070 20578
rect 1710 20514 1762 20526
rect 2494 20514 2546 20526
rect 21198 20514 21250 20526
rect 37662 20514 37714 20526
rect 37886 20578 37938 20590
rect 37886 20514 37938 20526
rect 1344 20410 38800 20444
rect 1344 20358 10538 20410
rect 10590 20358 10642 20410
rect 10694 20358 10746 20410
rect 10798 20358 19862 20410
rect 19914 20358 19966 20410
rect 20018 20358 20070 20410
rect 20122 20358 29186 20410
rect 29238 20358 29290 20410
rect 29342 20358 29394 20410
rect 29446 20358 38510 20410
rect 38562 20358 38614 20410
rect 38666 20358 38718 20410
rect 38770 20358 38800 20410
rect 1344 20324 38800 20358
rect 25790 20242 25842 20254
rect 22082 20190 22094 20242
rect 22146 20190 22158 20242
rect 25790 20178 25842 20190
rect 2046 20130 2098 20142
rect 21310 20130 21362 20142
rect 18162 20078 18174 20130
rect 18226 20078 18238 20130
rect 2046 20066 2098 20078
rect 21310 20066 21362 20078
rect 21758 20130 21810 20142
rect 21758 20066 21810 20078
rect 22542 20130 22594 20142
rect 22542 20066 22594 20078
rect 23214 20130 23266 20142
rect 37886 20130 37938 20142
rect 24658 20078 24670 20130
rect 24722 20078 24734 20130
rect 23214 20066 23266 20078
rect 37886 20066 37938 20078
rect 1710 20018 1762 20030
rect 21534 20018 21586 20030
rect 12338 19966 12350 20018
rect 12402 19966 12414 20018
rect 13570 19966 13582 20018
rect 13634 19966 13646 20018
rect 14914 19966 14926 20018
rect 14978 19966 14990 20018
rect 15362 19966 15374 20018
rect 15426 19966 15438 20018
rect 17602 19966 17614 20018
rect 17666 19966 17678 20018
rect 19282 19966 19294 20018
rect 19346 19966 19358 20018
rect 1710 19954 1762 19966
rect 21534 19954 21586 19966
rect 21646 20018 21698 20030
rect 21646 19954 21698 19966
rect 22654 20018 22706 20030
rect 22654 19954 22706 19966
rect 22766 20018 22818 20030
rect 23774 20018 23826 20030
rect 38222 20018 38274 20030
rect 23426 19966 23438 20018
rect 23490 19966 23502 20018
rect 24434 19966 24446 20018
rect 24498 19966 24510 20018
rect 26898 19966 26910 20018
rect 26962 19966 26974 20018
rect 27458 19966 27470 20018
rect 27522 19966 27534 20018
rect 28802 19966 28814 20018
rect 28866 19966 28878 20018
rect 29922 19966 29934 20018
rect 29986 19966 29998 20018
rect 22766 19954 22818 19966
rect 23774 19954 23826 19966
rect 38222 19954 38274 19966
rect 2494 19906 2546 19918
rect 25230 19906 25282 19918
rect 15810 19854 15822 19906
rect 15874 19854 15886 19906
rect 19170 19854 19182 19906
rect 19234 19854 19246 19906
rect 2494 19842 2546 19854
rect 25230 19842 25282 19854
rect 26238 19906 26290 19918
rect 26238 19842 26290 19854
rect 26574 19906 26626 19918
rect 26574 19842 26626 19854
rect 27694 19906 27746 19918
rect 27694 19842 27746 19854
rect 37662 19906 37714 19918
rect 37662 19842 37714 19854
rect 23102 19794 23154 19806
rect 15698 19742 15710 19794
rect 15762 19742 15774 19794
rect 18722 19742 18734 19794
rect 18786 19742 18798 19794
rect 23102 19730 23154 19742
rect 28478 19794 28530 19806
rect 28478 19730 28530 19742
rect 1344 19626 38640 19660
rect 1344 19574 5876 19626
rect 5928 19574 5980 19626
rect 6032 19574 6084 19626
rect 6136 19574 15200 19626
rect 15252 19574 15304 19626
rect 15356 19574 15408 19626
rect 15460 19574 24524 19626
rect 24576 19574 24628 19626
rect 24680 19574 24732 19626
rect 24784 19574 33848 19626
rect 33900 19574 33952 19626
rect 34004 19574 34056 19626
rect 34108 19574 38640 19626
rect 1344 19540 38640 19574
rect 18946 19406 18958 19458
rect 19010 19406 19022 19458
rect 1934 19346 1986 19358
rect 12910 19346 12962 19358
rect 25342 19346 25394 19358
rect 12226 19294 12238 19346
rect 12290 19294 12302 19346
rect 15586 19294 15598 19346
rect 15650 19294 15662 19346
rect 17042 19294 17054 19346
rect 17106 19294 17118 19346
rect 1934 19282 1986 19294
rect 12910 19282 12962 19294
rect 25342 19282 25394 19294
rect 12574 19234 12626 19246
rect 18174 19234 18226 19246
rect 19630 19234 19682 19246
rect 4274 19182 4286 19234
rect 4338 19182 4350 19234
rect 13458 19182 13470 19234
rect 13522 19182 13534 19234
rect 13794 19182 13806 19234
rect 13858 19182 13870 19234
rect 15362 19182 15374 19234
rect 15426 19182 15438 19234
rect 16818 19182 16830 19234
rect 16882 19182 16894 19234
rect 19394 19182 19406 19234
rect 19458 19182 19470 19234
rect 12574 19170 12626 19182
rect 18174 19170 18226 19182
rect 19630 19170 19682 19182
rect 20302 19234 20354 19246
rect 20302 19170 20354 19182
rect 21646 19234 21698 19246
rect 21646 19170 21698 19182
rect 21982 19234 22034 19246
rect 25778 19182 25790 19234
rect 25842 19182 25854 19234
rect 26226 19182 26238 19234
rect 26290 19182 26302 19234
rect 26898 19182 26910 19234
rect 26962 19182 26974 19234
rect 27570 19182 27582 19234
rect 27634 19182 27646 19234
rect 28466 19182 28478 19234
rect 28530 19182 28542 19234
rect 21982 19170 22034 19182
rect 18510 19122 18562 19134
rect 18510 19058 18562 19070
rect 19966 19122 20018 19134
rect 19966 19058 20018 19070
rect 21870 19122 21922 19134
rect 37886 19122 37938 19134
rect 26338 19070 26350 19122
rect 26402 19070 26414 19122
rect 21870 19058 21922 19070
rect 37886 19058 37938 19070
rect 38222 19122 38274 19134
rect 38222 19058 38274 19070
rect 18398 19010 18450 19022
rect 18398 18946 18450 18958
rect 37662 19010 37714 19022
rect 37662 18946 37714 18958
rect 1344 18842 38800 18876
rect 1344 18790 10538 18842
rect 10590 18790 10642 18842
rect 10694 18790 10746 18842
rect 10798 18790 19862 18842
rect 19914 18790 19966 18842
rect 20018 18790 20070 18842
rect 20122 18790 29186 18842
rect 29238 18790 29290 18842
rect 29342 18790 29394 18842
rect 29446 18790 38510 18842
rect 38562 18790 38614 18842
rect 38666 18790 38718 18842
rect 38770 18790 38800 18842
rect 1344 18756 38800 18790
rect 37886 18674 37938 18686
rect 37886 18610 37938 18622
rect 22206 18562 22258 18574
rect 2034 18510 2046 18562
rect 2098 18510 2110 18562
rect 16258 18510 16270 18562
rect 16322 18510 16334 18562
rect 22206 18498 22258 18510
rect 1710 18450 1762 18462
rect 17950 18450 18002 18462
rect 13458 18398 13470 18450
rect 13522 18398 13534 18450
rect 14690 18398 14702 18450
rect 14754 18398 14766 18450
rect 15586 18398 15598 18450
rect 15650 18398 15662 18450
rect 1710 18386 1762 18398
rect 17950 18386 18002 18398
rect 18958 18450 19010 18462
rect 20414 18450 20466 18462
rect 22542 18450 22594 18462
rect 19730 18398 19742 18450
rect 19794 18398 19806 18450
rect 21522 18398 21534 18450
rect 21586 18398 21598 18450
rect 18958 18386 19010 18398
rect 20414 18386 20466 18398
rect 22542 18386 22594 18398
rect 22878 18450 22930 18462
rect 22878 18386 22930 18398
rect 25230 18450 25282 18462
rect 25230 18386 25282 18398
rect 38222 18450 38274 18462
rect 38222 18386 38274 18398
rect 2494 18338 2546 18350
rect 2494 18274 2546 18286
rect 17390 18338 17442 18350
rect 17390 18274 17442 18286
rect 18398 18338 18450 18350
rect 18398 18274 18450 18286
rect 19294 18338 19346 18350
rect 19294 18274 19346 18286
rect 21086 18338 21138 18350
rect 21086 18274 21138 18286
rect 22990 18338 23042 18350
rect 22990 18274 23042 18286
rect 25790 18338 25842 18350
rect 25790 18274 25842 18286
rect 37662 18338 37714 18350
rect 37662 18274 37714 18286
rect 15922 18174 15934 18226
rect 15986 18174 15998 18226
rect 1344 18058 38640 18092
rect 1344 18006 5876 18058
rect 5928 18006 5980 18058
rect 6032 18006 6084 18058
rect 6136 18006 15200 18058
rect 15252 18006 15304 18058
rect 15356 18006 15408 18058
rect 15460 18006 24524 18058
rect 24576 18006 24628 18058
rect 24680 18006 24732 18058
rect 24784 18006 33848 18058
rect 33900 18006 33952 18058
rect 34004 18006 34056 18058
rect 34108 18006 38640 18058
rect 1344 17972 38640 18006
rect 12798 17890 12850 17902
rect 16818 17838 16830 17890
rect 16882 17838 16894 17890
rect 12798 17826 12850 17838
rect 1934 17778 1986 17790
rect 1934 17714 1986 17726
rect 11790 17778 11842 17790
rect 14802 17726 14814 17778
rect 14866 17726 14878 17778
rect 11790 17714 11842 17726
rect 19406 17666 19458 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 12226 17614 12238 17666
rect 12290 17614 12302 17666
rect 13010 17614 13022 17666
rect 13074 17614 13086 17666
rect 13794 17614 13806 17666
rect 13858 17614 13870 17666
rect 14018 17614 14030 17666
rect 14082 17614 14094 17666
rect 14914 17614 14926 17666
rect 14978 17614 14990 17666
rect 15474 17614 15486 17666
rect 15538 17614 15550 17666
rect 16594 17614 16606 17666
rect 16658 17614 16670 17666
rect 17714 17614 17726 17666
rect 17778 17614 17790 17666
rect 19406 17602 19458 17614
rect 19630 17666 19682 17678
rect 19630 17602 19682 17614
rect 19966 17666 20018 17678
rect 19966 17602 20018 17614
rect 21646 17666 21698 17678
rect 21646 17602 21698 17614
rect 22990 17666 23042 17678
rect 23426 17614 23438 17666
rect 23490 17614 23502 17666
rect 25778 17614 25790 17666
rect 25842 17614 25854 17666
rect 26226 17614 26238 17666
rect 26290 17614 26302 17666
rect 26898 17614 26910 17666
rect 26962 17614 26974 17666
rect 27346 17614 27358 17666
rect 27410 17614 27422 17666
rect 28466 17614 28478 17666
rect 28530 17614 28542 17666
rect 22990 17602 23042 17614
rect 19854 17554 19906 17566
rect 18162 17502 18174 17554
rect 18226 17502 18238 17554
rect 19058 17502 19070 17554
rect 19122 17502 19134 17554
rect 19854 17490 19906 17502
rect 20414 17554 20466 17566
rect 20414 17490 20466 17502
rect 20526 17554 20578 17566
rect 20526 17490 20578 17502
rect 25342 17554 25394 17566
rect 29262 17554 29314 17566
rect 26338 17502 26350 17554
rect 26402 17502 26414 17554
rect 25342 17490 25394 17502
rect 29262 17490 29314 17502
rect 36542 17554 36594 17566
rect 36542 17490 36594 17502
rect 37550 17554 37602 17566
rect 37550 17490 37602 17502
rect 37886 17554 37938 17566
rect 37886 17490 37938 17502
rect 38222 17554 38274 17566
rect 38222 17490 38274 17502
rect 20190 17442 20242 17454
rect 22654 17442 22706 17454
rect 21298 17390 21310 17442
rect 21362 17390 21374 17442
rect 22306 17390 22318 17442
rect 22370 17390 22382 17442
rect 20190 17378 20242 17390
rect 22654 17378 22706 17390
rect 23886 17442 23938 17454
rect 37214 17442 37266 17454
rect 24210 17390 24222 17442
rect 24274 17390 24286 17442
rect 23886 17378 23938 17390
rect 37214 17378 37266 17390
rect 1344 17274 38800 17308
rect 1344 17222 10538 17274
rect 10590 17222 10642 17274
rect 10694 17222 10746 17274
rect 10798 17222 19862 17274
rect 19914 17222 19966 17274
rect 20018 17222 20070 17274
rect 20122 17222 29186 17274
rect 29238 17222 29290 17274
rect 29342 17222 29394 17274
rect 29446 17222 38510 17274
rect 38562 17222 38614 17274
rect 38666 17222 38718 17274
rect 38770 17222 38800 17274
rect 1344 17188 38800 17222
rect 2718 17106 2770 17118
rect 2718 17042 2770 17054
rect 18622 17106 18674 17118
rect 18622 17042 18674 17054
rect 19742 17106 19794 17118
rect 19742 17042 19794 17054
rect 20414 17106 20466 17118
rect 26898 17054 26910 17106
rect 26962 17054 26974 17106
rect 20414 17042 20466 17054
rect 2046 16994 2098 17006
rect 19070 16994 19122 17006
rect 16258 16942 16270 16994
rect 16322 16942 16334 16994
rect 2046 16930 2098 16942
rect 19070 16930 19122 16942
rect 20526 16994 20578 17006
rect 37550 16994 37602 17006
rect 22418 16942 22430 16994
rect 22482 16942 22494 16994
rect 20526 16930 20578 16942
rect 37550 16930 37602 16942
rect 37886 16994 37938 17006
rect 37886 16930 37938 16942
rect 1710 16882 1762 16894
rect 1710 16818 1762 16830
rect 2382 16882 2434 16894
rect 2382 16818 2434 16830
rect 3166 16882 3218 16894
rect 3166 16818 3218 16830
rect 12798 16882 12850 16894
rect 12798 16818 12850 16830
rect 13134 16882 13186 16894
rect 18062 16882 18114 16894
rect 14690 16830 14702 16882
rect 14754 16830 14766 16882
rect 15698 16830 15710 16882
rect 15762 16830 15774 16882
rect 13134 16818 13186 16830
rect 18062 16818 18114 16830
rect 19966 16882 20018 16894
rect 19966 16818 20018 16830
rect 20190 16882 20242 16894
rect 23102 16882 23154 16894
rect 37214 16882 37266 16894
rect 21858 16830 21870 16882
rect 21922 16830 21934 16882
rect 22306 16830 22318 16882
rect 22370 16830 22382 16882
rect 23650 16830 23662 16882
rect 23714 16830 23726 16882
rect 24546 16830 24558 16882
rect 24610 16830 24622 16882
rect 26226 16830 26238 16882
rect 26290 16830 26302 16882
rect 26786 16830 26798 16882
rect 26850 16830 26862 16882
rect 27458 16830 27470 16882
rect 27522 16830 27534 16882
rect 28130 16830 28142 16882
rect 28194 16830 28206 16882
rect 29026 16830 29038 16882
rect 29090 16830 29102 16882
rect 20190 16818 20242 16830
rect 23102 16818 23154 16830
rect 37214 16818 37266 16830
rect 38222 16882 38274 16894
rect 38222 16818 38274 16830
rect 19294 16770 19346 16782
rect 12450 16718 12462 16770
rect 12514 16718 12526 16770
rect 14578 16718 14590 16770
rect 14642 16718 14654 16770
rect 18946 16718 18958 16770
rect 19010 16718 19022 16770
rect 19294 16706 19346 16718
rect 21422 16770 21474 16782
rect 21422 16706 21474 16718
rect 25902 16770 25954 16782
rect 25902 16706 25954 16718
rect 19630 16658 19682 16670
rect 13906 16606 13918 16658
rect 13970 16606 13982 16658
rect 19630 16594 19682 16606
rect 1344 16490 38640 16524
rect 1344 16438 5876 16490
rect 5928 16438 5980 16490
rect 6032 16438 6084 16490
rect 6136 16438 15200 16490
rect 15252 16438 15304 16490
rect 15356 16438 15408 16490
rect 15460 16438 24524 16490
rect 24576 16438 24628 16490
rect 24680 16438 24732 16490
rect 24784 16438 33848 16490
rect 33900 16438 33952 16490
rect 34004 16438 34056 16490
rect 34108 16438 38640 16490
rect 1344 16404 38640 16438
rect 15586 16270 15598 16322
rect 15650 16270 15662 16322
rect 2494 16210 2546 16222
rect 14478 16210 14530 16222
rect 13794 16158 13806 16210
rect 13858 16158 13870 16210
rect 15362 16158 15374 16210
rect 15426 16158 15438 16210
rect 2494 16146 2546 16158
rect 14478 16146 14530 16158
rect 14142 16098 14194 16110
rect 17390 16098 17442 16110
rect 15138 16046 15150 16098
rect 15202 16046 15214 16098
rect 15810 16046 15822 16098
rect 15874 16046 15886 16098
rect 14142 16034 14194 16046
rect 17390 16034 17442 16046
rect 17950 16098 18002 16110
rect 17950 16034 18002 16046
rect 18174 16098 18226 16110
rect 18174 16034 18226 16046
rect 18510 16098 18562 16110
rect 18510 16034 18562 16046
rect 18846 16098 18898 16110
rect 19518 16098 19570 16110
rect 19170 16046 19182 16098
rect 19234 16046 19246 16098
rect 18846 16034 18898 16046
rect 19518 16034 19570 16046
rect 1710 15986 1762 15998
rect 1710 15922 1762 15934
rect 18398 15986 18450 15998
rect 18398 15922 18450 15934
rect 38222 15986 38274 15998
rect 38222 15922 38274 15934
rect 2046 15874 2098 15886
rect 2046 15810 2098 15822
rect 2942 15874 2994 15886
rect 2942 15810 2994 15822
rect 19294 15874 19346 15886
rect 19294 15810 19346 15822
rect 19406 15874 19458 15886
rect 19406 15810 19458 15822
rect 37662 15874 37714 15886
rect 37662 15810 37714 15822
rect 37886 15874 37938 15886
rect 37886 15810 37938 15822
rect 1344 15706 38800 15740
rect 1344 15654 10538 15706
rect 10590 15654 10642 15706
rect 10694 15654 10746 15706
rect 10798 15654 19862 15706
rect 19914 15654 19966 15706
rect 20018 15654 20070 15706
rect 20122 15654 29186 15706
rect 29238 15654 29290 15706
rect 29342 15654 29394 15706
rect 29446 15654 38510 15706
rect 38562 15654 38614 15706
rect 38666 15654 38718 15706
rect 38770 15654 38800 15706
rect 1344 15620 38800 15654
rect 19070 15538 19122 15550
rect 19070 15474 19122 15486
rect 21646 15538 21698 15550
rect 21646 15474 21698 15486
rect 2046 15426 2098 15438
rect 16382 15426 16434 15438
rect 37886 15426 37938 15438
rect 14578 15374 14590 15426
rect 14642 15374 14654 15426
rect 19506 15374 19518 15426
rect 19570 15374 19582 15426
rect 2046 15362 2098 15374
rect 16382 15362 16434 15374
rect 37886 15362 37938 15374
rect 1710 15314 1762 15326
rect 16046 15314 16098 15326
rect 14018 15262 14030 15314
rect 14082 15262 14094 15314
rect 14242 15262 14254 15314
rect 14306 15262 14318 15314
rect 15362 15262 15374 15314
rect 15426 15262 15438 15314
rect 1710 15250 1762 15262
rect 16046 15250 16098 15262
rect 18622 15314 18674 15326
rect 18622 15250 18674 15262
rect 18846 15314 18898 15326
rect 21198 15314 21250 15326
rect 20066 15262 20078 15314
rect 20130 15262 20142 15314
rect 20626 15262 20638 15314
rect 20690 15262 20702 15314
rect 18846 15250 18898 15262
rect 21198 15250 21250 15262
rect 21422 15314 21474 15326
rect 21422 15250 21474 15262
rect 21534 15314 21586 15326
rect 21534 15250 21586 15262
rect 38222 15314 38274 15326
rect 38222 15250 38274 15262
rect 2494 15202 2546 15214
rect 18958 15202 19010 15214
rect 37662 15202 37714 15214
rect 15698 15150 15710 15202
rect 15762 15150 15774 15202
rect 20178 15150 20190 15202
rect 20242 15150 20254 15202
rect 2494 15138 2546 15150
rect 18958 15138 19010 15150
rect 37662 15138 37714 15150
rect 18398 15090 18450 15102
rect 18398 15026 18450 15038
rect 20974 15090 21026 15102
rect 20974 15026 21026 15038
rect 1344 14922 38640 14956
rect 1344 14870 5876 14922
rect 5928 14870 5980 14922
rect 6032 14870 6084 14922
rect 6136 14870 15200 14922
rect 15252 14870 15304 14922
rect 15356 14870 15408 14922
rect 15460 14870 24524 14922
rect 24576 14870 24628 14922
rect 24680 14870 24732 14922
rect 24784 14870 33848 14922
rect 33900 14870 33952 14922
rect 34004 14870 34056 14922
rect 34108 14870 38640 14922
rect 1344 14836 38640 14870
rect 19506 14478 19518 14530
rect 19570 14478 19582 14530
rect 20626 14478 20638 14530
rect 20690 14478 20702 14530
rect 21298 14478 21310 14530
rect 21362 14478 21374 14530
rect 22194 14478 22206 14530
rect 22258 14478 22270 14530
rect 23202 14478 23214 14530
rect 23266 14478 23278 14530
rect 23650 14478 23662 14530
rect 23714 14478 23726 14530
rect 24994 14478 25006 14530
rect 25058 14478 25070 14530
rect 25890 14478 25902 14530
rect 25954 14478 25966 14530
rect 1710 14418 1762 14430
rect 1710 14354 1762 14366
rect 2046 14418 2098 14430
rect 22766 14418 22818 14430
rect 19954 14366 19966 14418
rect 20018 14366 20030 14418
rect 21410 14366 21422 14418
rect 21474 14366 21486 14418
rect 2046 14354 2098 14366
rect 22766 14354 22818 14366
rect 24222 14418 24274 14430
rect 24222 14354 24274 14366
rect 37662 14418 37714 14430
rect 37662 14354 37714 14366
rect 38222 14418 38274 14430
rect 38222 14354 38274 14366
rect 2494 14306 2546 14318
rect 37886 14306 37938 14318
rect 20402 14254 20414 14306
rect 20466 14254 20478 14306
rect 22306 14254 22318 14306
rect 22370 14254 22382 14306
rect 23762 14254 23774 14306
rect 23826 14254 23838 14306
rect 2494 14242 2546 14254
rect 37886 14242 37938 14254
rect 1344 14138 38800 14172
rect 1344 14086 10538 14138
rect 10590 14086 10642 14138
rect 10694 14086 10746 14138
rect 10798 14086 19862 14138
rect 19914 14086 19966 14138
rect 20018 14086 20070 14138
rect 20122 14086 29186 14138
rect 29238 14086 29290 14138
rect 29342 14086 29394 14138
rect 29446 14086 38510 14138
rect 38562 14086 38614 14138
rect 38666 14086 38718 14138
rect 38770 14086 38800 14138
rect 1344 14052 38800 14086
rect 2046 13970 2098 13982
rect 2046 13906 2098 13918
rect 17950 13970 18002 13982
rect 17950 13906 18002 13918
rect 18062 13970 18114 13982
rect 18062 13906 18114 13918
rect 37886 13970 37938 13982
rect 37886 13906 37938 13918
rect 2718 13858 2770 13870
rect 22878 13858 22930 13870
rect 20066 13806 20078 13858
rect 20130 13806 20142 13858
rect 22418 13806 22430 13858
rect 22482 13806 22494 13858
rect 2718 13794 2770 13806
rect 22878 13794 22930 13806
rect 1710 13746 1762 13758
rect 1710 13682 1762 13694
rect 2382 13746 2434 13758
rect 2382 13682 2434 13694
rect 17838 13746 17890 13758
rect 25454 13746 25506 13758
rect 19730 13694 19742 13746
rect 19794 13694 19806 13746
rect 21858 13694 21870 13746
rect 21922 13694 21934 13746
rect 22194 13694 22206 13746
rect 22258 13694 22270 13746
rect 23538 13694 23550 13746
rect 23602 13694 23614 13746
rect 24546 13694 24558 13746
rect 24610 13694 24622 13746
rect 17838 13682 17890 13694
rect 25454 13682 25506 13694
rect 38222 13746 38274 13758
rect 38222 13682 38274 13694
rect 3166 13634 3218 13646
rect 3166 13570 3218 13582
rect 3614 13634 3666 13646
rect 3614 13570 3666 13582
rect 18286 13634 18338 13646
rect 18286 13570 18338 13582
rect 18958 13634 19010 13646
rect 18958 13570 19010 13582
rect 21422 13634 21474 13646
rect 21422 13570 21474 13582
rect 37662 13634 37714 13646
rect 37662 13570 37714 13582
rect 18510 13522 18562 13534
rect 18510 13458 18562 13470
rect 19294 13522 19346 13534
rect 19294 13458 19346 13470
rect 1344 13354 38640 13388
rect 1344 13302 5876 13354
rect 5928 13302 5980 13354
rect 6032 13302 6084 13354
rect 6136 13302 15200 13354
rect 15252 13302 15304 13354
rect 15356 13302 15408 13354
rect 15460 13302 24524 13354
rect 24576 13302 24628 13354
rect 24680 13302 24732 13354
rect 24784 13302 33848 13354
rect 33900 13302 33952 13354
rect 34004 13302 34056 13354
rect 34108 13302 38640 13354
rect 1344 13268 38640 13302
rect 21310 13186 21362 13198
rect 21310 13122 21362 13134
rect 1934 13074 1986 13086
rect 1934 13010 1986 13022
rect 21870 13074 21922 13086
rect 21870 13010 21922 13022
rect 19294 12962 19346 12974
rect 21534 12962 21586 12974
rect 4274 12910 4286 12962
rect 4338 12910 4350 12962
rect 19730 12910 19742 12962
rect 19794 12910 19806 12962
rect 19294 12898 19346 12910
rect 21534 12898 21586 12910
rect 21982 12962 22034 12974
rect 24222 12962 24274 12974
rect 23202 12910 23214 12962
rect 23266 12910 23278 12962
rect 23650 12910 23662 12962
rect 23714 12910 23726 12962
rect 24994 12910 25006 12962
rect 25058 12910 25070 12962
rect 25890 12910 25902 12962
rect 25954 12910 25966 12962
rect 21982 12898 22034 12910
rect 24222 12898 24274 12910
rect 22766 12850 22818 12862
rect 20066 12798 20078 12850
rect 20130 12798 20142 12850
rect 22766 12786 22818 12798
rect 37214 12850 37266 12862
rect 37214 12786 37266 12798
rect 37550 12850 37602 12862
rect 37550 12786 37602 12798
rect 37886 12850 37938 12862
rect 37886 12786 37938 12798
rect 38222 12850 38274 12862
rect 38222 12786 38274 12798
rect 18958 12738 19010 12750
rect 18958 12674 19010 12686
rect 21758 12738 21810 12750
rect 36542 12738 36594 12750
rect 23762 12686 23774 12738
rect 23826 12686 23838 12738
rect 21758 12674 21810 12686
rect 36542 12674 36594 12686
rect 1344 12570 38800 12604
rect 1344 12518 10538 12570
rect 10590 12518 10642 12570
rect 10694 12518 10746 12570
rect 10798 12518 19862 12570
rect 19914 12518 19966 12570
rect 20018 12518 20070 12570
rect 20122 12518 29186 12570
rect 29238 12518 29290 12570
rect 29342 12518 29394 12570
rect 29446 12518 38510 12570
rect 38562 12518 38614 12570
rect 38666 12518 38718 12570
rect 38770 12518 38800 12570
rect 1344 12484 38800 12518
rect 18958 12402 19010 12414
rect 18958 12338 19010 12350
rect 20974 12402 21026 12414
rect 20974 12338 21026 12350
rect 21086 12402 21138 12414
rect 21086 12338 21138 12350
rect 21198 12402 21250 12414
rect 21198 12338 21250 12350
rect 37886 12290 37938 12302
rect 19842 12238 19854 12290
rect 19906 12238 19918 12290
rect 37886 12226 37938 12238
rect 20526 12178 20578 12190
rect 4274 12126 4286 12178
rect 4338 12126 4350 12178
rect 19730 12126 19742 12178
rect 19794 12126 19806 12178
rect 20526 12114 20578 12126
rect 20750 12178 20802 12190
rect 20750 12114 20802 12126
rect 37550 12178 37602 12190
rect 37550 12114 37602 12126
rect 38222 12178 38274 12190
rect 38222 12114 38274 12126
rect 37214 12066 37266 12078
rect 37214 12002 37266 12014
rect 1934 11954 1986 11966
rect 1934 11890 1986 11902
rect 19294 11954 19346 11966
rect 19294 11890 19346 11902
rect 1344 11786 38640 11820
rect 1344 11734 5876 11786
rect 5928 11734 5980 11786
rect 6032 11734 6084 11786
rect 6136 11734 15200 11786
rect 15252 11734 15304 11786
rect 15356 11734 15408 11786
rect 15460 11734 24524 11786
rect 24576 11734 24628 11786
rect 24680 11734 24732 11786
rect 24784 11734 33848 11786
rect 33900 11734 33952 11786
rect 34004 11734 34056 11786
rect 34108 11734 38640 11786
rect 1344 11700 38640 11734
rect 37886 11282 37938 11294
rect 37886 11218 37938 11230
rect 38222 11282 38274 11294
rect 38222 11218 38274 11230
rect 37662 11170 37714 11182
rect 37662 11106 37714 11118
rect 1344 11002 38800 11036
rect 1344 10950 10538 11002
rect 10590 10950 10642 11002
rect 10694 10950 10746 11002
rect 10798 10950 19862 11002
rect 19914 10950 19966 11002
rect 20018 10950 20070 11002
rect 20122 10950 29186 11002
rect 29238 10950 29290 11002
rect 29342 10950 29394 11002
rect 29446 10950 38510 11002
rect 38562 10950 38614 11002
rect 38666 10950 38718 11002
rect 38770 10950 38800 11002
rect 1344 10916 38800 10950
rect 37886 10722 37938 10734
rect 37886 10658 37938 10670
rect 37662 10610 37714 10622
rect 37662 10546 37714 10558
rect 38222 10610 38274 10622
rect 38222 10546 38274 10558
rect 1344 10218 38640 10252
rect 1344 10166 5876 10218
rect 5928 10166 5980 10218
rect 6032 10166 6084 10218
rect 6136 10166 15200 10218
rect 15252 10166 15304 10218
rect 15356 10166 15408 10218
rect 15460 10166 24524 10218
rect 24576 10166 24628 10218
rect 24680 10166 24732 10218
rect 24784 10166 33848 10218
rect 33900 10166 33952 10218
rect 34004 10166 34056 10218
rect 34108 10166 38640 10218
rect 1344 10132 38640 10166
rect 1344 9434 38800 9468
rect 1344 9382 10538 9434
rect 10590 9382 10642 9434
rect 10694 9382 10746 9434
rect 10798 9382 19862 9434
rect 19914 9382 19966 9434
rect 20018 9382 20070 9434
rect 20122 9382 29186 9434
rect 29238 9382 29290 9434
rect 29342 9382 29394 9434
rect 29446 9382 38510 9434
rect 38562 9382 38614 9434
rect 38666 9382 38718 9434
rect 38770 9382 38800 9434
rect 1344 9348 38800 9382
rect 1344 8650 38640 8684
rect 1344 8598 5876 8650
rect 5928 8598 5980 8650
rect 6032 8598 6084 8650
rect 6136 8598 15200 8650
rect 15252 8598 15304 8650
rect 15356 8598 15408 8650
rect 15460 8598 24524 8650
rect 24576 8598 24628 8650
rect 24680 8598 24732 8650
rect 24784 8598 33848 8650
rect 33900 8598 33952 8650
rect 34004 8598 34056 8650
rect 34108 8598 38640 8650
rect 1344 8564 38640 8598
rect 1344 7866 38800 7900
rect 1344 7814 10538 7866
rect 10590 7814 10642 7866
rect 10694 7814 10746 7866
rect 10798 7814 19862 7866
rect 19914 7814 19966 7866
rect 20018 7814 20070 7866
rect 20122 7814 29186 7866
rect 29238 7814 29290 7866
rect 29342 7814 29394 7866
rect 29446 7814 38510 7866
rect 38562 7814 38614 7866
rect 38666 7814 38718 7866
rect 38770 7814 38800 7866
rect 1344 7780 38800 7814
rect 1344 7082 38640 7116
rect 1344 7030 5876 7082
rect 5928 7030 5980 7082
rect 6032 7030 6084 7082
rect 6136 7030 15200 7082
rect 15252 7030 15304 7082
rect 15356 7030 15408 7082
rect 15460 7030 24524 7082
rect 24576 7030 24628 7082
rect 24680 7030 24732 7082
rect 24784 7030 33848 7082
rect 33900 7030 33952 7082
rect 34004 7030 34056 7082
rect 34108 7030 38640 7082
rect 1344 6996 38640 7030
rect 1344 6298 38800 6332
rect 1344 6246 10538 6298
rect 10590 6246 10642 6298
rect 10694 6246 10746 6298
rect 10798 6246 19862 6298
rect 19914 6246 19966 6298
rect 20018 6246 20070 6298
rect 20122 6246 29186 6298
rect 29238 6246 29290 6298
rect 29342 6246 29394 6298
rect 29446 6246 38510 6298
rect 38562 6246 38614 6298
rect 38666 6246 38718 6298
rect 38770 6246 38800 6298
rect 1344 6212 38800 6246
rect 1344 5514 38640 5548
rect 1344 5462 5876 5514
rect 5928 5462 5980 5514
rect 6032 5462 6084 5514
rect 6136 5462 15200 5514
rect 15252 5462 15304 5514
rect 15356 5462 15408 5514
rect 15460 5462 24524 5514
rect 24576 5462 24628 5514
rect 24680 5462 24732 5514
rect 24784 5462 33848 5514
rect 33900 5462 33952 5514
rect 34004 5462 34056 5514
rect 34108 5462 38640 5514
rect 1344 5428 38640 5462
rect 13694 5122 13746 5134
rect 13694 5058 13746 5070
rect 14366 5122 14418 5134
rect 14366 5058 14418 5070
rect 15038 5122 15090 5134
rect 15038 5058 15090 5070
rect 14702 5010 14754 5022
rect 14702 4946 14754 4958
rect 15374 5010 15426 5022
rect 15374 4946 15426 4958
rect 14142 4898 14194 4910
rect 14142 4834 14194 4846
rect 16606 4898 16658 4910
rect 16606 4834 16658 4846
rect 22206 4898 22258 4910
rect 22206 4834 22258 4846
rect 1344 4730 38800 4764
rect 1344 4678 10538 4730
rect 10590 4678 10642 4730
rect 10694 4678 10746 4730
rect 10798 4678 19862 4730
rect 19914 4678 19966 4730
rect 20018 4678 20070 4730
rect 20122 4678 29186 4730
rect 29238 4678 29290 4730
rect 29342 4678 29394 4730
rect 29446 4678 38510 4730
rect 38562 4678 38614 4730
rect 38666 4678 38718 4730
rect 38770 4678 38800 4730
rect 1344 4644 38800 4678
rect 16046 4562 16098 4574
rect 16046 4498 16098 4510
rect 21086 4562 21138 4574
rect 21086 4498 21138 4510
rect 21758 4562 21810 4574
rect 21758 4498 21810 4510
rect 22430 4562 22482 4574
rect 22430 4498 22482 4510
rect 27134 4562 27186 4574
rect 27134 4498 27186 4510
rect 29486 4562 29538 4574
rect 29486 4498 29538 4510
rect 15710 4338 15762 4350
rect 14914 4286 14926 4338
rect 14978 4286 14990 4338
rect 15710 4274 15762 4286
rect 20862 4338 20914 4350
rect 21298 4286 21310 4338
rect 21362 4286 21374 4338
rect 21970 4286 21982 4338
rect 22034 4286 22046 4338
rect 22642 4286 22654 4338
rect 22706 4286 22718 4338
rect 27346 4286 27358 4338
rect 27410 4286 27422 4338
rect 20862 4274 20914 4286
rect 15486 4226 15538 4238
rect 15486 4162 15538 4174
rect 16830 4226 16882 4238
rect 16830 4162 16882 4174
rect 17614 4226 17666 4238
rect 17614 4162 17666 4174
rect 18174 4226 18226 4238
rect 18174 4162 18226 4174
rect 18846 4226 18898 4238
rect 18846 4162 18898 4174
rect 19966 4226 20018 4238
rect 19966 4162 20018 4174
rect 20414 4226 20466 4238
rect 20414 4162 20466 4174
rect 23438 4226 23490 4238
rect 23438 4162 23490 4174
rect 24334 4226 24386 4238
rect 24334 4162 24386 4174
rect 25454 4226 25506 4238
rect 25454 4162 25506 4174
rect 25902 4226 25954 4238
rect 25902 4162 25954 4174
rect 26350 4226 26402 4238
rect 26350 4162 26402 4174
rect 26910 4226 26962 4238
rect 26910 4162 26962 4174
rect 27918 4226 27970 4238
rect 27918 4162 27970 4174
rect 28478 4226 28530 4238
rect 28478 4162 28530 4174
rect 28926 4226 28978 4238
rect 28926 4162 28978 4174
rect 30158 4226 30210 4238
rect 30158 4162 30210 4174
rect 30830 4226 30882 4238
rect 30830 4162 30882 4174
rect 12574 4114 12626 4126
rect 25554 4062 25566 4114
rect 25618 4111 25630 4114
rect 26338 4111 26350 4114
rect 25618 4065 26350 4111
rect 25618 4062 25630 4065
rect 26338 4062 26350 4065
rect 26402 4111 26414 4114
rect 26786 4111 26798 4114
rect 26402 4065 26798 4111
rect 26402 4062 26414 4065
rect 26786 4062 26798 4065
rect 26850 4062 26862 4114
rect 12574 4050 12626 4062
rect 1344 3946 38640 3980
rect 1344 3894 5876 3946
rect 5928 3894 5980 3946
rect 6032 3894 6084 3946
rect 6136 3894 15200 3946
rect 15252 3894 15304 3946
rect 15356 3894 15408 3946
rect 15460 3894 24524 3946
rect 24576 3894 24628 3946
rect 24680 3894 24732 3946
rect 24784 3894 33848 3946
rect 33900 3894 33952 3946
rect 34004 3894 34056 3946
rect 34108 3894 38640 3946
rect 1344 3860 38640 3894
rect 13358 3666 13410 3678
rect 13358 3602 13410 3614
rect 20974 3666 21026 3678
rect 20974 3602 21026 3614
rect 17054 3554 17106 3566
rect 12338 3502 12350 3554
rect 12402 3502 12414 3554
rect 15698 3502 15710 3554
rect 15762 3502 15774 3554
rect 16146 3502 16158 3554
rect 16210 3502 16222 3554
rect 17054 3490 17106 3502
rect 17726 3554 17778 3566
rect 26238 3554 26290 3566
rect 18610 3502 18622 3554
rect 18674 3502 18686 3554
rect 19282 3502 19294 3554
rect 19346 3502 19358 3554
rect 20066 3502 20078 3554
rect 20130 3502 20142 3554
rect 22866 3502 22878 3554
rect 22930 3502 22942 3554
rect 23874 3502 23886 3554
rect 23938 3502 23950 3554
rect 24770 3502 24782 3554
rect 24834 3502 24846 3554
rect 25442 3502 25454 3554
rect 25506 3502 25518 3554
rect 26786 3502 26798 3554
rect 26850 3502 26862 3554
rect 27458 3502 27470 3554
rect 27522 3502 27534 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 29922 3502 29934 3554
rect 29986 3502 29998 3554
rect 30594 3502 30606 3554
rect 30658 3502 30670 3554
rect 31266 3502 31278 3554
rect 31330 3502 31342 3554
rect 17726 3490 17778 3502
rect 26238 3490 26290 3502
rect 12014 3442 12066 3454
rect 12014 3378 12066 3390
rect 12574 3442 12626 3454
rect 12574 3378 12626 3390
rect 17390 3442 17442 3454
rect 17390 3378 17442 3390
rect 18062 3442 18114 3454
rect 18062 3378 18114 3390
rect 18398 3442 18450 3454
rect 18398 3378 18450 3390
rect 19070 3442 19122 3454
rect 19070 3378 19122 3390
rect 19854 3442 19906 3454
rect 19854 3378 19906 3390
rect 23662 3442 23714 3454
rect 23662 3378 23714 3390
rect 24558 3442 24610 3454
rect 24558 3378 24610 3390
rect 25230 3442 25282 3454
rect 25230 3378 25282 3390
rect 25902 3442 25954 3454
rect 25902 3378 25954 3390
rect 26574 3442 26626 3454
rect 26574 3378 26626 3390
rect 27246 3442 27298 3454
rect 27246 3378 27298 3390
rect 28366 3442 28418 3454
rect 28366 3378 28418 3390
rect 29374 3442 29426 3454
rect 29374 3378 29426 3390
rect 29710 3442 29762 3454
rect 29710 3378 29762 3390
rect 30382 3442 30434 3454
rect 30382 3378 30434 3390
rect 31054 3442 31106 3454
rect 31054 3378 31106 3390
rect 16382 3330 16434 3342
rect 16382 3266 16434 3278
rect 29038 3330 29090 3342
rect 29038 3266 29090 3278
rect 1344 3162 38800 3196
rect 1344 3110 10538 3162
rect 10590 3110 10642 3162
rect 10694 3110 10746 3162
rect 10798 3110 19862 3162
rect 19914 3110 19966 3162
rect 20018 3110 20070 3162
rect 20122 3110 29186 3162
rect 29238 3110 29290 3162
rect 29342 3110 29394 3162
rect 29446 3110 38510 3162
rect 38562 3110 38614 3162
rect 38666 3110 38718 3162
rect 38770 3110 38800 3162
rect 1344 3076 38800 3110
rect 28914 2830 28926 2882
rect 28978 2879 28990 2882
rect 29922 2879 29934 2882
rect 28978 2833 29934 2879
rect 28978 2830 28990 2833
rect 29922 2830 29934 2833
rect 29986 2830 29998 2882
<< via1 >>
rect 5876 36822 5928 36874
rect 5980 36822 6032 36874
rect 6084 36822 6136 36874
rect 15200 36822 15252 36874
rect 15304 36822 15356 36874
rect 15408 36822 15460 36874
rect 24524 36822 24576 36874
rect 24628 36822 24680 36874
rect 24732 36822 24784 36874
rect 33848 36822 33900 36874
rect 33952 36822 34004 36874
rect 34056 36822 34108 36874
rect 17166 36654 17218 36706
rect 22094 36654 22146 36706
rect 10222 36542 10274 36594
rect 28478 36542 28530 36594
rect 11006 36430 11058 36482
rect 11678 36430 11730 36482
rect 12350 36430 12402 36482
rect 13470 36430 13522 36482
rect 14142 36430 14194 36482
rect 14814 36430 14866 36482
rect 15486 36430 15538 36482
rect 16158 36430 16210 36482
rect 19182 36430 19234 36482
rect 19854 36430 19906 36482
rect 21086 36430 21138 36482
rect 24782 36430 24834 36482
rect 25454 36430 25506 36482
rect 26238 36430 26290 36482
rect 26798 36430 26850 36482
rect 27470 36430 27522 36482
rect 10670 36318 10722 36370
rect 11230 36206 11282 36258
rect 11902 36206 11954 36258
rect 12574 36206 12626 36258
rect 13694 36206 13746 36258
rect 14366 36206 14418 36258
rect 15038 36206 15090 36258
rect 15710 36206 15762 36258
rect 16382 36206 16434 36258
rect 20190 36206 20242 36258
rect 24558 36206 24610 36258
rect 25230 36206 25282 36258
rect 25902 36206 25954 36258
rect 26574 36206 26626 36258
rect 27246 36206 27298 36258
rect 10538 36038 10590 36090
rect 10642 36038 10694 36090
rect 10746 36038 10798 36090
rect 19862 36038 19914 36090
rect 19966 36038 20018 36090
rect 20070 36038 20122 36090
rect 29186 36038 29238 36090
rect 29290 36038 29342 36090
rect 29394 36038 29446 36090
rect 38510 36038 38562 36090
rect 38614 36038 38666 36090
rect 38718 36038 38770 36090
rect 14030 35870 14082 35922
rect 14590 35870 14642 35922
rect 15262 35870 15314 35922
rect 15934 35870 15986 35922
rect 16494 35870 16546 35922
rect 16942 35870 16994 35922
rect 19854 35870 19906 35922
rect 21422 35870 21474 35922
rect 25454 35870 25506 35922
rect 25902 35870 25954 35922
rect 26350 35870 26402 35922
rect 26910 35870 26962 35922
rect 17726 35758 17778 35810
rect 18062 35758 18114 35810
rect 18398 35758 18450 35810
rect 18734 35758 18786 35810
rect 19070 35758 19122 35810
rect 19406 35758 19458 35810
rect 23326 35758 23378 35810
rect 23998 35758 24050 35810
rect 27134 35758 27186 35810
rect 13358 35646 13410 35698
rect 20526 35646 20578 35698
rect 23550 35646 23602 35698
rect 24222 35646 24274 35698
rect 27358 35646 27410 35698
rect 11454 35534 11506 35586
rect 5876 35254 5928 35306
rect 5980 35254 6032 35306
rect 6084 35254 6136 35306
rect 15200 35254 15252 35306
rect 15304 35254 15356 35306
rect 15408 35254 15460 35306
rect 24524 35254 24576 35306
rect 24628 35254 24680 35306
rect 24732 35254 24784 35306
rect 33848 35254 33900 35306
rect 33952 35254 34004 35306
rect 34056 35254 34108 35306
rect 12798 34974 12850 35026
rect 18174 34974 18226 35026
rect 18846 34974 18898 35026
rect 21534 34974 21586 35026
rect 23102 34974 23154 35026
rect 23774 34974 23826 35026
rect 21758 34862 21810 34914
rect 22094 34638 22146 34690
rect 24334 34638 24386 34690
rect 10538 34470 10590 34522
rect 10642 34470 10694 34522
rect 10746 34470 10798 34522
rect 19862 34470 19914 34522
rect 19966 34470 20018 34522
rect 20070 34470 20122 34522
rect 29186 34470 29238 34522
rect 29290 34470 29342 34522
rect 29394 34470 29446 34522
rect 38510 34470 38562 34522
rect 38614 34470 38666 34522
rect 38718 34470 38770 34522
rect 5876 33686 5928 33738
rect 5980 33686 6032 33738
rect 6084 33686 6136 33738
rect 15200 33686 15252 33738
rect 15304 33686 15356 33738
rect 15408 33686 15460 33738
rect 24524 33686 24576 33738
rect 24628 33686 24680 33738
rect 24732 33686 24784 33738
rect 33848 33686 33900 33738
rect 33952 33686 34004 33738
rect 34056 33686 34108 33738
rect 10538 32902 10590 32954
rect 10642 32902 10694 32954
rect 10746 32902 10798 32954
rect 19862 32902 19914 32954
rect 19966 32902 20018 32954
rect 20070 32902 20122 32954
rect 29186 32902 29238 32954
rect 29290 32902 29342 32954
rect 29394 32902 29446 32954
rect 38510 32902 38562 32954
rect 38614 32902 38666 32954
rect 38718 32902 38770 32954
rect 5876 32118 5928 32170
rect 5980 32118 6032 32170
rect 6084 32118 6136 32170
rect 15200 32118 15252 32170
rect 15304 32118 15356 32170
rect 15408 32118 15460 32170
rect 24524 32118 24576 32170
rect 24628 32118 24680 32170
rect 24732 32118 24784 32170
rect 33848 32118 33900 32170
rect 33952 32118 34004 32170
rect 34056 32118 34108 32170
rect 10538 31334 10590 31386
rect 10642 31334 10694 31386
rect 10746 31334 10798 31386
rect 19862 31334 19914 31386
rect 19966 31334 20018 31386
rect 20070 31334 20122 31386
rect 29186 31334 29238 31386
rect 29290 31334 29342 31386
rect 29394 31334 29446 31386
rect 38510 31334 38562 31386
rect 38614 31334 38666 31386
rect 38718 31334 38770 31386
rect 37886 31054 37938 31106
rect 38222 30942 38274 30994
rect 37662 30830 37714 30882
rect 5876 30550 5928 30602
rect 5980 30550 6032 30602
rect 6084 30550 6136 30602
rect 15200 30550 15252 30602
rect 15304 30550 15356 30602
rect 15408 30550 15460 30602
rect 24524 30550 24576 30602
rect 24628 30550 24680 30602
rect 24732 30550 24784 30602
rect 33848 30550 33900 30602
rect 33952 30550 34004 30602
rect 34056 30550 34108 30602
rect 37662 30046 37714 30098
rect 38222 30046 38274 30098
rect 37886 29934 37938 29986
rect 10538 29766 10590 29818
rect 10642 29766 10694 29818
rect 10746 29766 10798 29818
rect 19862 29766 19914 29818
rect 19966 29766 20018 29818
rect 20070 29766 20122 29818
rect 29186 29766 29238 29818
rect 29290 29766 29342 29818
rect 29394 29766 29446 29818
rect 38510 29766 38562 29818
rect 38614 29766 38666 29818
rect 38718 29766 38770 29818
rect 37886 29486 37938 29538
rect 4286 29374 4338 29426
rect 38222 29374 38274 29426
rect 37662 29262 37714 29314
rect 1934 29150 1986 29202
rect 5876 28982 5928 29034
rect 5980 28982 6032 29034
rect 6084 28982 6136 29034
rect 15200 28982 15252 29034
rect 15304 28982 15356 29034
rect 15408 28982 15460 29034
rect 24524 28982 24576 29034
rect 24628 28982 24680 29034
rect 24732 28982 24784 29034
rect 33848 28982 33900 29034
rect 33952 28982 34004 29034
rect 34056 28982 34108 29034
rect 1710 28590 1762 28642
rect 2494 28590 2546 28642
rect 37662 28590 37714 28642
rect 38110 28590 38162 28642
rect 37886 28478 37938 28530
rect 2046 28366 2098 28418
rect 10538 28198 10590 28250
rect 10642 28198 10694 28250
rect 10746 28198 10798 28250
rect 19862 28198 19914 28250
rect 19966 28198 20018 28250
rect 20070 28198 20122 28250
rect 29186 28198 29238 28250
rect 29290 28198 29342 28250
rect 29394 28198 29446 28250
rect 38510 28198 38562 28250
rect 38614 28198 38666 28250
rect 38718 28198 38770 28250
rect 20526 28030 20578 28082
rect 2046 27918 2098 27970
rect 19854 27918 19906 27970
rect 20302 27918 20354 27970
rect 37886 27918 37938 27970
rect 1710 27806 1762 27858
rect 19518 27806 19570 27858
rect 38222 27806 38274 27858
rect 2494 27694 2546 27746
rect 2942 27694 2994 27746
rect 37214 27694 37266 27746
rect 37662 27694 37714 27746
rect 5876 27414 5928 27466
rect 5980 27414 6032 27466
rect 6084 27414 6136 27466
rect 15200 27414 15252 27466
rect 15304 27414 15356 27466
rect 15408 27414 15460 27466
rect 24524 27414 24576 27466
rect 24628 27414 24680 27466
rect 24732 27414 24784 27466
rect 33848 27414 33900 27466
rect 33952 27414 34004 27466
rect 34056 27414 34108 27466
rect 19854 27246 19906 27298
rect 17502 27134 17554 27186
rect 1822 27022 1874 27074
rect 16270 27022 16322 27074
rect 16494 27022 16546 27074
rect 17614 27022 17666 27074
rect 18734 27022 18786 27074
rect 19742 27022 19794 27074
rect 20190 27022 20242 27074
rect 20638 27022 20690 27074
rect 37662 27022 37714 27074
rect 38110 27022 38162 27074
rect 2046 26910 2098 26962
rect 2382 26910 2434 26962
rect 3166 26910 3218 26962
rect 17054 26910 17106 26962
rect 18174 26910 18226 26962
rect 18510 26910 18562 26962
rect 21310 26910 21362 26962
rect 21646 26910 21698 26962
rect 37326 26910 37378 26962
rect 2718 26798 2770 26850
rect 21534 26798 21586 26850
rect 36990 26798 37042 26850
rect 10538 26630 10590 26682
rect 10642 26630 10694 26682
rect 10746 26630 10798 26682
rect 19862 26630 19914 26682
rect 19966 26630 20018 26682
rect 20070 26630 20122 26682
rect 29186 26630 29238 26682
rect 29290 26630 29342 26682
rect 29394 26630 29446 26682
rect 38510 26630 38562 26682
rect 38614 26630 38666 26682
rect 38718 26630 38770 26682
rect 15038 26462 15090 26514
rect 17726 26462 17778 26514
rect 37662 26462 37714 26514
rect 2046 26350 2098 26402
rect 14814 26350 14866 26402
rect 37886 26350 37938 26402
rect 1710 26238 1762 26290
rect 14702 26238 14754 26290
rect 15598 26238 15650 26290
rect 16606 26238 16658 26290
rect 18510 26238 18562 26290
rect 19518 26238 19570 26290
rect 20302 26238 20354 26290
rect 20974 26238 21026 26290
rect 38222 26238 38274 26290
rect 2494 26126 2546 26178
rect 15822 26126 15874 26178
rect 16382 26126 16434 26178
rect 21422 26126 21474 26178
rect 37214 26126 37266 26178
rect 19630 26014 19682 26066
rect 5876 25846 5928 25898
rect 5980 25846 6032 25898
rect 6084 25846 6136 25898
rect 15200 25846 15252 25898
rect 15304 25846 15356 25898
rect 15408 25846 15460 25898
rect 24524 25846 24576 25898
rect 24628 25846 24680 25898
rect 24732 25846 24784 25898
rect 33848 25846 33900 25898
rect 33952 25846 34004 25898
rect 34056 25846 34108 25898
rect 14366 25678 14418 25730
rect 14702 25678 14754 25730
rect 15710 25566 15762 25618
rect 16494 25566 16546 25618
rect 19182 25566 19234 25618
rect 21870 25566 21922 25618
rect 13694 25454 13746 25506
rect 15598 25454 15650 25506
rect 16606 25454 16658 25506
rect 17390 25454 17442 25506
rect 18622 25454 18674 25506
rect 19630 25454 19682 25506
rect 22206 25454 22258 25506
rect 22654 25454 22706 25506
rect 23438 25454 23490 25506
rect 23998 25454 24050 25506
rect 24894 25454 24946 25506
rect 1710 25342 1762 25394
rect 13582 25342 13634 25394
rect 20078 25342 20130 25394
rect 21422 25342 21474 25394
rect 21534 25342 21586 25394
rect 22878 25342 22930 25394
rect 37662 25342 37714 25394
rect 38222 25342 38274 25394
rect 2046 25230 2098 25282
rect 2494 25230 2546 25282
rect 21198 25230 21250 25282
rect 37886 25230 37938 25282
rect 10538 25062 10590 25114
rect 10642 25062 10694 25114
rect 10746 25062 10798 25114
rect 19862 25062 19914 25114
rect 19966 25062 20018 25114
rect 20070 25062 20122 25114
rect 29186 25062 29238 25114
rect 29290 25062 29342 25114
rect 29394 25062 29446 25114
rect 38510 25062 38562 25114
rect 38614 25062 38666 25114
rect 38718 25062 38770 25114
rect 22878 24894 22930 24946
rect 2046 24782 2098 24834
rect 16270 24782 16322 24834
rect 22654 24782 22706 24834
rect 22990 24782 23042 24834
rect 26574 24782 26626 24834
rect 37886 24782 37938 24834
rect 1710 24670 1762 24722
rect 12350 24670 12402 24722
rect 12574 24670 12626 24722
rect 13134 24670 13186 24722
rect 14702 24670 14754 24722
rect 15710 24670 15762 24722
rect 17950 24670 18002 24722
rect 18734 24670 18786 24722
rect 20302 24670 20354 24722
rect 20974 24670 21026 24722
rect 25902 24670 25954 24722
rect 26462 24670 26514 24722
rect 27022 24670 27074 24722
rect 27806 24670 27858 24722
rect 28702 24670 28754 24722
rect 38222 24670 38274 24722
rect 2494 24558 2546 24610
rect 14590 24558 14642 24610
rect 21758 24558 21810 24610
rect 25566 24558 25618 24610
rect 37662 24558 37714 24610
rect 15822 24446 15874 24498
rect 19630 24446 19682 24498
rect 5876 24278 5928 24330
rect 5980 24278 6032 24330
rect 6084 24278 6136 24330
rect 15200 24278 15252 24330
rect 15304 24278 15356 24330
rect 15408 24278 15460 24330
rect 24524 24278 24576 24330
rect 24628 24278 24680 24330
rect 24732 24278 24784 24330
rect 33848 24278 33900 24330
rect 33952 24278 34004 24330
rect 34056 24278 34108 24330
rect 14590 24110 14642 24162
rect 17838 24110 17890 24162
rect 12462 23998 12514 24050
rect 16718 23998 16770 24050
rect 21870 23998 21922 24050
rect 14366 23886 14418 23938
rect 14702 23886 14754 23938
rect 15598 23886 15650 23938
rect 17502 23886 17554 23938
rect 18622 23886 18674 23938
rect 19630 23886 19682 23938
rect 21198 23886 21250 23938
rect 22206 23886 22258 23938
rect 22766 23886 22818 23938
rect 23438 23886 23490 23938
rect 24110 23886 24162 23938
rect 25006 23886 25058 23938
rect 20078 23774 20130 23826
rect 21422 23774 21474 23826
rect 21534 23774 21586 23826
rect 38222 23774 38274 23826
rect 1710 23662 1762 23714
rect 2046 23662 2098 23714
rect 2494 23662 2546 23714
rect 12910 23662 12962 23714
rect 13918 23662 13970 23714
rect 16270 23662 16322 23714
rect 22878 23662 22930 23714
rect 37662 23662 37714 23714
rect 37886 23662 37938 23714
rect 10538 23494 10590 23546
rect 10642 23494 10694 23546
rect 10746 23494 10798 23546
rect 19862 23494 19914 23546
rect 19966 23494 20018 23546
rect 20070 23494 20122 23546
rect 29186 23494 29238 23546
rect 29290 23494 29342 23546
rect 29394 23494 29446 23546
rect 38510 23494 38562 23546
rect 38614 23494 38666 23546
rect 38718 23494 38770 23546
rect 21422 23326 21474 23378
rect 26462 23326 26514 23378
rect 2046 23214 2098 23266
rect 16718 23214 16770 23266
rect 18622 23214 18674 23266
rect 23550 23214 23602 23266
rect 37886 23214 37938 23266
rect 1710 23102 1762 23154
rect 13582 23102 13634 23154
rect 15038 23102 15090 23154
rect 15598 23102 15650 23154
rect 17390 23102 17442 23154
rect 17838 23102 17890 23154
rect 19182 23102 19234 23154
rect 19742 23102 19794 23154
rect 20078 23102 20130 23154
rect 20414 23102 20466 23154
rect 21086 23102 21138 23154
rect 23326 23102 23378 23154
rect 25790 23102 25842 23154
rect 26350 23102 26402 23154
rect 27022 23102 27074 23154
rect 27694 23102 27746 23154
rect 28478 23102 28530 23154
rect 38222 23102 38274 23154
rect 2494 22990 2546 23042
rect 13134 22990 13186 23042
rect 14478 22990 14530 23042
rect 25454 22990 25506 23042
rect 37662 22990 37714 23042
rect 20190 22878 20242 22930
rect 5876 22710 5928 22762
rect 5980 22710 6032 22762
rect 6084 22710 6136 22762
rect 15200 22710 15252 22762
rect 15304 22710 15356 22762
rect 15408 22710 15460 22762
rect 24524 22710 24576 22762
rect 24628 22710 24680 22762
rect 24732 22710 24784 22762
rect 33848 22710 33900 22762
rect 33952 22710 34004 22762
rect 34056 22710 34108 22762
rect 20414 22542 20466 22594
rect 20862 22542 20914 22594
rect 15598 22430 15650 22482
rect 17726 22430 17778 22482
rect 20078 22430 20130 22482
rect 13806 22318 13858 22370
rect 15934 22318 15986 22370
rect 16830 22318 16882 22370
rect 17614 22318 17666 22370
rect 18510 22318 18562 22370
rect 19630 22318 19682 22370
rect 1710 22206 1762 22258
rect 2046 22206 2098 22258
rect 21534 22206 21586 22258
rect 21870 22206 21922 22258
rect 21982 22206 22034 22258
rect 36542 22206 36594 22258
rect 37550 22206 37602 22258
rect 38222 22206 38274 22258
rect 2382 22094 2434 22146
rect 2718 22094 2770 22146
rect 3166 22094 3218 22146
rect 14478 22094 14530 22146
rect 20638 22094 20690 22146
rect 21198 22094 21250 22146
rect 21422 22094 21474 22146
rect 22206 22094 22258 22146
rect 23438 22094 23490 22146
rect 24222 22094 24274 22146
rect 37214 22094 37266 22146
rect 37886 22094 37938 22146
rect 10538 21926 10590 21978
rect 10642 21926 10694 21978
rect 10746 21926 10798 21978
rect 19862 21926 19914 21978
rect 19966 21926 20018 21978
rect 20070 21926 20122 21978
rect 29186 21926 29238 21978
rect 29290 21926 29342 21978
rect 29394 21926 29446 21978
rect 38510 21926 38562 21978
rect 38614 21926 38666 21978
rect 38718 21926 38770 21978
rect 2494 21758 2546 21810
rect 17390 21758 17442 21810
rect 2046 21646 2098 21698
rect 19742 21646 19794 21698
rect 20414 21646 20466 21698
rect 21086 21646 21138 21698
rect 23998 21646 24050 21698
rect 37886 21646 37938 21698
rect 1710 21534 1762 21586
rect 12350 21534 12402 21586
rect 13582 21534 13634 21586
rect 14926 21534 14978 21586
rect 15374 21534 15426 21586
rect 19518 21534 19570 21586
rect 20526 21534 20578 21586
rect 21422 21534 21474 21586
rect 22094 21534 22146 21586
rect 23774 21534 23826 21586
rect 25230 21534 25282 21586
rect 25790 21534 25842 21586
rect 37550 21534 37602 21586
rect 38222 21534 38274 21586
rect 2942 21422 2994 21474
rect 12126 21422 12178 21474
rect 15822 21422 15874 21474
rect 17950 21422 18002 21474
rect 18510 21422 18562 21474
rect 20302 21422 20354 21474
rect 22878 21422 22930 21474
rect 23214 21422 23266 21474
rect 24446 21422 24498 21474
rect 37214 21422 37266 21474
rect 15710 21310 15762 21362
rect 24334 21310 24386 21362
rect 5876 21142 5928 21194
rect 5980 21142 6032 21194
rect 6084 21142 6136 21194
rect 15200 21142 15252 21194
rect 15304 21142 15356 21194
rect 15408 21142 15460 21194
rect 24524 21142 24576 21194
rect 24628 21142 24680 21194
rect 24732 21142 24784 21194
rect 33848 21142 33900 21194
rect 33952 21142 34004 21194
rect 34056 21142 34108 21194
rect 17390 20974 17442 21026
rect 20638 20974 20690 21026
rect 12462 20862 12514 20914
rect 16942 20862 16994 20914
rect 28254 20862 28306 20914
rect 11342 20750 11394 20802
rect 12910 20750 12962 20802
rect 13470 20750 13522 20802
rect 13806 20750 13858 20802
rect 15374 20750 15426 20802
rect 16830 20750 16882 20802
rect 18958 20750 19010 20802
rect 20078 20750 20130 20802
rect 20190 20750 20242 20802
rect 20526 20750 20578 20802
rect 21310 20750 21362 20802
rect 22318 20750 22370 20802
rect 23438 20750 23490 20802
rect 24334 20750 24386 20802
rect 24894 20750 24946 20802
rect 25566 20750 25618 20802
rect 26238 20750 26290 20802
rect 27134 20750 27186 20802
rect 11790 20638 11842 20690
rect 18286 20638 18338 20690
rect 22542 20638 22594 20690
rect 23102 20638 23154 20690
rect 23998 20638 24050 20690
rect 27806 20638 27858 20690
rect 38222 20638 38274 20690
rect 1710 20526 1762 20578
rect 2046 20526 2098 20578
rect 2494 20526 2546 20578
rect 18622 20526 18674 20578
rect 21198 20526 21250 20578
rect 25006 20526 25058 20578
rect 37662 20526 37714 20578
rect 37886 20526 37938 20578
rect 10538 20358 10590 20410
rect 10642 20358 10694 20410
rect 10746 20358 10798 20410
rect 19862 20358 19914 20410
rect 19966 20358 20018 20410
rect 20070 20358 20122 20410
rect 29186 20358 29238 20410
rect 29290 20358 29342 20410
rect 29394 20358 29446 20410
rect 38510 20358 38562 20410
rect 38614 20358 38666 20410
rect 38718 20358 38770 20410
rect 22094 20190 22146 20242
rect 25790 20190 25842 20242
rect 2046 20078 2098 20130
rect 18174 20078 18226 20130
rect 21310 20078 21362 20130
rect 21758 20078 21810 20130
rect 22542 20078 22594 20130
rect 23214 20078 23266 20130
rect 24670 20078 24722 20130
rect 37886 20078 37938 20130
rect 1710 19966 1762 20018
rect 12350 19966 12402 20018
rect 13582 19966 13634 20018
rect 14926 19966 14978 20018
rect 15374 19966 15426 20018
rect 17614 19966 17666 20018
rect 19294 19966 19346 20018
rect 21534 19966 21586 20018
rect 21646 19966 21698 20018
rect 22654 19966 22706 20018
rect 22766 19966 22818 20018
rect 23438 19966 23490 20018
rect 23774 19966 23826 20018
rect 24446 19966 24498 20018
rect 26910 19966 26962 20018
rect 27470 19966 27522 20018
rect 28814 19966 28866 20018
rect 29934 19966 29986 20018
rect 38222 19966 38274 20018
rect 2494 19854 2546 19906
rect 15822 19854 15874 19906
rect 19182 19854 19234 19906
rect 25230 19854 25282 19906
rect 26238 19854 26290 19906
rect 26574 19854 26626 19906
rect 27694 19854 27746 19906
rect 37662 19854 37714 19906
rect 15710 19742 15762 19794
rect 18734 19742 18786 19794
rect 23102 19742 23154 19794
rect 28478 19742 28530 19794
rect 5876 19574 5928 19626
rect 5980 19574 6032 19626
rect 6084 19574 6136 19626
rect 15200 19574 15252 19626
rect 15304 19574 15356 19626
rect 15408 19574 15460 19626
rect 24524 19574 24576 19626
rect 24628 19574 24680 19626
rect 24732 19574 24784 19626
rect 33848 19574 33900 19626
rect 33952 19574 34004 19626
rect 34056 19574 34108 19626
rect 18958 19406 19010 19458
rect 1934 19294 1986 19346
rect 12238 19294 12290 19346
rect 12910 19294 12962 19346
rect 15598 19294 15650 19346
rect 17054 19294 17106 19346
rect 25342 19294 25394 19346
rect 4286 19182 4338 19234
rect 12574 19182 12626 19234
rect 13470 19182 13522 19234
rect 13806 19182 13858 19234
rect 15374 19182 15426 19234
rect 16830 19182 16882 19234
rect 18174 19182 18226 19234
rect 19406 19182 19458 19234
rect 19630 19182 19682 19234
rect 20302 19182 20354 19234
rect 21646 19182 21698 19234
rect 21982 19182 22034 19234
rect 25790 19182 25842 19234
rect 26238 19182 26290 19234
rect 26910 19182 26962 19234
rect 27582 19182 27634 19234
rect 28478 19182 28530 19234
rect 18510 19070 18562 19122
rect 19966 19070 20018 19122
rect 21870 19070 21922 19122
rect 26350 19070 26402 19122
rect 37886 19070 37938 19122
rect 38222 19070 38274 19122
rect 18398 18958 18450 19010
rect 37662 18958 37714 19010
rect 10538 18790 10590 18842
rect 10642 18790 10694 18842
rect 10746 18790 10798 18842
rect 19862 18790 19914 18842
rect 19966 18790 20018 18842
rect 20070 18790 20122 18842
rect 29186 18790 29238 18842
rect 29290 18790 29342 18842
rect 29394 18790 29446 18842
rect 38510 18790 38562 18842
rect 38614 18790 38666 18842
rect 38718 18790 38770 18842
rect 37886 18622 37938 18674
rect 2046 18510 2098 18562
rect 16270 18510 16322 18562
rect 22206 18510 22258 18562
rect 1710 18398 1762 18450
rect 13470 18398 13522 18450
rect 14702 18398 14754 18450
rect 15598 18398 15650 18450
rect 17950 18398 18002 18450
rect 18958 18398 19010 18450
rect 19742 18398 19794 18450
rect 20414 18398 20466 18450
rect 21534 18398 21586 18450
rect 22542 18398 22594 18450
rect 22878 18398 22930 18450
rect 25230 18398 25282 18450
rect 38222 18398 38274 18450
rect 2494 18286 2546 18338
rect 17390 18286 17442 18338
rect 18398 18286 18450 18338
rect 19294 18286 19346 18338
rect 21086 18286 21138 18338
rect 22990 18286 23042 18338
rect 25790 18286 25842 18338
rect 37662 18286 37714 18338
rect 15934 18174 15986 18226
rect 5876 18006 5928 18058
rect 5980 18006 6032 18058
rect 6084 18006 6136 18058
rect 15200 18006 15252 18058
rect 15304 18006 15356 18058
rect 15408 18006 15460 18058
rect 24524 18006 24576 18058
rect 24628 18006 24680 18058
rect 24732 18006 24784 18058
rect 33848 18006 33900 18058
rect 33952 18006 34004 18058
rect 34056 18006 34108 18058
rect 12798 17838 12850 17890
rect 16830 17838 16882 17890
rect 1934 17726 1986 17778
rect 11790 17726 11842 17778
rect 14814 17726 14866 17778
rect 4286 17614 4338 17666
rect 12238 17614 12290 17666
rect 13022 17614 13074 17666
rect 13806 17614 13858 17666
rect 14030 17614 14082 17666
rect 14926 17614 14978 17666
rect 15486 17614 15538 17666
rect 16606 17614 16658 17666
rect 17726 17614 17778 17666
rect 19406 17614 19458 17666
rect 19630 17614 19682 17666
rect 19966 17614 20018 17666
rect 21646 17614 21698 17666
rect 22990 17614 23042 17666
rect 23438 17614 23490 17666
rect 25790 17614 25842 17666
rect 26238 17614 26290 17666
rect 26910 17614 26962 17666
rect 27358 17614 27410 17666
rect 28478 17614 28530 17666
rect 18174 17502 18226 17554
rect 19070 17502 19122 17554
rect 19854 17502 19906 17554
rect 20414 17502 20466 17554
rect 20526 17502 20578 17554
rect 25342 17502 25394 17554
rect 26350 17502 26402 17554
rect 29262 17502 29314 17554
rect 36542 17502 36594 17554
rect 37550 17502 37602 17554
rect 37886 17502 37938 17554
rect 38222 17502 38274 17554
rect 20190 17390 20242 17442
rect 21310 17390 21362 17442
rect 22318 17390 22370 17442
rect 22654 17390 22706 17442
rect 23886 17390 23938 17442
rect 24222 17390 24274 17442
rect 37214 17390 37266 17442
rect 10538 17222 10590 17274
rect 10642 17222 10694 17274
rect 10746 17222 10798 17274
rect 19862 17222 19914 17274
rect 19966 17222 20018 17274
rect 20070 17222 20122 17274
rect 29186 17222 29238 17274
rect 29290 17222 29342 17274
rect 29394 17222 29446 17274
rect 38510 17222 38562 17274
rect 38614 17222 38666 17274
rect 38718 17222 38770 17274
rect 2718 17054 2770 17106
rect 18622 17054 18674 17106
rect 19742 17054 19794 17106
rect 20414 17054 20466 17106
rect 26910 17054 26962 17106
rect 2046 16942 2098 16994
rect 16270 16942 16322 16994
rect 19070 16942 19122 16994
rect 20526 16942 20578 16994
rect 22430 16942 22482 16994
rect 37550 16942 37602 16994
rect 37886 16942 37938 16994
rect 1710 16830 1762 16882
rect 2382 16830 2434 16882
rect 3166 16830 3218 16882
rect 12798 16830 12850 16882
rect 13134 16830 13186 16882
rect 14702 16830 14754 16882
rect 15710 16830 15762 16882
rect 18062 16830 18114 16882
rect 19966 16830 20018 16882
rect 20190 16830 20242 16882
rect 21870 16830 21922 16882
rect 22318 16830 22370 16882
rect 23102 16830 23154 16882
rect 23662 16830 23714 16882
rect 24558 16830 24610 16882
rect 26238 16830 26290 16882
rect 26798 16830 26850 16882
rect 27470 16830 27522 16882
rect 28142 16830 28194 16882
rect 29038 16830 29090 16882
rect 37214 16830 37266 16882
rect 38222 16830 38274 16882
rect 12462 16718 12514 16770
rect 14590 16718 14642 16770
rect 18958 16718 19010 16770
rect 19294 16718 19346 16770
rect 21422 16718 21474 16770
rect 25902 16718 25954 16770
rect 13918 16606 13970 16658
rect 19630 16606 19682 16658
rect 5876 16438 5928 16490
rect 5980 16438 6032 16490
rect 6084 16438 6136 16490
rect 15200 16438 15252 16490
rect 15304 16438 15356 16490
rect 15408 16438 15460 16490
rect 24524 16438 24576 16490
rect 24628 16438 24680 16490
rect 24732 16438 24784 16490
rect 33848 16438 33900 16490
rect 33952 16438 34004 16490
rect 34056 16438 34108 16490
rect 15598 16270 15650 16322
rect 2494 16158 2546 16210
rect 13806 16158 13858 16210
rect 14478 16158 14530 16210
rect 15374 16158 15426 16210
rect 14142 16046 14194 16098
rect 15150 16046 15202 16098
rect 15822 16046 15874 16098
rect 17390 16046 17442 16098
rect 17950 16046 18002 16098
rect 18174 16046 18226 16098
rect 18510 16046 18562 16098
rect 18846 16046 18898 16098
rect 19182 16046 19234 16098
rect 19518 16046 19570 16098
rect 1710 15934 1762 15986
rect 18398 15934 18450 15986
rect 38222 15934 38274 15986
rect 2046 15822 2098 15874
rect 2942 15822 2994 15874
rect 19294 15822 19346 15874
rect 19406 15822 19458 15874
rect 37662 15822 37714 15874
rect 37886 15822 37938 15874
rect 10538 15654 10590 15706
rect 10642 15654 10694 15706
rect 10746 15654 10798 15706
rect 19862 15654 19914 15706
rect 19966 15654 20018 15706
rect 20070 15654 20122 15706
rect 29186 15654 29238 15706
rect 29290 15654 29342 15706
rect 29394 15654 29446 15706
rect 38510 15654 38562 15706
rect 38614 15654 38666 15706
rect 38718 15654 38770 15706
rect 19070 15486 19122 15538
rect 21646 15486 21698 15538
rect 2046 15374 2098 15426
rect 14590 15374 14642 15426
rect 16382 15374 16434 15426
rect 19518 15374 19570 15426
rect 37886 15374 37938 15426
rect 1710 15262 1762 15314
rect 14030 15262 14082 15314
rect 14254 15262 14306 15314
rect 15374 15262 15426 15314
rect 16046 15262 16098 15314
rect 18622 15262 18674 15314
rect 18846 15262 18898 15314
rect 20078 15262 20130 15314
rect 20638 15262 20690 15314
rect 21198 15262 21250 15314
rect 21422 15262 21474 15314
rect 21534 15262 21586 15314
rect 38222 15262 38274 15314
rect 2494 15150 2546 15202
rect 15710 15150 15762 15202
rect 18958 15150 19010 15202
rect 20190 15150 20242 15202
rect 37662 15150 37714 15202
rect 18398 15038 18450 15090
rect 20974 15038 21026 15090
rect 5876 14870 5928 14922
rect 5980 14870 6032 14922
rect 6084 14870 6136 14922
rect 15200 14870 15252 14922
rect 15304 14870 15356 14922
rect 15408 14870 15460 14922
rect 24524 14870 24576 14922
rect 24628 14870 24680 14922
rect 24732 14870 24784 14922
rect 33848 14870 33900 14922
rect 33952 14870 34004 14922
rect 34056 14870 34108 14922
rect 19518 14478 19570 14530
rect 20638 14478 20690 14530
rect 21310 14478 21362 14530
rect 22206 14478 22258 14530
rect 23214 14478 23266 14530
rect 23662 14478 23714 14530
rect 25006 14478 25058 14530
rect 25902 14478 25954 14530
rect 1710 14366 1762 14418
rect 2046 14366 2098 14418
rect 19966 14366 20018 14418
rect 21422 14366 21474 14418
rect 22766 14366 22818 14418
rect 24222 14366 24274 14418
rect 37662 14366 37714 14418
rect 38222 14366 38274 14418
rect 2494 14254 2546 14306
rect 20414 14254 20466 14306
rect 22318 14254 22370 14306
rect 23774 14254 23826 14306
rect 37886 14254 37938 14306
rect 10538 14086 10590 14138
rect 10642 14086 10694 14138
rect 10746 14086 10798 14138
rect 19862 14086 19914 14138
rect 19966 14086 20018 14138
rect 20070 14086 20122 14138
rect 29186 14086 29238 14138
rect 29290 14086 29342 14138
rect 29394 14086 29446 14138
rect 38510 14086 38562 14138
rect 38614 14086 38666 14138
rect 38718 14086 38770 14138
rect 2046 13918 2098 13970
rect 17950 13918 18002 13970
rect 18062 13918 18114 13970
rect 37886 13918 37938 13970
rect 2718 13806 2770 13858
rect 20078 13806 20130 13858
rect 22430 13806 22482 13858
rect 22878 13806 22930 13858
rect 1710 13694 1762 13746
rect 2382 13694 2434 13746
rect 17838 13694 17890 13746
rect 19742 13694 19794 13746
rect 21870 13694 21922 13746
rect 22206 13694 22258 13746
rect 23550 13694 23602 13746
rect 24558 13694 24610 13746
rect 25454 13694 25506 13746
rect 38222 13694 38274 13746
rect 3166 13582 3218 13634
rect 3614 13582 3666 13634
rect 18286 13582 18338 13634
rect 18958 13582 19010 13634
rect 21422 13582 21474 13634
rect 37662 13582 37714 13634
rect 18510 13470 18562 13522
rect 19294 13470 19346 13522
rect 5876 13302 5928 13354
rect 5980 13302 6032 13354
rect 6084 13302 6136 13354
rect 15200 13302 15252 13354
rect 15304 13302 15356 13354
rect 15408 13302 15460 13354
rect 24524 13302 24576 13354
rect 24628 13302 24680 13354
rect 24732 13302 24784 13354
rect 33848 13302 33900 13354
rect 33952 13302 34004 13354
rect 34056 13302 34108 13354
rect 21310 13134 21362 13186
rect 1934 13022 1986 13074
rect 21870 13022 21922 13074
rect 4286 12910 4338 12962
rect 19294 12910 19346 12962
rect 19742 12910 19794 12962
rect 21534 12910 21586 12962
rect 21982 12910 22034 12962
rect 23214 12910 23266 12962
rect 23662 12910 23714 12962
rect 24222 12910 24274 12962
rect 25006 12910 25058 12962
rect 25902 12910 25954 12962
rect 20078 12798 20130 12850
rect 22766 12798 22818 12850
rect 37214 12798 37266 12850
rect 37550 12798 37602 12850
rect 37886 12798 37938 12850
rect 38222 12798 38274 12850
rect 18958 12686 19010 12738
rect 21758 12686 21810 12738
rect 23774 12686 23826 12738
rect 36542 12686 36594 12738
rect 10538 12518 10590 12570
rect 10642 12518 10694 12570
rect 10746 12518 10798 12570
rect 19862 12518 19914 12570
rect 19966 12518 20018 12570
rect 20070 12518 20122 12570
rect 29186 12518 29238 12570
rect 29290 12518 29342 12570
rect 29394 12518 29446 12570
rect 38510 12518 38562 12570
rect 38614 12518 38666 12570
rect 38718 12518 38770 12570
rect 18958 12350 19010 12402
rect 20974 12350 21026 12402
rect 21086 12350 21138 12402
rect 21198 12350 21250 12402
rect 19854 12238 19906 12290
rect 37886 12238 37938 12290
rect 4286 12126 4338 12178
rect 19742 12126 19794 12178
rect 20526 12126 20578 12178
rect 20750 12126 20802 12178
rect 37550 12126 37602 12178
rect 38222 12126 38274 12178
rect 37214 12014 37266 12066
rect 1934 11902 1986 11954
rect 19294 11902 19346 11954
rect 5876 11734 5928 11786
rect 5980 11734 6032 11786
rect 6084 11734 6136 11786
rect 15200 11734 15252 11786
rect 15304 11734 15356 11786
rect 15408 11734 15460 11786
rect 24524 11734 24576 11786
rect 24628 11734 24680 11786
rect 24732 11734 24784 11786
rect 33848 11734 33900 11786
rect 33952 11734 34004 11786
rect 34056 11734 34108 11786
rect 37886 11230 37938 11282
rect 38222 11230 38274 11282
rect 37662 11118 37714 11170
rect 10538 10950 10590 11002
rect 10642 10950 10694 11002
rect 10746 10950 10798 11002
rect 19862 10950 19914 11002
rect 19966 10950 20018 11002
rect 20070 10950 20122 11002
rect 29186 10950 29238 11002
rect 29290 10950 29342 11002
rect 29394 10950 29446 11002
rect 38510 10950 38562 11002
rect 38614 10950 38666 11002
rect 38718 10950 38770 11002
rect 37886 10670 37938 10722
rect 37662 10558 37714 10610
rect 38222 10558 38274 10610
rect 5876 10166 5928 10218
rect 5980 10166 6032 10218
rect 6084 10166 6136 10218
rect 15200 10166 15252 10218
rect 15304 10166 15356 10218
rect 15408 10166 15460 10218
rect 24524 10166 24576 10218
rect 24628 10166 24680 10218
rect 24732 10166 24784 10218
rect 33848 10166 33900 10218
rect 33952 10166 34004 10218
rect 34056 10166 34108 10218
rect 10538 9382 10590 9434
rect 10642 9382 10694 9434
rect 10746 9382 10798 9434
rect 19862 9382 19914 9434
rect 19966 9382 20018 9434
rect 20070 9382 20122 9434
rect 29186 9382 29238 9434
rect 29290 9382 29342 9434
rect 29394 9382 29446 9434
rect 38510 9382 38562 9434
rect 38614 9382 38666 9434
rect 38718 9382 38770 9434
rect 5876 8598 5928 8650
rect 5980 8598 6032 8650
rect 6084 8598 6136 8650
rect 15200 8598 15252 8650
rect 15304 8598 15356 8650
rect 15408 8598 15460 8650
rect 24524 8598 24576 8650
rect 24628 8598 24680 8650
rect 24732 8598 24784 8650
rect 33848 8598 33900 8650
rect 33952 8598 34004 8650
rect 34056 8598 34108 8650
rect 10538 7814 10590 7866
rect 10642 7814 10694 7866
rect 10746 7814 10798 7866
rect 19862 7814 19914 7866
rect 19966 7814 20018 7866
rect 20070 7814 20122 7866
rect 29186 7814 29238 7866
rect 29290 7814 29342 7866
rect 29394 7814 29446 7866
rect 38510 7814 38562 7866
rect 38614 7814 38666 7866
rect 38718 7814 38770 7866
rect 5876 7030 5928 7082
rect 5980 7030 6032 7082
rect 6084 7030 6136 7082
rect 15200 7030 15252 7082
rect 15304 7030 15356 7082
rect 15408 7030 15460 7082
rect 24524 7030 24576 7082
rect 24628 7030 24680 7082
rect 24732 7030 24784 7082
rect 33848 7030 33900 7082
rect 33952 7030 34004 7082
rect 34056 7030 34108 7082
rect 10538 6246 10590 6298
rect 10642 6246 10694 6298
rect 10746 6246 10798 6298
rect 19862 6246 19914 6298
rect 19966 6246 20018 6298
rect 20070 6246 20122 6298
rect 29186 6246 29238 6298
rect 29290 6246 29342 6298
rect 29394 6246 29446 6298
rect 38510 6246 38562 6298
rect 38614 6246 38666 6298
rect 38718 6246 38770 6298
rect 5876 5462 5928 5514
rect 5980 5462 6032 5514
rect 6084 5462 6136 5514
rect 15200 5462 15252 5514
rect 15304 5462 15356 5514
rect 15408 5462 15460 5514
rect 24524 5462 24576 5514
rect 24628 5462 24680 5514
rect 24732 5462 24784 5514
rect 33848 5462 33900 5514
rect 33952 5462 34004 5514
rect 34056 5462 34108 5514
rect 13694 5070 13746 5122
rect 14366 5070 14418 5122
rect 15038 5070 15090 5122
rect 14702 4958 14754 5010
rect 15374 4958 15426 5010
rect 14142 4846 14194 4898
rect 16606 4846 16658 4898
rect 22206 4846 22258 4898
rect 10538 4678 10590 4730
rect 10642 4678 10694 4730
rect 10746 4678 10798 4730
rect 19862 4678 19914 4730
rect 19966 4678 20018 4730
rect 20070 4678 20122 4730
rect 29186 4678 29238 4730
rect 29290 4678 29342 4730
rect 29394 4678 29446 4730
rect 38510 4678 38562 4730
rect 38614 4678 38666 4730
rect 38718 4678 38770 4730
rect 16046 4510 16098 4562
rect 21086 4510 21138 4562
rect 21758 4510 21810 4562
rect 22430 4510 22482 4562
rect 27134 4510 27186 4562
rect 29486 4510 29538 4562
rect 14926 4286 14978 4338
rect 15710 4286 15762 4338
rect 20862 4286 20914 4338
rect 21310 4286 21362 4338
rect 21982 4286 22034 4338
rect 22654 4286 22706 4338
rect 27358 4286 27410 4338
rect 15486 4174 15538 4226
rect 16830 4174 16882 4226
rect 17614 4174 17666 4226
rect 18174 4174 18226 4226
rect 18846 4174 18898 4226
rect 19966 4174 20018 4226
rect 20414 4174 20466 4226
rect 23438 4174 23490 4226
rect 24334 4174 24386 4226
rect 25454 4174 25506 4226
rect 25902 4174 25954 4226
rect 26350 4174 26402 4226
rect 26910 4174 26962 4226
rect 27918 4174 27970 4226
rect 28478 4174 28530 4226
rect 28926 4174 28978 4226
rect 30158 4174 30210 4226
rect 30830 4174 30882 4226
rect 12574 4062 12626 4114
rect 25566 4062 25618 4114
rect 26350 4062 26402 4114
rect 26798 4062 26850 4114
rect 5876 3894 5928 3946
rect 5980 3894 6032 3946
rect 6084 3894 6136 3946
rect 15200 3894 15252 3946
rect 15304 3894 15356 3946
rect 15408 3894 15460 3946
rect 24524 3894 24576 3946
rect 24628 3894 24680 3946
rect 24732 3894 24784 3946
rect 33848 3894 33900 3946
rect 33952 3894 34004 3946
rect 34056 3894 34108 3946
rect 13358 3614 13410 3666
rect 20974 3614 21026 3666
rect 12350 3502 12402 3554
rect 15710 3502 15762 3554
rect 16158 3502 16210 3554
rect 17054 3502 17106 3554
rect 17726 3502 17778 3554
rect 18622 3502 18674 3554
rect 19294 3502 19346 3554
rect 20078 3502 20130 3554
rect 22878 3502 22930 3554
rect 23886 3502 23938 3554
rect 24782 3502 24834 3554
rect 25454 3502 25506 3554
rect 26238 3502 26290 3554
rect 26798 3502 26850 3554
rect 27470 3502 27522 3554
rect 28590 3502 28642 3554
rect 29934 3502 29986 3554
rect 30606 3502 30658 3554
rect 31278 3502 31330 3554
rect 12014 3390 12066 3442
rect 12574 3390 12626 3442
rect 17390 3390 17442 3442
rect 18062 3390 18114 3442
rect 18398 3390 18450 3442
rect 19070 3390 19122 3442
rect 19854 3390 19906 3442
rect 23662 3390 23714 3442
rect 24558 3390 24610 3442
rect 25230 3390 25282 3442
rect 25902 3390 25954 3442
rect 26574 3390 26626 3442
rect 27246 3390 27298 3442
rect 28366 3390 28418 3442
rect 29374 3390 29426 3442
rect 29710 3390 29762 3442
rect 30382 3390 30434 3442
rect 31054 3390 31106 3442
rect 16382 3278 16434 3330
rect 29038 3278 29090 3330
rect 10538 3110 10590 3162
rect 10642 3110 10694 3162
rect 10746 3110 10798 3162
rect 19862 3110 19914 3162
rect 19966 3110 20018 3162
rect 20070 3110 20122 3162
rect 29186 3110 29238 3162
rect 29290 3110 29342 3162
rect 29394 3110 29446 3162
rect 38510 3110 38562 3162
rect 38614 3110 38666 3162
rect 38718 3110 38770 3162
rect 28926 2830 28978 2882
rect 29934 2830 29986 2882
<< metal2 >>
rect 10752 39200 10864 40000
rect 11424 39200 11536 40000
rect 12096 39200 12208 40000
rect 12768 39200 12880 40000
rect 13440 39200 13552 40000
rect 14112 39200 14224 40000
rect 14784 39200 14896 40000
rect 15456 39200 15568 40000
rect 16128 39200 16240 40000
rect 16800 39200 16912 40000
rect 17472 39200 17584 40000
rect 18144 39200 18256 40000
rect 18816 39200 18928 40000
rect 19488 39200 19600 40000
rect 20160 39200 20272 40000
rect 20832 39200 20944 40000
rect 21504 39200 21616 40000
rect 22176 39200 22288 40000
rect 22848 39200 22960 40000
rect 23520 39200 23632 40000
rect 24192 39200 24304 40000
rect 24864 39200 24976 40000
rect 25536 39200 25648 40000
rect 26208 39200 26320 40000
rect 26880 39200 26992 40000
rect 10780 36932 10836 39200
rect 11452 37156 11508 39200
rect 12124 37268 12180 39200
rect 5874 36876 6138 36886
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 10780 36866 10836 36876
rect 11004 37100 11508 37156
rect 11788 37212 12180 37268
rect 5874 36810 6138 36820
rect 10220 36596 10276 36606
rect 11004 36596 11060 37100
rect 10220 36594 11060 36596
rect 10220 36542 10222 36594
rect 10274 36542 11060 36594
rect 10220 36540 11060 36542
rect 10220 36530 10276 36540
rect 11004 36482 11060 36540
rect 11004 36430 11006 36482
rect 11058 36430 11060 36482
rect 11004 36418 11060 36430
rect 11452 36932 11508 36942
rect 10668 36372 10724 36382
rect 10668 36278 10724 36316
rect 11228 36260 11284 36270
rect 11116 36258 11284 36260
rect 11116 36206 11230 36258
rect 11282 36206 11284 36258
rect 11116 36204 11284 36206
rect 10536 36092 10800 36102
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10536 36026 10800 36036
rect 5874 35308 6138 35318
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 5874 35242 6138 35252
rect 10536 34524 10800 34534
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10536 34458 10800 34468
rect 5874 33740 6138 33750
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 5874 33674 6138 33684
rect 10536 32956 10800 32966
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10536 32890 10800 32900
rect 5874 32172 6138 32182
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 5874 32106 6138 32116
rect 11116 31948 11172 36204
rect 11228 36194 11284 36204
rect 11452 35586 11508 36876
rect 11676 36484 11732 36494
rect 11788 36484 11844 37212
rect 11676 36482 11844 36484
rect 11676 36430 11678 36482
rect 11730 36430 11844 36482
rect 11676 36428 11844 36430
rect 12348 36484 12404 36494
rect 12796 36484 12852 39200
rect 12348 36482 12852 36484
rect 12348 36430 12350 36482
rect 12402 36430 12852 36482
rect 12348 36428 12852 36430
rect 11676 36372 11732 36428
rect 12348 36418 12404 36428
rect 11676 36306 11732 36316
rect 11900 36260 11956 36270
rect 11900 36166 11956 36204
rect 12572 36258 12628 36270
rect 12572 36206 12574 36258
rect 12626 36206 12628 36258
rect 11452 35534 11454 35586
rect 11506 35534 11508 35586
rect 11452 35522 11508 35534
rect 11116 31892 11284 31948
rect 10536 31388 10800 31398
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10536 31322 10800 31332
rect 5874 30604 6138 30614
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 5874 30538 6138 30548
rect 10536 29820 10800 29830
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10536 29754 10800 29764
rect 4284 29428 4340 29438
rect 4284 29334 4340 29372
rect 1932 29204 1988 29214
rect 1932 29110 1988 29148
rect 5874 29036 6138 29046
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 5874 28970 6138 28980
rect 1708 28642 1764 28654
rect 1708 28590 1710 28642
rect 1762 28590 1764 28642
rect 1708 28308 1764 28590
rect 2492 28642 2548 28654
rect 2492 28590 2494 28642
rect 2546 28590 2548 28642
rect 2044 28420 2100 28430
rect 2044 28418 2436 28420
rect 2044 28366 2046 28418
rect 2098 28366 2436 28418
rect 2044 28364 2436 28366
rect 2044 28354 2100 28364
rect 1708 28242 1764 28252
rect 2380 28084 2436 28364
rect 2492 28308 2548 28590
rect 2492 28242 2548 28252
rect 10536 28252 10800 28262
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10536 28186 10800 28196
rect 2380 28028 2884 28084
rect 2044 27972 2100 27982
rect 2044 27970 2660 27972
rect 2044 27918 2046 27970
rect 2098 27918 2660 27970
rect 2044 27916 2660 27918
rect 2044 27906 2100 27916
rect 1708 27858 1764 27870
rect 1708 27806 1710 27858
rect 1762 27806 1764 27858
rect 1708 27636 1764 27806
rect 1708 27570 1764 27580
rect 2492 27746 2548 27758
rect 2492 27694 2494 27746
rect 2546 27694 2548 27746
rect 2492 27524 2548 27694
rect 1932 27468 2548 27524
rect 1820 27076 1876 27086
rect 1932 27076 1988 27468
rect 1820 27074 1988 27076
rect 1820 27022 1822 27074
rect 1874 27022 1988 27074
rect 1820 27020 1988 27022
rect 2044 27300 2100 27310
rect 1708 26290 1764 26302
rect 1708 26238 1710 26290
rect 1762 26238 1764 26290
rect 1708 26180 1764 26238
rect 1820 26292 1876 27020
rect 2044 26962 2100 27244
rect 2044 26910 2046 26962
rect 2098 26910 2100 26962
rect 2044 26898 2100 26910
rect 2380 26964 2436 26974
rect 2380 26870 2436 26908
rect 2044 26404 2100 26414
rect 2044 26310 2100 26348
rect 1820 26226 1876 26236
rect 1708 25620 1764 26124
rect 2492 26180 2548 26190
rect 2492 26086 2548 26124
rect 1708 25554 1764 25564
rect 1708 25394 1764 25406
rect 1708 25342 1710 25394
rect 1762 25342 1764 25394
rect 1708 24948 1764 25342
rect 2044 25284 2100 25294
rect 2044 25190 2100 25228
rect 2492 25282 2548 25294
rect 2492 25230 2494 25282
rect 2546 25230 2548 25282
rect 1708 24882 1764 24892
rect 2492 24948 2548 25230
rect 2492 24882 2548 24892
rect 2044 24836 2100 24846
rect 2044 24834 2324 24836
rect 2044 24782 2046 24834
rect 2098 24782 2324 24834
rect 2044 24780 2324 24782
rect 2044 24770 2100 24780
rect 1708 24722 1764 24734
rect 1708 24670 1710 24722
rect 1762 24670 1764 24722
rect 1708 24276 1764 24670
rect 1708 24210 1764 24220
rect 1708 23714 1764 23726
rect 1708 23662 1710 23714
rect 1762 23662 1764 23714
rect 1708 23604 1764 23662
rect 2044 23716 2100 23726
rect 2044 23622 2100 23660
rect 1708 23538 1764 23548
rect 2044 23268 2100 23278
rect 2044 23174 2100 23212
rect 1708 23154 1764 23166
rect 1708 23102 1710 23154
rect 1762 23102 1764 23154
rect 1708 22932 1764 23102
rect 1708 22866 1764 22876
rect 2044 22372 2100 22382
rect 1708 22260 1764 22270
rect 1708 22166 1764 22204
rect 2044 22258 2100 22316
rect 2044 22206 2046 22258
rect 2098 22206 2100 22258
rect 2044 22194 2100 22206
rect 2044 21700 2100 21710
rect 2044 21606 2100 21644
rect 1708 21586 1764 21598
rect 1708 21534 1710 21586
rect 1762 21534 1764 21586
rect 1708 21476 1764 21534
rect 1708 20916 1764 21420
rect 1708 20850 1764 20860
rect 1708 20578 1764 20590
rect 1708 20526 1710 20578
rect 1762 20526 1764 20578
rect 1708 20244 1764 20526
rect 2044 20580 2100 20590
rect 2268 20580 2324 24780
rect 2492 24610 2548 24622
rect 2492 24558 2494 24610
rect 2546 24558 2548 24610
rect 2492 24276 2548 24558
rect 2492 24210 2548 24220
rect 2492 23714 2548 23726
rect 2492 23662 2494 23714
rect 2546 23662 2548 23714
rect 2492 23604 2548 23662
rect 2492 23538 2548 23548
rect 2492 23042 2548 23054
rect 2492 22990 2494 23042
rect 2546 22990 2548 23042
rect 2492 22932 2548 22990
rect 2492 22866 2548 22876
rect 2492 22260 2548 22270
rect 2380 22146 2436 22158
rect 2380 22094 2382 22146
rect 2434 22094 2436 22146
rect 2380 21588 2436 22094
rect 2492 21810 2548 22204
rect 2492 21758 2494 21810
rect 2546 21758 2548 21810
rect 2492 21746 2548 21758
rect 2380 21522 2436 21532
rect 2604 21364 2660 27916
rect 2716 26850 2772 26862
rect 2716 26798 2718 26850
rect 2770 26798 2772 26850
rect 2716 24052 2772 26798
rect 2716 23986 2772 23996
rect 2604 21298 2660 21308
rect 2716 22146 2772 22158
rect 2716 22094 2718 22146
rect 2770 22094 2772 22146
rect 2044 20578 2212 20580
rect 2044 20526 2046 20578
rect 2098 20526 2212 20578
rect 2044 20524 2212 20526
rect 2044 20514 2100 20524
rect 1708 20178 1764 20188
rect 2044 20132 2100 20142
rect 2044 20038 2100 20076
rect 1708 20018 1764 20030
rect 1708 19966 1710 20018
rect 1762 19966 1764 20018
rect 1708 19572 1764 19966
rect 2156 19796 2212 20524
rect 2268 20514 2324 20524
rect 2492 20578 2548 20590
rect 2492 20526 2494 20578
rect 2546 20526 2548 20578
rect 2492 20244 2548 20526
rect 2492 20178 2548 20188
rect 2156 19730 2212 19740
rect 2492 19906 2548 19918
rect 2492 19854 2494 19906
rect 2546 19854 2548 19906
rect 1708 19506 1764 19516
rect 2492 19572 2548 19854
rect 2492 19506 2548 19516
rect 1932 19346 1988 19358
rect 1932 19294 1934 19346
rect 1986 19294 1988 19346
rect 1932 18900 1988 19294
rect 2716 19348 2772 22094
rect 2828 20916 2884 28028
rect 2940 27746 2996 27758
rect 2940 27694 2942 27746
rect 2994 27694 2996 27746
rect 2940 27636 2996 27694
rect 2940 27570 2996 27580
rect 5874 27468 6138 27478
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 5874 27402 6138 27412
rect 3164 26964 3220 26974
rect 3164 26870 3220 26908
rect 10536 26684 10800 26694
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10536 26618 10800 26628
rect 11228 26516 11284 31892
rect 12572 27188 12628 36206
rect 12796 35026 12852 36428
rect 13468 36484 13524 39200
rect 14140 36484 14196 39200
rect 14812 36484 14868 39200
rect 15484 37044 15540 39200
rect 15484 36988 15652 37044
rect 15198 36876 15462 36886
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15198 36810 15462 36820
rect 15484 36484 15540 36494
rect 15596 36484 15652 36988
rect 16156 36708 16212 39200
rect 16156 36642 16212 36652
rect 16156 36484 16212 36494
rect 13468 36482 14084 36484
rect 13468 36430 13470 36482
rect 13522 36430 14084 36482
rect 13468 36428 14084 36430
rect 13468 36418 13524 36428
rect 13692 36258 13748 36270
rect 13692 36206 13694 36258
rect 13746 36206 13748 36258
rect 12796 34974 12798 35026
rect 12850 34974 12852 35026
rect 12796 34962 12852 34974
rect 13356 35698 13412 35710
rect 13356 35646 13358 35698
rect 13410 35646 13412 35698
rect 12572 27122 12628 27132
rect 11228 26450 11284 26460
rect 12572 26964 12628 26974
rect 5874 25900 6138 25910
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 5874 25834 6138 25844
rect 12348 25284 12404 25294
rect 10536 25116 10800 25126
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10536 25050 10800 25060
rect 12348 24722 12404 25228
rect 12348 24670 12350 24722
rect 12402 24670 12404 24722
rect 12348 24658 12404 24670
rect 12572 24722 12628 26908
rect 12572 24670 12574 24722
rect 12626 24670 12628 24722
rect 12460 24500 12516 24510
rect 5874 24332 6138 24342
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 5874 24266 6138 24276
rect 12460 24050 12516 24444
rect 12460 23998 12462 24050
rect 12514 23998 12516 24050
rect 12460 23986 12516 23998
rect 12348 23604 12404 23614
rect 10536 23548 10800 23558
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10536 23482 10800 23492
rect 5874 22764 6138 22774
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 5874 22698 6138 22708
rect 3164 22146 3220 22158
rect 3164 22094 3166 22146
rect 3218 22094 3220 22146
rect 3164 21588 3220 22094
rect 10536 21980 10800 21990
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10536 21914 10800 21924
rect 3164 21522 3220 21532
rect 12236 21700 12292 21710
rect 2940 21476 2996 21486
rect 2940 21382 2996 21420
rect 12124 21474 12180 21486
rect 12124 21422 12126 21474
rect 12178 21422 12180 21474
rect 12124 21364 12180 21422
rect 12124 21298 12180 21308
rect 5874 21196 6138 21206
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 5874 21130 6138 21140
rect 12236 21140 12292 21644
rect 12348 21586 12404 23548
rect 12348 21534 12350 21586
rect 12402 21534 12404 21586
rect 12348 21522 12404 21534
rect 12236 21084 12404 21140
rect 2828 20850 2884 20860
rect 11340 20804 11396 20814
rect 11340 20710 11396 20748
rect 11788 20692 11844 20702
rect 11788 20598 11844 20636
rect 10536 20412 10800 20422
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10536 20346 10800 20356
rect 12236 20132 12292 20142
rect 5874 19628 6138 19638
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 5874 19562 6138 19572
rect 2716 19282 2772 19292
rect 12236 19346 12292 20076
rect 12348 20018 12404 21084
rect 12460 20916 12516 20926
rect 12460 20822 12516 20860
rect 12348 19966 12350 20018
rect 12402 19966 12404 20018
rect 12348 19954 12404 19966
rect 12236 19294 12238 19346
rect 12290 19294 12292 19346
rect 12236 19282 12292 19294
rect 4284 19236 4340 19246
rect 4284 19142 4340 19180
rect 12572 19234 12628 24670
rect 12908 25396 12964 25406
rect 12908 23714 12964 25340
rect 13132 24724 13188 24734
rect 13132 24630 13188 24668
rect 13356 24164 13412 35646
rect 13692 31948 13748 36206
rect 14028 35922 14084 36428
rect 14140 36482 14644 36484
rect 14140 36430 14142 36482
rect 14194 36430 14644 36482
rect 14140 36428 14644 36430
rect 14140 36418 14196 36428
rect 14028 35870 14030 35922
rect 14082 35870 14084 35922
rect 14028 35858 14084 35870
rect 14364 36258 14420 36270
rect 14364 36206 14366 36258
rect 14418 36206 14420 36258
rect 13692 31892 13860 31948
rect 13580 27300 13636 27310
rect 13580 25394 13636 27244
rect 13580 25342 13582 25394
rect 13634 25342 13636 25394
rect 13580 25330 13636 25342
rect 13692 25506 13748 25518
rect 13692 25454 13694 25506
rect 13746 25454 13748 25506
rect 13692 25396 13748 25454
rect 13692 25330 13748 25340
rect 13804 24948 13860 31892
rect 14364 29204 14420 36206
rect 14588 35922 14644 36428
rect 14812 36482 15316 36484
rect 14812 36430 14814 36482
rect 14866 36430 15316 36482
rect 14812 36428 15316 36430
rect 14812 36418 14868 36428
rect 14588 35870 14590 35922
rect 14642 35870 14644 35922
rect 14588 35858 14644 35870
rect 15036 36258 15092 36270
rect 15036 36206 15038 36258
rect 15090 36206 15092 36258
rect 14364 29138 14420 29148
rect 15036 28868 15092 36206
rect 15260 35922 15316 36428
rect 15484 36482 15988 36484
rect 15484 36430 15486 36482
rect 15538 36430 15988 36482
rect 15484 36428 15988 36430
rect 15484 36418 15540 36428
rect 15260 35870 15262 35922
rect 15314 35870 15316 35922
rect 15260 35858 15316 35870
rect 15708 36258 15764 36270
rect 15708 36206 15710 36258
rect 15762 36206 15764 36258
rect 15198 35308 15462 35318
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15198 35242 15462 35252
rect 15198 33740 15462 33750
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15198 33674 15462 33684
rect 15198 32172 15462 32182
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15198 32106 15462 32116
rect 15198 30604 15462 30614
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15198 30538 15462 30548
rect 15708 29428 15764 36206
rect 15932 35922 15988 36428
rect 16156 36390 16212 36428
rect 16492 36484 16548 36494
rect 15932 35870 15934 35922
rect 15986 35870 15988 35922
rect 15932 35858 15988 35870
rect 16380 36258 16436 36270
rect 16380 36206 16382 36258
rect 16434 36206 16436 36258
rect 15708 29372 16324 29428
rect 15820 29204 15876 29214
rect 15198 29036 15462 29046
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15198 28970 15462 28980
rect 15036 28802 15092 28812
rect 15708 28868 15764 28878
rect 15036 27860 15092 27870
rect 15036 26514 15092 27804
rect 15198 27468 15462 27478
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15198 27402 15462 27412
rect 15036 26462 15038 26514
rect 15090 26462 15092 26514
rect 15036 26450 15092 26462
rect 14364 26404 14420 26414
rect 14364 25730 14420 26348
rect 14812 26402 14868 26414
rect 14812 26350 14814 26402
rect 14866 26350 14868 26402
rect 14364 25678 14366 25730
rect 14418 25678 14420 25730
rect 14364 25666 14420 25678
rect 14700 26290 14756 26302
rect 14700 26238 14702 26290
rect 14754 26238 14756 26290
rect 14700 25730 14756 26238
rect 14812 26292 14868 26350
rect 14812 26226 14868 26236
rect 15596 26290 15652 26302
rect 15596 26238 15598 26290
rect 15650 26238 15652 26290
rect 15198 25900 15462 25910
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15198 25834 15462 25844
rect 14700 25678 14702 25730
rect 14754 25678 14756 25730
rect 14700 25666 14756 25678
rect 13804 24882 13860 24892
rect 15596 25506 15652 26238
rect 15708 25618 15764 28812
rect 15820 26178 15876 29148
rect 15820 26126 15822 26178
rect 15874 26126 15876 26178
rect 15820 26114 15876 26126
rect 15932 29092 15988 29102
rect 15708 25566 15710 25618
rect 15762 25566 15764 25618
rect 15708 25554 15764 25566
rect 15596 25454 15598 25506
rect 15650 25454 15652 25506
rect 14700 24724 14756 24734
rect 14700 24630 14756 24668
rect 13356 24098 13412 24108
rect 14588 24610 14644 24622
rect 14588 24558 14590 24610
rect 14642 24558 14644 24610
rect 14588 24162 14644 24558
rect 14588 24110 14590 24162
rect 14642 24110 14644 24162
rect 14588 24098 14644 24110
rect 14700 24500 14756 24510
rect 14364 24052 14420 24062
rect 14364 23938 14420 23996
rect 14364 23886 14366 23938
rect 14418 23886 14420 23938
rect 14364 23874 14420 23886
rect 14700 23938 14756 24444
rect 15596 24500 15652 25454
rect 15198 24332 15462 24342
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15198 24266 15462 24276
rect 15596 24164 15652 24444
rect 14700 23886 14702 23938
rect 14754 23886 14756 23938
rect 14700 23874 14756 23886
rect 15484 24108 15652 24164
rect 15708 24722 15764 24734
rect 15708 24670 15710 24722
rect 15762 24670 15764 24722
rect 12908 23662 12910 23714
rect 12962 23662 12964 23714
rect 12908 23156 12964 23662
rect 13916 23714 13972 23726
rect 13916 23662 13918 23714
rect 13970 23662 13972 23714
rect 13916 23380 13972 23662
rect 13692 23324 13972 23380
rect 13132 23156 13188 23166
rect 12908 23100 13132 23156
rect 13132 23042 13188 23100
rect 13132 22990 13134 23042
rect 13186 22990 13188 23042
rect 13132 22978 13188 22990
rect 13580 23156 13636 23166
rect 13692 23156 13748 23324
rect 13580 23154 13748 23156
rect 13580 23102 13582 23154
rect 13634 23102 13748 23154
rect 13580 23100 13748 23102
rect 13804 23156 13860 23166
rect 13580 22148 13636 23100
rect 13804 22370 13860 23100
rect 15036 23154 15092 23166
rect 15036 23102 15038 23154
rect 15090 23102 15092 23154
rect 14476 23044 14532 23054
rect 14476 23042 14644 23044
rect 14476 22990 14478 23042
rect 14530 22990 14644 23042
rect 14476 22988 14644 22990
rect 14476 22978 14532 22988
rect 13804 22318 13806 22370
rect 13858 22318 13860 22370
rect 13804 22306 13860 22318
rect 13580 22082 13636 22092
rect 14476 22146 14532 22158
rect 14476 22094 14478 22146
rect 14530 22094 14532 22146
rect 14476 21700 14532 22094
rect 14476 21634 14532 21644
rect 13580 21586 13636 21598
rect 13580 21534 13582 21586
rect 13634 21534 13636 21586
rect 12908 21028 12964 21038
rect 12908 20802 12964 20972
rect 13580 20916 13636 21534
rect 14588 21588 14644 22988
rect 15036 22484 15092 23102
rect 15484 22932 15540 24108
rect 15596 23938 15652 23950
rect 15596 23886 15598 23938
rect 15650 23886 15652 23938
rect 15596 23492 15652 23886
rect 15596 23426 15652 23436
rect 15596 23156 15652 23166
rect 15596 23062 15652 23100
rect 15484 22876 15652 22932
rect 15198 22764 15462 22774
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15198 22698 15462 22708
rect 15036 22418 15092 22428
rect 15596 22482 15652 22876
rect 15596 22430 15598 22482
rect 15650 22430 15652 22482
rect 15596 22418 15652 22430
rect 14924 21588 14980 21598
rect 14588 21586 14980 21588
rect 14588 21534 14926 21586
rect 14978 21534 14980 21586
rect 14588 21532 14980 21534
rect 12908 20750 12910 20802
rect 12962 20750 12964 20802
rect 12908 20738 12964 20750
rect 13468 20804 13524 20814
rect 13580 20804 13636 20860
rect 13804 20804 13860 20814
rect 13580 20802 13860 20804
rect 13580 20750 13806 20802
rect 13858 20750 13860 20802
rect 13580 20748 13860 20750
rect 13468 20710 13524 20748
rect 13580 20020 13636 20030
rect 13804 20020 13860 20748
rect 13580 20018 13860 20020
rect 13580 19966 13582 20018
rect 13634 19966 13860 20018
rect 13580 19964 13860 19966
rect 13580 19954 13636 19964
rect 12908 19460 12964 19470
rect 12908 19346 12964 19404
rect 12908 19294 12910 19346
rect 12962 19294 12964 19346
rect 12908 19282 12964 19294
rect 12572 19182 12574 19234
rect 12626 19182 12628 19234
rect 1932 18834 1988 18844
rect 10536 18844 10800 18854
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10536 18778 10800 18788
rect 2044 18562 2100 18574
rect 2044 18510 2046 18562
rect 2098 18510 2100 18562
rect 1708 18450 1764 18462
rect 1708 18398 1710 18450
rect 1762 18398 1764 18450
rect 1708 18228 1764 18398
rect 2044 18452 2100 18510
rect 2044 18386 2100 18396
rect 1708 18162 1764 18172
rect 2492 18338 2548 18350
rect 2492 18286 2494 18338
rect 2546 18286 2548 18338
rect 2492 18228 2548 18286
rect 2492 18162 2548 18172
rect 12572 18228 12628 19182
rect 13468 19236 13524 19246
rect 13468 19142 13524 19180
rect 13804 19234 13860 19964
rect 13804 19182 13806 19234
rect 13858 19182 13860 19234
rect 13804 19170 13860 19182
rect 14924 20188 14980 21532
rect 15372 21586 15428 21598
rect 15372 21534 15374 21586
rect 15426 21534 15428 21586
rect 15372 21364 15428 21534
rect 15372 21298 15428 21308
rect 15708 21362 15764 24670
rect 15820 24500 15876 24510
rect 15932 24500 15988 29036
rect 16268 27074 16324 29372
rect 16268 27022 16270 27074
rect 16322 27022 16324 27074
rect 16268 27010 16324 27022
rect 16380 26908 16436 36206
rect 16492 35922 16548 36428
rect 16828 36484 16884 39200
rect 17164 36708 17220 36718
rect 17164 36614 17220 36652
rect 16828 36418 16884 36428
rect 16492 35870 16494 35922
rect 16546 35870 16548 35922
rect 16492 35858 16548 35870
rect 16940 35924 16996 35934
rect 17500 35924 17556 39200
rect 16940 35922 17556 35924
rect 16940 35870 16942 35922
rect 16994 35870 17556 35922
rect 16940 35868 17556 35870
rect 16940 35858 16996 35868
rect 17500 35812 17556 35868
rect 17724 35812 17780 35822
rect 17500 35810 17780 35812
rect 17500 35758 17726 35810
rect 17778 35758 17780 35810
rect 17500 35756 17780 35758
rect 17724 35746 17780 35756
rect 18060 35812 18116 35822
rect 18060 35718 18116 35756
rect 18172 35812 18228 39200
rect 18396 35812 18452 35822
rect 18172 35810 18452 35812
rect 18172 35758 18398 35810
rect 18450 35758 18452 35810
rect 18172 35756 18452 35758
rect 18172 35026 18228 35756
rect 18396 35746 18452 35756
rect 18732 35810 18788 35822
rect 18732 35758 18734 35810
rect 18786 35758 18788 35810
rect 18172 34974 18174 35026
rect 18226 34974 18228 35026
rect 18172 34962 18228 34974
rect 17500 27188 17556 27198
rect 16492 27076 16548 27114
rect 17500 27094 17556 27132
rect 16492 27010 16548 27020
rect 17612 27076 17668 27086
rect 17612 26982 17668 27020
rect 18732 27074 18788 35758
rect 18844 35812 18900 39200
rect 19516 37044 19572 39200
rect 19516 36988 19908 37044
rect 19180 36482 19236 36494
rect 19852 36484 19908 36988
rect 20188 36932 20244 39200
rect 20188 36866 20244 36876
rect 20860 36708 20916 39200
rect 20860 36642 20916 36652
rect 21420 36932 21476 36942
rect 21084 36484 21140 36494
rect 19180 36430 19182 36482
rect 19234 36430 19236 36482
rect 19068 35812 19124 35822
rect 18844 35810 19124 35812
rect 18844 35758 19070 35810
rect 19122 35758 19124 35810
rect 18844 35756 19124 35758
rect 18844 35026 18900 35756
rect 19068 35746 19124 35756
rect 18844 34974 18846 35026
rect 18898 34974 18900 35026
rect 18844 34962 18900 34974
rect 18732 27022 18734 27074
rect 18786 27022 18788 27074
rect 18732 27010 18788 27022
rect 17052 26962 17108 26974
rect 17052 26910 17054 26962
rect 17106 26910 17108 26962
rect 16380 26852 16772 26908
rect 16604 26292 16660 26302
rect 16380 26178 16436 26190
rect 16380 26126 16382 26178
rect 16434 26126 16436 26178
rect 16268 24836 16324 24846
rect 16268 24742 16324 24780
rect 15820 24498 15988 24500
rect 15820 24446 15822 24498
rect 15874 24446 15988 24498
rect 15820 24444 15988 24446
rect 15820 24434 15876 24444
rect 16380 23940 16436 26126
rect 16492 25618 16548 25630
rect 16492 25566 16494 25618
rect 16546 25566 16548 25618
rect 16492 25508 16548 25566
rect 16492 25442 16548 25452
rect 16604 25506 16660 26236
rect 16604 25454 16606 25506
rect 16658 25454 16660 25506
rect 16380 23874 16436 23884
rect 16268 23714 16324 23726
rect 16268 23662 16270 23714
rect 16322 23662 16324 23714
rect 15932 22372 15988 22382
rect 15932 22278 15988 22316
rect 15708 21310 15710 21362
rect 15762 21310 15764 21362
rect 15708 21298 15764 21310
rect 15820 21700 15876 21710
rect 15820 21474 15876 21644
rect 15820 21422 15822 21474
rect 15874 21422 15876 21474
rect 15198 21196 15462 21206
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15198 21130 15462 21140
rect 15820 20916 15876 21422
rect 16268 21028 16324 23662
rect 16492 23492 16548 23502
rect 16604 23492 16660 25454
rect 16716 24612 16772 26852
rect 17052 25284 17108 26910
rect 18172 26962 18228 26974
rect 18172 26910 18174 26962
rect 18226 26910 18228 26962
rect 17724 26516 17780 26526
rect 17724 26422 17780 26460
rect 17388 25508 17444 25518
rect 18172 25508 18228 26910
rect 18508 26962 18564 26974
rect 18508 26910 18510 26962
rect 18562 26910 18564 26962
rect 18508 26292 18564 26910
rect 18508 26290 18788 26292
rect 18508 26238 18510 26290
rect 18562 26238 18788 26290
rect 18508 26236 18788 26238
rect 18508 26226 18564 26236
rect 18620 25508 18676 25518
rect 18172 25506 18676 25508
rect 18172 25454 18622 25506
rect 18674 25454 18676 25506
rect 18172 25452 18676 25454
rect 17388 25414 17444 25452
rect 18620 25442 18676 25452
rect 17052 25218 17108 25228
rect 18620 25284 18676 25294
rect 17948 24948 18004 24958
rect 17948 24722 18004 24892
rect 17948 24670 17950 24722
rect 18002 24670 18004 24722
rect 17948 24658 18004 24670
rect 16716 24546 16772 24556
rect 17836 24164 17892 24174
rect 17836 24070 17892 24108
rect 16716 24052 16772 24062
rect 16716 23958 16772 23996
rect 17500 23940 17556 23950
rect 17500 23846 17556 23884
rect 18620 23938 18676 25228
rect 18620 23886 18622 23938
rect 18674 23886 18676 23938
rect 18620 23874 18676 23886
rect 18732 24722 18788 26236
rect 19180 25618 19236 36430
rect 19740 36482 19908 36484
rect 19740 36430 19854 36482
rect 19906 36430 19908 36482
rect 19740 36428 19908 36430
rect 19628 36260 19684 36270
rect 19180 25566 19182 25618
rect 19234 25566 19236 25618
rect 19180 25554 19236 25566
rect 19292 35812 19348 35822
rect 18732 24670 18734 24722
rect 18786 24670 18788 24722
rect 18732 24052 18788 24670
rect 18732 23716 18788 23996
rect 18620 23660 18788 23716
rect 16548 23436 16660 23492
rect 17388 23492 17444 23502
rect 16492 23426 16548 23436
rect 16716 23268 16772 23278
rect 16716 23174 16772 23212
rect 17388 23154 17444 23436
rect 18620 23266 18676 23660
rect 18620 23214 18622 23266
rect 18674 23214 18676 23266
rect 18620 23202 18676 23214
rect 17388 23102 17390 23154
rect 17442 23102 17444 23154
rect 17388 23090 17444 23102
rect 17836 23154 17892 23166
rect 17836 23102 17838 23154
rect 17890 23102 17892 23154
rect 17612 22932 17668 22942
rect 16828 22484 16884 22494
rect 16828 22370 16884 22428
rect 16828 22318 16830 22370
rect 16882 22318 16884 22370
rect 16828 22306 16884 22318
rect 17388 22484 17444 22494
rect 17388 21810 17444 22428
rect 17612 22370 17668 22876
rect 17612 22318 17614 22370
rect 17666 22318 17668 22370
rect 17612 22306 17668 22318
rect 17724 22482 17780 22494
rect 17724 22430 17726 22482
rect 17778 22430 17780 22482
rect 17388 21758 17390 21810
rect 17442 21758 17444 21810
rect 17388 21746 17444 21758
rect 16268 20962 16324 20972
rect 17388 21026 17444 21038
rect 17388 20974 17390 21026
rect 17442 20974 17444 21026
rect 15372 20802 15428 20814
rect 15372 20750 15374 20802
rect 15426 20750 15428 20802
rect 15372 20188 15428 20750
rect 14924 20132 15428 20188
rect 14924 20018 14980 20132
rect 14924 19966 14926 20018
rect 14978 19966 14980 20018
rect 14924 19236 14980 19966
rect 15372 20020 15428 20030
rect 15372 19926 15428 19964
rect 15820 19906 15876 20860
rect 16940 20916 16996 20926
rect 16996 20860 17108 20916
rect 16940 20822 16996 20860
rect 16828 20802 16884 20814
rect 16828 20750 16830 20802
rect 16882 20750 16884 20802
rect 16828 20692 16884 20750
rect 16828 20626 16884 20636
rect 15820 19854 15822 19906
rect 15874 19854 15876 19906
rect 15820 19842 15876 19854
rect 15708 19794 15764 19806
rect 15708 19742 15710 19794
rect 15762 19742 15764 19794
rect 15198 19628 15462 19638
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15198 19562 15462 19572
rect 15596 19346 15652 19358
rect 15596 19294 15598 19346
rect 15650 19294 15652 19346
rect 15372 19236 15428 19246
rect 14924 19234 15428 19236
rect 14924 19182 15374 19234
rect 15426 19182 15428 19234
rect 14924 19180 15428 19182
rect 15372 19170 15428 19180
rect 14924 18676 14980 18686
rect 14812 18620 14924 18676
rect 13468 18450 13524 18462
rect 14700 18452 14756 18462
rect 13468 18398 13470 18450
rect 13522 18398 13524 18450
rect 12572 18162 12628 18172
rect 13020 18340 13076 18350
rect 5874 18060 6138 18070
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 5874 17994 6138 18004
rect 12796 17892 12852 17902
rect 12796 17798 12852 17836
rect 1932 17780 1988 17790
rect 2156 17780 2212 17790
rect 1932 17686 1988 17724
rect 2044 17724 2156 17780
rect 2044 17220 2100 17724
rect 2156 17714 2212 17724
rect 11788 17778 11844 17790
rect 11788 17726 11790 17778
rect 11842 17726 11844 17778
rect 1932 17164 2100 17220
rect 2716 17668 2772 17678
rect 1708 16884 1764 16894
rect 1708 16790 1764 16828
rect 1708 15986 1764 15998
rect 1708 15934 1710 15986
rect 1762 15934 1764 15986
rect 1708 15540 1764 15934
rect 1708 15474 1764 15484
rect 1708 15314 1764 15326
rect 1708 15262 1710 15314
rect 1762 15262 1764 15314
rect 1708 14868 1764 15262
rect 1708 14802 1764 14812
rect 1708 14418 1764 14430
rect 1708 14366 1710 14418
rect 1762 14366 1764 14418
rect 1708 14196 1764 14366
rect 1932 14420 1988 17164
rect 2716 17106 2772 17612
rect 2716 17054 2718 17106
rect 2770 17054 2772 17106
rect 2716 17042 2772 17054
rect 4284 17666 4340 17678
rect 4284 17614 4286 17666
rect 4338 17614 4340 17666
rect 2044 16994 2100 17006
rect 2044 16942 2046 16994
rect 2098 16942 2100 16994
rect 2044 16324 2100 16942
rect 2380 16882 2436 16894
rect 2380 16830 2382 16882
rect 2434 16830 2436 16882
rect 2380 16772 2436 16830
rect 2268 16660 2324 16670
rect 2044 16258 2100 16268
rect 2156 16604 2268 16660
rect 2044 15876 2100 15886
rect 2044 15782 2100 15820
rect 2044 15428 2100 15438
rect 2044 15334 2100 15372
rect 2044 14420 2100 14430
rect 1932 14418 2100 14420
rect 1932 14366 2046 14418
rect 2098 14366 2100 14418
rect 1932 14364 2100 14366
rect 2044 14354 2100 14364
rect 1708 14130 1764 14140
rect 2044 13972 2100 13982
rect 2156 13972 2212 16604
rect 2268 16594 2324 16604
rect 2380 16212 2436 16716
rect 2380 16146 2436 16156
rect 2492 16884 2548 16894
rect 2492 16210 2548 16828
rect 3164 16882 3220 16894
rect 3164 16830 3166 16882
rect 3218 16830 3220 16882
rect 3164 16772 3220 16830
rect 3164 16706 3220 16716
rect 4284 16660 4340 17614
rect 11788 17668 11844 17726
rect 11788 17602 11844 17612
rect 12236 17668 12292 17678
rect 12236 17574 12292 17612
rect 13020 17666 13076 18284
rect 13468 17892 13524 18398
rect 13468 17826 13524 17836
rect 14476 18450 14756 18452
rect 14476 18398 14702 18450
rect 14754 18398 14756 18450
rect 14476 18396 14756 18398
rect 13020 17614 13022 17666
rect 13074 17614 13076 17666
rect 13020 17602 13076 17614
rect 13804 17780 13860 17790
rect 13804 17666 13860 17724
rect 13804 17614 13806 17666
rect 13858 17614 13860 17666
rect 13804 17602 13860 17614
rect 14028 17668 14084 17678
rect 14084 17612 14308 17668
rect 14028 17574 14084 17612
rect 10536 17276 10800 17286
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10536 17210 10800 17220
rect 12796 16882 12852 16894
rect 12796 16830 12798 16882
rect 12850 16830 12852 16882
rect 12460 16772 12516 16782
rect 12460 16678 12516 16716
rect 4284 16594 4340 16604
rect 5874 16492 6138 16502
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 5874 16426 6138 16436
rect 12796 16436 12852 16830
rect 13132 16884 13188 16894
rect 13132 16790 13188 16828
rect 13916 16660 13972 16670
rect 13916 16566 13972 16604
rect 12796 16370 12852 16380
rect 14140 16436 14196 16446
rect 2492 16158 2494 16210
rect 2546 16158 2548 16210
rect 2492 16146 2548 16158
rect 13804 16212 13860 16222
rect 13804 16118 13860 16156
rect 14140 16098 14196 16380
rect 14140 16046 14142 16098
rect 14194 16046 14196 16098
rect 2940 15874 2996 15886
rect 2940 15822 2942 15874
rect 2994 15822 2996 15874
rect 2940 15540 2996 15822
rect 10536 15708 10800 15718
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10536 15642 10800 15652
rect 2940 15474 2996 15484
rect 14140 15428 14196 16046
rect 14140 15362 14196 15372
rect 14252 16100 14308 17612
rect 14476 16210 14532 18396
rect 14700 18386 14756 18396
rect 14812 17778 14868 18620
rect 14924 18610 14980 18620
rect 15596 18450 15652 19294
rect 15596 18398 15598 18450
rect 15650 18398 15652 18450
rect 15596 18386 15652 18398
rect 14812 17726 14814 17778
rect 14866 17726 14868 17778
rect 14812 17714 14868 17726
rect 14924 18340 14980 18350
rect 14924 17666 14980 18284
rect 15198 18060 15462 18070
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15198 17994 15462 18004
rect 14924 17614 14926 17666
rect 14978 17614 14980 17666
rect 14924 17602 14980 17614
rect 15484 17668 15540 17678
rect 15484 17666 15652 17668
rect 15484 17614 15486 17666
rect 15538 17614 15652 17666
rect 15484 17612 15652 17614
rect 15484 17602 15540 17612
rect 14700 16884 14756 16894
rect 14700 16790 14756 16828
rect 14476 16158 14478 16210
rect 14530 16158 14532 16210
rect 14476 16146 14532 16158
rect 14588 16770 14644 16782
rect 14588 16718 14590 16770
rect 14642 16718 14644 16770
rect 14028 15316 14084 15326
rect 14028 15222 14084 15260
rect 14252 15314 14308 16044
rect 14588 15426 14644 16718
rect 15198 16492 15462 16502
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15198 16426 15462 16436
rect 15596 16322 15652 17612
rect 15708 16882 15764 19742
rect 17052 19346 17108 20860
rect 17388 20188 17444 20974
rect 17388 20132 17668 20188
rect 17612 20018 17668 20132
rect 17612 19966 17614 20018
rect 17666 19966 17668 20018
rect 17612 19954 17668 19966
rect 17052 19294 17054 19346
rect 17106 19294 17108 19346
rect 17052 19282 17108 19294
rect 16828 19234 16884 19246
rect 16828 19182 16830 19234
rect 16882 19182 16884 19234
rect 16268 18562 16324 18574
rect 16268 18510 16270 18562
rect 16322 18510 16324 18562
rect 15708 16830 15710 16882
rect 15762 16830 15764 16882
rect 15708 16818 15764 16830
rect 15820 18340 15876 18350
rect 15596 16270 15598 16322
rect 15650 16270 15652 16322
rect 15596 16258 15652 16270
rect 15372 16210 15428 16222
rect 15372 16158 15374 16210
rect 15426 16158 15428 16210
rect 15148 16100 15204 16110
rect 15148 16006 15204 16044
rect 15372 15876 15428 16158
rect 15820 16100 15876 18284
rect 15372 15810 15428 15820
rect 15484 16098 15876 16100
rect 15484 16046 15822 16098
rect 15874 16046 15876 16098
rect 15484 16044 15876 16046
rect 14588 15374 14590 15426
rect 14642 15374 14644 15426
rect 14588 15362 14644 15374
rect 14252 15262 14254 15314
rect 14306 15262 14308 15314
rect 14252 15250 14308 15262
rect 15372 15316 15428 15326
rect 15484 15316 15540 16044
rect 15820 16034 15876 16044
rect 15932 18226 15988 18238
rect 15932 18174 15934 18226
rect 15986 18174 15988 18226
rect 15372 15314 15540 15316
rect 15372 15262 15374 15314
rect 15426 15262 15540 15314
rect 15372 15260 15540 15262
rect 15372 15250 15428 15260
rect 2492 15202 2548 15214
rect 2492 15150 2494 15202
rect 2546 15150 2548 15202
rect 2492 14868 2548 15150
rect 15708 15202 15764 15214
rect 15708 15150 15710 15202
rect 15762 15150 15764 15202
rect 5874 14924 6138 14934
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 5874 14858 6138 14868
rect 15198 14924 15462 14934
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15198 14858 15462 14868
rect 2492 14802 2548 14812
rect 2492 14306 2548 14318
rect 2492 14254 2494 14306
rect 2546 14254 2548 14306
rect 2492 14196 2548 14254
rect 2492 14130 2548 14140
rect 10536 14140 10800 14150
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10536 14074 10800 14084
rect 2044 13970 2212 13972
rect 2044 13918 2046 13970
rect 2098 13918 2212 13970
rect 2044 13916 2212 13918
rect 2044 13906 2100 13916
rect 2716 13860 2772 13870
rect 2716 13766 2772 13804
rect 15708 13860 15764 15150
rect 15708 13794 15764 13804
rect 15820 14308 15876 14318
rect 1708 13746 1764 13758
rect 1708 13694 1710 13746
rect 1762 13694 1764 13746
rect 1708 13524 1764 13694
rect 1708 13458 1764 13468
rect 2380 13746 2436 13758
rect 2380 13694 2382 13746
rect 2434 13694 2436 13746
rect 2380 13412 2436 13694
rect 1932 13074 1988 13086
rect 1932 13022 1934 13074
rect 1986 13022 1988 13074
rect 1932 12180 1988 13022
rect 2380 12852 2436 13356
rect 3164 13634 3220 13646
rect 3164 13582 3166 13634
rect 3218 13582 3220 13634
rect 3164 13412 3220 13582
rect 3612 13634 3668 13646
rect 3612 13582 3614 13634
rect 3666 13582 3668 13634
rect 3612 13524 3668 13582
rect 3612 13458 3668 13468
rect 3164 13346 3220 13356
rect 5874 13356 6138 13366
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 5874 13290 6138 13300
rect 15198 13356 15462 13366
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15198 13290 15462 13300
rect 14700 13188 14756 13198
rect 4284 13076 4340 13086
rect 4284 12962 4340 13020
rect 4284 12910 4286 12962
rect 4338 12910 4340 12962
rect 4284 12898 4340 12910
rect 12684 12964 12740 12974
rect 2380 12786 2436 12796
rect 10536 12572 10800 12582
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10536 12506 10800 12516
rect 1932 12114 1988 12124
rect 4284 12180 4340 12190
rect 4284 12086 4340 12124
rect 1932 11954 1988 11966
rect 1932 11902 1934 11954
rect 1986 11902 1988 11954
rect 1932 11508 1988 11902
rect 5874 11788 6138 11798
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 5874 11722 6138 11732
rect 1932 11442 1988 11452
rect 10536 11004 10800 11014
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10536 10938 10800 10948
rect 5874 10220 6138 10230
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 5874 10154 6138 10164
rect 10536 9436 10800 9446
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10536 9370 10800 9380
rect 5874 8652 6138 8662
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 5874 8586 6138 8596
rect 10536 7868 10800 7878
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10536 7802 10800 7812
rect 5874 7084 6138 7094
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 5874 7018 6138 7028
rect 10536 6300 10800 6310
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10536 6234 10800 6244
rect 5874 5516 6138 5526
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 5874 5450 6138 5460
rect 10536 4732 10800 4742
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10536 4666 10800 4676
rect 12572 4116 12628 4126
rect 12460 4114 12628 4116
rect 12460 4062 12574 4114
rect 12626 4062 12628 4114
rect 12460 4060 12628 4062
rect 5874 3948 6138 3958
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 5874 3882 6138 3892
rect 12348 3554 12404 3566
rect 12348 3502 12350 3554
rect 12402 3502 12404 3554
rect 12012 3444 12068 3454
rect 12348 3444 12404 3502
rect 12012 3442 12348 3444
rect 12012 3390 12014 3442
rect 12066 3390 12348 3442
rect 12012 3388 12348 3390
rect 12012 3378 12068 3388
rect 12348 3378 12404 3388
rect 10536 3164 10800 3174
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10536 3098 10800 3108
rect 12460 980 12516 4060
rect 12572 4050 12628 4060
rect 12572 3444 12628 3454
rect 12684 3444 12740 12908
rect 13692 5124 13748 5134
rect 14364 5124 14420 5134
rect 13692 5122 14420 5124
rect 13692 5070 13694 5122
rect 13746 5070 14366 5122
rect 14418 5070 14420 5122
rect 13692 5068 14420 5070
rect 13692 5058 13748 5068
rect 14140 4900 14196 4910
rect 14140 4806 14196 4844
rect 14364 4228 14420 5068
rect 14700 5010 14756 13132
rect 15198 11788 15462 11798
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15198 11722 15462 11732
rect 15198 10220 15462 10230
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15198 10154 15462 10164
rect 15596 10164 15652 10174
rect 15198 8652 15462 8662
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15198 8586 15462 8596
rect 15198 7084 15462 7094
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15198 7018 15462 7028
rect 15198 5516 15462 5526
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15198 5450 15462 5460
rect 15596 5348 15652 10108
rect 15372 5292 15652 5348
rect 14700 4958 14702 5010
rect 14754 4958 14756 5010
rect 14700 4946 14756 4958
rect 14812 5124 14868 5134
rect 15036 5124 15092 5134
rect 14868 5122 15092 5124
rect 14868 5070 15038 5122
rect 15090 5070 15092 5122
rect 14868 5068 15092 5070
rect 14140 4172 14420 4228
rect 13356 3668 13412 3678
rect 12572 3442 12740 3444
rect 12572 3390 12574 3442
rect 12626 3390 12740 3442
rect 12572 3388 12740 3390
rect 13020 3666 13412 3668
rect 13020 3614 13358 3666
rect 13410 3614 13412 3666
rect 13020 3612 13412 3614
rect 12572 3378 12628 3388
rect 13020 980 13076 3612
rect 13356 3602 13412 3612
rect 12124 924 12516 980
rect 12796 924 13076 980
rect 13468 3444 13524 3454
rect 12124 800 12180 924
rect 12796 800 12852 924
rect 13468 800 13524 3388
rect 14140 800 14196 4172
rect 14812 800 14868 5068
rect 15036 5058 15092 5068
rect 15372 5010 15428 5292
rect 15372 4958 15374 5010
rect 15426 4958 15428 5010
rect 15372 4946 15428 4958
rect 14924 4340 14980 4350
rect 14924 4246 14980 4284
rect 15708 4338 15764 4350
rect 15708 4286 15710 4338
rect 15762 4286 15764 4338
rect 15484 4228 15540 4238
rect 15708 4228 15764 4286
rect 15484 4226 15764 4228
rect 15484 4174 15486 4226
rect 15538 4174 15764 4226
rect 15484 4172 15764 4174
rect 15484 4162 15540 4172
rect 15198 3948 15462 3958
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15198 3882 15462 3892
rect 15596 3388 15652 4172
rect 15708 3556 15764 3566
rect 15820 3556 15876 14252
rect 15932 12180 15988 18174
rect 16268 17892 16324 18510
rect 16828 18452 16884 19182
rect 16828 18386 16884 18396
rect 17388 18340 17444 18350
rect 17388 18246 17444 18284
rect 16268 17826 16324 17836
rect 16828 17890 16884 17902
rect 16828 17838 16830 17890
rect 16882 17838 16884 17890
rect 16604 17668 16660 17678
rect 16380 17666 16660 17668
rect 16380 17614 16606 17666
rect 16658 17614 16660 17666
rect 16380 17612 16660 17614
rect 16268 17444 16324 17454
rect 16268 16994 16324 17388
rect 16268 16942 16270 16994
rect 16322 16942 16324 16994
rect 16268 16930 16324 16942
rect 16380 15426 16436 17612
rect 16604 17602 16660 17612
rect 16380 15374 16382 15426
rect 16434 15374 16436 15426
rect 16380 15362 16436 15374
rect 16044 15316 16100 15326
rect 16044 15222 16100 15260
rect 16828 13076 16884 17838
rect 17724 17666 17780 22430
rect 17836 20188 17892 23102
rect 19180 23156 19236 23166
rect 19292 23156 19348 35756
rect 19404 35810 19460 35822
rect 19404 35758 19406 35810
rect 19458 35758 19460 35810
rect 19404 35364 19460 35758
rect 19404 35298 19460 35308
rect 19516 27860 19572 27870
rect 19516 27766 19572 27804
rect 19628 26908 19684 36204
rect 19740 35924 19796 36428
rect 19852 36418 19908 36428
rect 20748 36482 21140 36484
rect 20748 36430 21086 36482
rect 21138 36430 21140 36482
rect 20748 36428 21140 36430
rect 20188 36258 20244 36270
rect 20188 36206 20190 36258
rect 20242 36206 20244 36258
rect 19860 36092 20124 36102
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 19860 36026 20124 36036
rect 19852 35924 19908 35934
rect 19740 35922 19908 35924
rect 19740 35870 19854 35922
rect 19906 35870 19908 35922
rect 19740 35868 19908 35870
rect 19852 35858 19908 35868
rect 19860 34524 20124 34534
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 19860 34458 20124 34468
rect 19860 32956 20124 32966
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 19860 32890 20124 32900
rect 19860 31388 20124 31398
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 19860 31322 20124 31332
rect 19860 29820 20124 29830
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 19860 29754 20124 29764
rect 19860 28252 20124 28262
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 19860 28186 20124 28196
rect 19852 27970 19908 27982
rect 19852 27918 19854 27970
rect 19906 27918 19908 27970
rect 19852 27298 19908 27918
rect 19852 27246 19854 27298
rect 19906 27246 19908 27298
rect 19852 27234 19908 27246
rect 19516 26852 19684 26908
rect 19740 27074 19796 27086
rect 19740 27022 19742 27074
rect 19794 27022 19796 27074
rect 19516 26290 19572 26852
rect 19516 26238 19518 26290
rect 19570 26238 19572 26290
rect 19516 26226 19572 26238
rect 19628 26066 19684 26078
rect 19628 26014 19630 26066
rect 19682 26014 19684 26066
rect 19628 25506 19684 26014
rect 19628 25454 19630 25506
rect 19682 25454 19684 25506
rect 19628 25442 19684 25454
rect 19740 24724 19796 27022
rect 20188 27074 20244 36206
rect 20524 35698 20580 35710
rect 20524 35646 20526 35698
rect 20578 35646 20580 35698
rect 20524 28082 20580 35646
rect 20524 28030 20526 28082
rect 20578 28030 20580 28082
rect 20524 28018 20580 28030
rect 20636 32004 20692 32014
rect 20300 27970 20356 27982
rect 20300 27918 20302 27970
rect 20354 27918 20356 27970
rect 20300 27300 20356 27918
rect 20412 27300 20468 27310
rect 20636 27300 20692 31948
rect 20300 27244 20412 27300
rect 20412 27234 20468 27244
rect 20524 27244 20692 27300
rect 20188 27022 20190 27074
rect 20242 27022 20244 27074
rect 20188 27010 20244 27022
rect 20300 26964 20356 26974
rect 19860 26684 20124 26694
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 19860 26618 20124 26628
rect 20300 26516 20356 26908
rect 20076 26460 20356 26516
rect 20076 25394 20132 26460
rect 20076 25342 20078 25394
rect 20130 25342 20132 25394
rect 20076 25330 20132 25342
rect 20300 26290 20356 26302
rect 20300 26238 20302 26290
rect 20354 26238 20356 26290
rect 20188 25284 20244 25294
rect 19860 25116 20124 25126
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 19860 25050 20124 25060
rect 20188 24948 20244 25228
rect 19628 24498 19684 24510
rect 19628 24446 19630 24498
rect 19682 24446 19684 24498
rect 19628 23938 19684 24446
rect 19628 23886 19630 23938
rect 19682 23886 19684 23938
rect 19628 23874 19684 23886
rect 19180 23154 19348 23156
rect 19180 23102 19182 23154
rect 19234 23102 19348 23154
rect 19180 23100 19348 23102
rect 19740 23156 19796 24668
rect 20076 24892 20244 24948
rect 20076 23826 20132 24892
rect 20300 24724 20356 26238
rect 20300 24630 20356 24668
rect 20076 23774 20078 23826
rect 20130 23774 20132 23826
rect 20076 23762 20132 23774
rect 19860 23548 20124 23558
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 19860 23482 20124 23492
rect 20188 23268 20244 23278
rect 20076 23156 20132 23166
rect 20188 23156 20244 23212
rect 19740 23154 20020 23156
rect 19740 23102 19742 23154
rect 19794 23102 20020 23154
rect 19740 23100 20020 23102
rect 19180 23090 19236 23100
rect 19740 23090 19796 23100
rect 19068 22484 19124 22494
rect 18508 22370 18564 22382
rect 18508 22318 18510 22370
rect 18562 22318 18564 22370
rect 18508 21700 18564 22318
rect 17948 21476 18004 21486
rect 17948 21382 18004 21420
rect 18508 21474 18564 21644
rect 18508 21422 18510 21474
rect 18562 21422 18564 21474
rect 18508 21028 18564 21422
rect 18508 20962 18564 20972
rect 18956 21476 19012 21486
rect 18956 20802 19012 21420
rect 18956 20750 18958 20802
rect 19010 20750 19012 20802
rect 18284 20692 18340 20702
rect 18284 20598 18340 20636
rect 18620 20580 18676 20590
rect 17836 20132 18004 20188
rect 17724 17614 17726 17666
rect 17778 17614 17780 17666
rect 17724 17602 17780 17614
rect 17948 18450 18004 20132
rect 18172 20130 18228 20142
rect 18172 20078 18174 20130
rect 18226 20078 18228 20130
rect 18172 19234 18228 20078
rect 18172 19182 18174 19234
rect 18226 19182 18228 19234
rect 18172 19170 18228 19182
rect 18508 19124 18564 19134
rect 18508 19030 18564 19068
rect 18396 19010 18452 19022
rect 18396 18958 18398 19010
rect 18450 18958 18452 19010
rect 18396 18564 18452 18958
rect 18620 18788 18676 20524
rect 18956 20188 19012 20750
rect 18844 20132 19012 20188
rect 18732 19794 18788 19806
rect 18732 19742 18734 19794
rect 18786 19742 18788 19794
rect 18732 19236 18788 19742
rect 18732 19170 18788 19180
rect 18620 18732 18788 18788
rect 18620 18564 18676 18574
rect 18396 18508 18564 18564
rect 17948 18398 17950 18450
rect 18002 18398 18004 18450
rect 17948 16772 18004 18398
rect 18396 18340 18452 18350
rect 18284 18338 18452 18340
rect 18284 18286 18398 18338
rect 18450 18286 18452 18338
rect 18284 18284 18452 18286
rect 18172 17554 18228 17566
rect 18172 17502 18174 17554
rect 18226 17502 18228 17554
rect 17948 16706 18004 16716
rect 18060 17108 18116 17118
rect 18060 16882 18116 17052
rect 18060 16830 18062 16882
rect 18114 16830 18116 16882
rect 17388 16100 17444 16110
rect 17388 16006 17444 16044
rect 17948 16100 18004 16110
rect 17948 16006 18004 16044
rect 18060 15316 18116 16830
rect 18172 16098 18228 17502
rect 18172 16046 18174 16098
rect 18226 16046 18228 16098
rect 18172 16034 18228 16046
rect 18284 16100 18340 18284
rect 18396 18274 18452 18284
rect 18508 17556 18564 18508
rect 18284 16034 18340 16044
rect 18396 17500 18508 17556
rect 18396 15986 18452 17500
rect 18508 17490 18564 17500
rect 18620 17106 18676 18508
rect 18620 17054 18622 17106
rect 18674 17054 18676 17106
rect 18620 17042 18676 17054
rect 18508 16996 18564 17006
rect 18508 16098 18564 16940
rect 18732 16436 18788 18732
rect 18732 16370 18788 16380
rect 18844 16324 18900 20132
rect 18956 19460 19012 19470
rect 19068 19460 19124 22428
rect 19628 22484 19684 22494
rect 19964 22484 20020 23100
rect 20076 23154 20244 23156
rect 20076 23102 20078 23154
rect 20130 23102 20244 23154
rect 20076 23100 20244 23102
rect 20412 23154 20468 23166
rect 20412 23102 20414 23154
rect 20466 23102 20468 23154
rect 20076 23090 20132 23100
rect 20188 22930 20244 22942
rect 20188 22878 20190 22930
rect 20242 22878 20244 22930
rect 20076 22484 20132 22494
rect 19964 22482 20132 22484
rect 19964 22430 20078 22482
rect 20130 22430 20132 22482
rect 19964 22428 20132 22430
rect 19628 22370 19684 22428
rect 20076 22418 20132 22428
rect 19628 22318 19630 22370
rect 19682 22318 19684 22370
rect 19628 22306 19684 22318
rect 19516 22148 19572 22158
rect 19516 21586 19572 22092
rect 19860 21980 20124 21990
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 19860 21914 20124 21924
rect 19516 21534 19518 21586
rect 19570 21534 19572 21586
rect 19516 21522 19572 21534
rect 19740 21698 19796 21710
rect 19740 21646 19742 21698
rect 19794 21646 19796 21698
rect 19740 20188 19796 21646
rect 20076 21476 20132 21486
rect 20076 20802 20132 21420
rect 20188 21252 20244 22878
rect 20412 22594 20468 23102
rect 20412 22542 20414 22594
rect 20466 22542 20468 22594
rect 20412 22530 20468 22542
rect 20412 21700 20468 21710
rect 20412 21606 20468 21644
rect 20524 21586 20580 27244
rect 20636 27074 20692 27086
rect 20636 27022 20638 27074
rect 20690 27022 20692 27074
rect 20636 26180 20692 27022
rect 20636 26114 20692 26124
rect 20636 22148 20692 22158
rect 20636 22054 20692 22092
rect 20524 21534 20526 21586
rect 20578 21534 20580 21586
rect 20524 21522 20580 21534
rect 20300 21476 20356 21486
rect 20300 21382 20356 21420
rect 20188 21196 20356 21252
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 20076 20738 20132 20750
rect 20188 20804 20244 20814
rect 20300 20804 20356 21196
rect 20636 21028 20692 21038
rect 20748 21028 20804 36428
rect 21084 36418 21140 36428
rect 21420 35922 21476 36876
rect 21420 35870 21422 35922
rect 21474 35870 21476 35922
rect 21420 35858 21476 35870
rect 20860 35364 20916 35374
rect 20860 26908 20916 35308
rect 21532 35028 21588 39200
rect 22092 36708 22148 36718
rect 22092 36614 22148 36652
rect 22204 35812 22260 39200
rect 22876 36484 22932 39200
rect 23548 36596 23604 39200
rect 24220 36820 24276 39200
rect 24522 36876 24786 36886
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24522 36810 24786 36820
rect 24220 36754 24276 36764
rect 24892 36596 24948 39200
rect 25564 36820 25620 39200
rect 26236 36932 26292 39200
rect 26236 36866 26292 36876
rect 26908 36820 26964 39200
rect 27468 36932 27524 36942
rect 25564 36764 26180 36820
rect 26908 36764 27076 36820
rect 23548 36540 24276 36596
rect 22876 36418 22932 36428
rect 22204 35746 22260 35756
rect 23100 35812 23156 35822
rect 22764 35700 22820 35710
rect 21532 35026 21812 35028
rect 21532 34974 21534 35026
rect 21586 34974 21812 35026
rect 21532 34972 21812 34974
rect 21532 34962 21588 34972
rect 21756 34914 21812 34972
rect 21756 34862 21758 34914
rect 21810 34862 21812 34914
rect 21756 34850 21812 34862
rect 22652 34916 22708 34926
rect 22092 34690 22148 34702
rect 22092 34638 22094 34690
rect 22146 34638 22148 34690
rect 21868 32340 21924 32350
rect 21084 27300 21140 27310
rect 20860 26852 21028 26908
rect 20972 26516 21028 26852
rect 20860 26460 21028 26516
rect 20860 22594 20916 26460
rect 20972 26292 21028 26302
rect 20972 26198 21028 26236
rect 20972 24724 21028 24734
rect 20972 24630 21028 24668
rect 21084 23940 21140 27244
rect 21308 26964 21364 27002
rect 21308 26898 21364 26908
rect 21644 26962 21700 26974
rect 21644 26910 21646 26962
rect 21698 26910 21700 26962
rect 21532 26850 21588 26862
rect 21532 26798 21534 26850
rect 21586 26798 21588 26850
rect 21420 26180 21476 26190
rect 21420 26086 21476 26124
rect 21532 25620 21588 26798
rect 21420 25564 21588 25620
rect 21420 25396 21476 25564
rect 21308 25394 21476 25396
rect 21308 25342 21422 25394
rect 21474 25342 21476 25394
rect 21308 25340 21476 25342
rect 21196 25284 21252 25294
rect 21196 25190 21252 25228
rect 21308 24948 21364 25340
rect 21420 25330 21476 25340
rect 21532 25396 21588 25406
rect 21532 25302 21588 25340
rect 21644 25284 21700 26910
rect 21644 25218 21700 25228
rect 21756 26180 21812 26190
rect 21196 23940 21252 23950
rect 21084 23938 21252 23940
rect 21084 23886 21198 23938
rect 21250 23886 21252 23938
rect 21084 23884 21252 23886
rect 21196 23874 21252 23884
rect 21308 23828 21364 24892
rect 21756 24610 21812 26124
rect 21868 25618 21924 32284
rect 22092 32004 22148 34638
rect 22092 31938 22148 31948
rect 22204 31556 22260 31566
rect 22652 31556 22708 34860
rect 21868 25566 21870 25618
rect 21922 25566 21924 25618
rect 21868 25554 21924 25566
rect 21980 31500 22204 31556
rect 21756 24558 21758 24610
rect 21810 24558 21812 24610
rect 21420 23828 21476 23838
rect 21308 23826 21476 23828
rect 21308 23774 21422 23826
rect 21474 23774 21476 23826
rect 21308 23772 21476 23774
rect 21420 23378 21476 23772
rect 21420 23326 21422 23378
rect 21474 23326 21476 23378
rect 21420 23314 21476 23326
rect 21532 23826 21588 23838
rect 21532 23774 21534 23826
rect 21586 23774 21588 23826
rect 21532 23380 21588 23774
rect 21532 23314 21588 23324
rect 21756 23268 21812 24558
rect 21868 24052 21924 24062
rect 21980 24052 22036 31500
rect 22204 31490 22260 31500
rect 22540 31500 22708 31556
rect 22540 26908 22596 31500
rect 22540 26852 22708 26908
rect 21868 24050 22036 24052
rect 21868 23998 21870 24050
rect 21922 23998 22036 24050
rect 21868 23996 22036 23998
rect 22204 25506 22260 25518
rect 22204 25454 22206 25506
rect 22258 25454 22260 25506
rect 21868 23986 21924 23996
rect 22204 23940 22260 25454
rect 22652 25506 22708 26852
rect 22652 25454 22654 25506
rect 22706 25454 22708 25506
rect 22652 25442 22708 25454
rect 21756 23202 21812 23212
rect 22092 23938 22260 23940
rect 22092 23886 22206 23938
rect 22258 23886 22260 23938
rect 22092 23884 22260 23886
rect 21084 23156 21140 23166
rect 20860 22542 20862 22594
rect 20914 22542 20916 22594
rect 20860 22530 20916 22542
rect 20972 23154 21140 23156
rect 20972 23102 21086 23154
rect 21138 23102 21140 23154
rect 20972 23100 21140 23102
rect 20636 21026 20804 21028
rect 20636 20974 20638 21026
rect 20690 20974 20804 21026
rect 20636 20972 20804 20974
rect 20860 22148 20916 22158
rect 20636 20962 20692 20972
rect 20524 20804 20580 20814
rect 20300 20802 20580 20804
rect 20300 20750 20526 20802
rect 20578 20750 20580 20802
rect 20300 20748 20580 20750
rect 20188 20710 20244 20748
rect 20524 20738 20580 20748
rect 19860 20412 20124 20422
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 19860 20346 20124 20356
rect 19404 20132 19796 20188
rect 19292 20018 19348 20030
rect 19292 19966 19294 20018
rect 19346 19966 19348 20018
rect 18956 19458 19124 19460
rect 18956 19406 18958 19458
rect 19010 19406 19124 19458
rect 18956 19404 19124 19406
rect 19180 19906 19236 19918
rect 19180 19854 19182 19906
rect 19234 19854 19236 19906
rect 18956 19394 19012 19404
rect 19180 18676 19236 19854
rect 19292 19460 19348 19966
rect 19292 19394 19348 19404
rect 19404 19234 19460 20132
rect 19740 20066 19796 20076
rect 19964 20244 20020 20254
rect 19404 19182 19406 19234
rect 19458 19182 19460 19234
rect 19404 19170 19460 19182
rect 19628 19236 19684 19246
rect 19628 19142 19684 19180
rect 19964 19124 20020 20188
rect 20300 20132 20356 20142
rect 20300 19234 20356 20076
rect 20300 19182 20302 19234
rect 20354 19182 20356 19234
rect 20300 19170 20356 19182
rect 20412 19348 20468 19358
rect 19740 19122 20020 19124
rect 19740 19070 19966 19122
rect 20018 19070 20020 19122
rect 19740 19068 20020 19070
rect 19740 18788 19796 19068
rect 19964 19058 20020 19068
rect 19180 18610 19236 18620
rect 19404 18732 19796 18788
rect 19860 18844 20124 18854
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 19860 18778 20124 18788
rect 18956 18452 19012 18462
rect 18956 18358 19012 18396
rect 19292 18338 19348 18350
rect 19292 18286 19294 18338
rect 19346 18286 19348 18338
rect 19292 18228 19348 18286
rect 19292 18162 19348 18172
rect 19404 17668 19460 18732
rect 19740 18564 19796 18574
rect 19740 18450 19796 18508
rect 19740 18398 19742 18450
rect 19794 18398 19796 18450
rect 19740 18386 19796 18398
rect 20412 18452 20468 19292
rect 20860 19348 20916 22092
rect 20972 20244 21028 23100
rect 21084 23090 21140 23100
rect 21532 22258 21588 22270
rect 21532 22206 21534 22258
rect 21586 22206 21588 22258
rect 21196 22148 21252 22158
rect 21420 22148 21476 22158
rect 21084 22146 21252 22148
rect 21084 22094 21198 22146
rect 21250 22094 21252 22146
rect 21084 22092 21252 22094
rect 21084 21698 21140 22092
rect 21196 22082 21252 22092
rect 21308 22146 21476 22148
rect 21308 22094 21422 22146
rect 21474 22094 21476 22146
rect 21308 22092 21476 22094
rect 21084 21646 21086 21698
rect 21138 21646 21140 21698
rect 21084 21634 21140 21646
rect 21196 20804 21252 20814
rect 21196 20578 21252 20748
rect 21196 20526 21198 20578
rect 21250 20526 21252 20578
rect 21196 20514 21252 20526
rect 21308 20802 21364 22092
rect 21420 22082 21476 22092
rect 21532 22148 21588 22206
rect 21532 22082 21588 22092
rect 21868 22258 21924 22270
rect 21868 22206 21870 22258
rect 21922 22206 21924 22258
rect 21308 20750 21310 20802
rect 21362 20750 21364 20802
rect 21308 20356 21364 20750
rect 21196 20300 21364 20356
rect 21420 21586 21476 21598
rect 21420 21534 21422 21586
rect 21474 21534 21476 21586
rect 21420 20692 21476 21534
rect 21196 20188 21252 20300
rect 20972 20178 21028 20188
rect 20860 19282 20916 19292
rect 21084 20132 21252 20188
rect 20412 18358 20468 18396
rect 21084 19236 21140 20132
rect 21084 18338 21140 19180
rect 21308 20130 21364 20142
rect 21308 20078 21310 20130
rect 21362 20078 21364 20130
rect 21308 18452 21364 20078
rect 21420 19236 21476 20636
rect 21756 20188 21812 20198
rect 21756 20130 21812 20132
rect 21756 20078 21758 20130
rect 21810 20078 21812 20130
rect 21756 20066 21812 20078
rect 21532 20018 21588 20030
rect 21532 19966 21534 20018
rect 21586 19966 21588 20018
rect 21532 19796 21588 19966
rect 21532 19730 21588 19740
rect 21644 20020 21700 20030
rect 21644 19572 21700 19964
rect 21868 19908 21924 22206
rect 21980 22260 22036 22270
rect 22092 22260 22148 23884
rect 22204 23874 22260 23884
rect 22540 25284 22596 25294
rect 22540 23716 22596 25228
rect 22652 24836 22708 24846
rect 22652 24742 22708 24780
rect 22764 23938 22820 35644
rect 23100 35026 23156 35756
rect 23100 34974 23102 35026
rect 23154 34974 23156 35026
rect 23100 34962 23156 34974
rect 23324 35810 23380 35822
rect 23324 35758 23326 35810
rect 23378 35758 23380 35810
rect 23324 31556 23380 35758
rect 23548 35812 23604 35822
rect 23548 35698 23604 35756
rect 23548 35646 23550 35698
rect 23602 35646 23604 35698
rect 23548 35634 23604 35646
rect 23772 35026 23828 36540
rect 23996 35812 24052 35822
rect 23996 35718 24052 35756
rect 24220 35698 24276 36540
rect 24892 36530 24948 36540
rect 25452 36708 25508 36718
rect 26124 36708 26180 36764
rect 26124 36652 26852 36708
rect 24780 36484 24836 36494
rect 24556 36260 24612 36270
rect 24220 35646 24222 35698
rect 24274 35646 24276 35698
rect 24220 35634 24276 35646
rect 24332 36258 24612 36260
rect 24332 36206 24558 36258
rect 24610 36206 24612 36258
rect 24332 36204 24612 36206
rect 23772 34974 23774 35026
rect 23826 34974 23828 35026
rect 23772 34962 23828 34974
rect 24220 35476 24276 35486
rect 23324 31490 23380 31500
rect 23996 33460 24052 33470
rect 23436 25506 23492 25518
rect 23436 25454 23438 25506
rect 23490 25454 23492 25506
rect 22876 25396 22932 25406
rect 22876 25302 22932 25340
rect 22876 24948 22932 24958
rect 22876 24854 22932 24892
rect 22988 24836 23044 24846
rect 22988 24742 23044 24780
rect 22764 23886 22766 23938
rect 22818 23886 22820 23938
rect 22764 23874 22820 23886
rect 23436 23938 23492 25454
rect 23996 25506 24052 33404
rect 24220 26908 24276 35420
rect 24332 34916 24388 36204
rect 24556 36194 24612 36204
rect 24780 35476 24836 36428
rect 25452 36482 25508 36652
rect 26236 36484 26292 36494
rect 25452 36430 25454 36482
rect 25506 36430 25508 36482
rect 25004 36260 25060 36270
rect 24780 35420 24948 35476
rect 24522 35308 24786 35318
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24522 35242 24786 35252
rect 24892 35140 24948 35420
rect 24332 34850 24388 34860
rect 24444 35084 24948 35140
rect 24332 34692 24388 34702
rect 24444 34692 24500 35084
rect 24332 34690 24500 34692
rect 24332 34638 24334 34690
rect 24386 34638 24500 34690
rect 24332 34636 24500 34638
rect 24332 34626 24388 34636
rect 24522 33740 24786 33750
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24522 33674 24786 33684
rect 24892 33572 24948 33582
rect 24522 32172 24786 32182
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24522 32106 24786 32116
rect 24522 30604 24786 30614
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24522 30538 24786 30548
rect 24522 29036 24786 29046
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24522 28970 24786 28980
rect 24522 27468 24786 27478
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24522 27402 24786 27412
rect 23996 25454 23998 25506
rect 24050 25454 24052 25506
rect 23996 25442 24052 25454
rect 24108 26852 24276 26908
rect 23436 23886 23438 23938
rect 23490 23886 23492 23938
rect 22876 23716 22932 23726
rect 22540 23714 22932 23716
rect 22540 23662 22878 23714
rect 22930 23662 22932 23714
rect 22540 23660 22932 23662
rect 22876 23650 22932 23660
rect 23436 23268 23492 23886
rect 24108 23938 24164 26852
rect 24522 25900 24786 25910
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24522 25834 24786 25844
rect 24892 25506 24948 33516
rect 24892 25454 24894 25506
rect 24946 25454 24948 25506
rect 24892 25442 24948 25454
rect 24522 24332 24786 24342
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24522 24266 24786 24276
rect 24108 23886 24110 23938
rect 24162 23886 24164 23938
rect 24108 23874 24164 23886
rect 25004 23938 25060 36204
rect 25228 36258 25284 36270
rect 25228 36206 25230 36258
rect 25282 36206 25284 36258
rect 25228 35476 25284 36206
rect 25452 35922 25508 36430
rect 26012 36428 26236 36484
rect 25900 36260 25956 36270
rect 25452 35870 25454 35922
rect 25506 35870 25508 35922
rect 25452 35858 25508 35870
rect 25788 36258 25956 36260
rect 25788 36206 25902 36258
rect 25954 36206 25956 36258
rect 25788 36204 25956 36206
rect 25228 35410 25284 35420
rect 25788 32340 25844 36204
rect 25900 36194 25956 36204
rect 25900 35924 25956 35934
rect 26012 35924 26068 36428
rect 26236 36390 26292 36428
rect 25900 35922 26068 35924
rect 25900 35870 25902 35922
rect 25954 35870 26068 35922
rect 25900 35868 26068 35870
rect 26348 35922 26404 36652
rect 26796 36482 26852 36652
rect 26796 36430 26798 36482
rect 26850 36430 26852 36482
rect 26796 36418 26852 36430
rect 26572 36260 26628 36270
rect 26572 36166 26628 36204
rect 27020 36036 27076 36764
rect 27468 36482 27524 36876
rect 28476 36932 28532 36942
rect 28476 36594 28532 36876
rect 33846 36876 34110 36886
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 33846 36810 34110 36820
rect 28476 36542 28478 36594
rect 28530 36542 28532 36594
rect 28476 36530 28532 36542
rect 27468 36430 27470 36482
rect 27522 36430 27524 36482
rect 27468 36418 27524 36430
rect 27244 36260 27300 36270
rect 27244 36258 27524 36260
rect 27244 36206 27246 36258
rect 27298 36206 27524 36258
rect 27244 36204 27524 36206
rect 27244 36194 27300 36204
rect 27020 35980 27412 36036
rect 26348 35870 26350 35922
rect 26402 35870 26404 35922
rect 25900 35858 25956 35868
rect 26348 35858 26404 35870
rect 26908 35924 26964 35934
rect 27020 35924 27076 35980
rect 26908 35922 27076 35924
rect 26908 35870 26910 35922
rect 26962 35870 27076 35922
rect 26908 35868 27076 35870
rect 26908 35858 26964 35868
rect 27132 35810 27188 35822
rect 27132 35758 27134 35810
rect 27186 35758 27188 35810
rect 27132 33460 27188 35758
rect 27356 35698 27412 35980
rect 27356 35646 27358 35698
rect 27410 35646 27412 35698
rect 27356 35634 27412 35646
rect 27468 33572 27524 36204
rect 29184 36092 29448 36102
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29184 36026 29448 36036
rect 38508 36092 38772 36102
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38508 36026 38772 36036
rect 33846 35308 34110 35318
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 33846 35242 34110 35252
rect 29184 34524 29448 34534
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29184 34458 29448 34468
rect 38508 34524 38772 34534
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38508 34458 38772 34468
rect 33846 33740 34110 33750
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 33846 33674 34110 33684
rect 27468 33506 27524 33516
rect 27132 33394 27188 33404
rect 29184 32956 29448 32966
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29184 32890 29448 32900
rect 38508 32956 38772 32966
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38508 32890 38772 32900
rect 25788 32274 25844 32284
rect 33846 32172 34110 32182
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 33846 32106 34110 32116
rect 29184 31388 29448 31398
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29184 31322 29448 31332
rect 38508 31388 38772 31398
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38508 31322 38772 31332
rect 37884 31108 37940 31118
rect 37324 31106 37940 31108
rect 37324 31054 37886 31106
rect 37938 31054 37940 31106
rect 37324 31052 37940 31054
rect 33846 30604 34110 30614
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 33846 30538 34110 30548
rect 29184 29820 29448 29830
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29184 29754 29448 29764
rect 33846 29036 34110 29046
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 33846 28970 34110 28980
rect 28700 28756 28756 28766
rect 26460 25284 26516 25294
rect 25900 24724 25956 24734
rect 25676 24722 25956 24724
rect 25676 24670 25902 24722
rect 25954 24670 25956 24722
rect 25676 24668 25956 24670
rect 25564 24612 25620 24622
rect 25564 24518 25620 24556
rect 25004 23886 25006 23938
rect 25058 23886 25060 23938
rect 25004 23874 25060 23886
rect 23548 23268 23604 23278
rect 23436 23212 23548 23268
rect 23548 23174 23604 23212
rect 22036 22204 22148 22260
rect 23324 23154 23380 23166
rect 23324 23102 23326 23154
rect 23378 23102 23380 23154
rect 21980 22166 22036 22204
rect 22204 22148 22260 22158
rect 22260 22092 22372 22148
rect 22204 22054 22260 22092
rect 22092 21588 22148 21598
rect 21980 21586 22148 21588
rect 21980 21534 22094 21586
rect 22146 21534 22148 21586
rect 21980 21532 22148 21534
rect 21980 19908 22036 21532
rect 22092 21522 22148 21532
rect 22316 20802 22372 22092
rect 22316 20750 22318 20802
rect 22370 20750 22372 20802
rect 22316 20738 22372 20750
rect 22876 21474 22932 21486
rect 22876 21422 22878 21474
rect 22930 21422 22932 21474
rect 22540 20690 22596 20702
rect 22540 20638 22542 20690
rect 22594 20638 22596 20690
rect 22540 20356 22596 20638
rect 22092 20300 22596 20356
rect 22764 20356 22820 20366
rect 22092 20242 22148 20300
rect 22092 20190 22094 20242
rect 22146 20190 22148 20242
rect 22092 20178 22148 20190
rect 22764 20188 22820 20300
rect 22540 20132 22820 20188
rect 22876 20132 22932 21422
rect 23212 21476 23268 21486
rect 23212 21382 23268 21420
rect 23100 20692 23156 20702
rect 23100 20598 23156 20636
rect 23324 20188 23380 23102
rect 25452 23044 25508 23054
rect 25452 22950 25508 22988
rect 24522 22764 24786 22774
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24522 22698 24786 22708
rect 23436 22146 23492 22158
rect 23436 22094 23438 22146
rect 23490 22094 23492 22146
rect 23436 21476 23492 22094
rect 24220 22146 24276 22158
rect 24220 22094 24222 22146
rect 24274 22094 24276 22146
rect 24220 21924 24276 22094
rect 23436 21410 23492 21420
rect 23772 21868 24276 21924
rect 23772 21586 23828 21868
rect 23996 21700 24052 21710
rect 23772 21534 23774 21586
rect 23826 21534 23828 21586
rect 23772 21476 23828 21534
rect 23772 21028 23828 21420
rect 23772 20962 23828 20972
rect 23884 21698 24052 21700
rect 23884 21646 23998 21698
rect 24050 21646 24052 21698
rect 23884 21644 24052 21646
rect 23436 20802 23492 20814
rect 23436 20750 23438 20802
rect 23490 20750 23492 20802
rect 23436 20692 23492 20750
rect 23436 20626 23492 20636
rect 23884 20188 23940 21644
rect 23996 21634 24052 21644
rect 25228 21586 25284 21598
rect 25228 21534 25230 21586
rect 25282 21534 25284 21586
rect 24444 21476 24500 21486
rect 24444 21382 24500 21420
rect 25004 21476 25060 21486
rect 24332 21364 24388 21374
rect 24220 21362 24388 21364
rect 24220 21310 24334 21362
rect 24386 21310 24388 21362
rect 24220 21308 24388 21310
rect 23996 20690 24052 20702
rect 23996 20638 23998 20690
rect 24050 20638 24052 20690
rect 23996 20580 24052 20638
rect 23996 20514 24052 20524
rect 22540 20130 22596 20132
rect 22540 20078 22542 20130
rect 22594 20078 22596 20130
rect 22540 20066 22596 20078
rect 22876 20066 22932 20076
rect 23212 20132 23268 20142
rect 23324 20132 23828 20188
rect 23884 20132 24052 20188
rect 22652 20018 22708 20030
rect 22652 19966 22654 20018
rect 22706 19966 22708 20018
rect 21980 19852 22148 19908
rect 21868 19796 21924 19852
rect 21644 19506 21700 19516
rect 21756 19740 21924 19796
rect 21644 19236 21700 19246
rect 21420 19234 21700 19236
rect 21420 19182 21646 19234
rect 21698 19182 21700 19234
rect 21420 19180 21700 19182
rect 21644 19170 21700 19180
rect 21532 18452 21588 18462
rect 21308 18396 21532 18452
rect 21532 18358 21588 18396
rect 21084 18286 21086 18338
rect 21138 18286 21140 18338
rect 19180 17666 19460 17668
rect 19180 17614 19406 17666
rect 19458 17614 19460 17666
rect 19180 17612 19460 17614
rect 19068 17556 19124 17566
rect 19068 17462 19124 17500
rect 19068 16996 19124 17006
rect 19180 16996 19236 17612
rect 19404 17602 19460 17612
rect 19628 17892 19684 17902
rect 19628 17666 19684 17836
rect 19628 17614 19630 17666
rect 19682 17614 19684 17666
rect 19628 17602 19684 17614
rect 19964 17668 20020 17678
rect 19964 17574 20020 17612
rect 19852 17556 19908 17566
rect 19852 17462 19908 17500
rect 20412 17556 20468 17566
rect 20412 17462 20468 17500
rect 20524 17554 20580 17566
rect 20524 17502 20526 17554
rect 20578 17502 20580 17554
rect 20188 17444 20244 17454
rect 20188 17350 20244 17388
rect 19860 17276 20124 17286
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 19860 17210 20124 17220
rect 20524 17220 20580 17502
rect 20524 17154 20580 17164
rect 19740 17108 19796 17118
rect 19740 17014 19796 17052
rect 20412 17108 20468 17118
rect 19068 16994 19236 16996
rect 19068 16942 19070 16994
rect 19122 16942 19236 16994
rect 19068 16940 19236 16942
rect 19068 16930 19124 16940
rect 19180 16884 19236 16940
rect 19180 16818 19236 16828
rect 19964 16884 20020 16894
rect 19964 16790 20020 16828
rect 20188 16884 20244 16894
rect 20188 16882 20356 16884
rect 20188 16830 20190 16882
rect 20242 16830 20356 16882
rect 20188 16828 20356 16830
rect 20188 16818 20244 16828
rect 18956 16772 19012 16782
rect 18956 16678 19012 16716
rect 19292 16772 19348 16782
rect 19292 16678 19348 16716
rect 19628 16660 19684 16670
rect 19404 16658 19684 16660
rect 19404 16606 19630 16658
rect 19682 16606 19684 16658
rect 19404 16604 19684 16606
rect 19068 16436 19124 16446
rect 18844 16268 19012 16324
rect 18844 16100 18900 16110
rect 18508 16046 18510 16098
rect 18562 16046 18564 16098
rect 18508 16034 18564 16046
rect 18732 16098 18900 16100
rect 18732 16046 18846 16098
rect 18898 16046 18900 16098
rect 18732 16044 18900 16046
rect 18396 15934 18398 15986
rect 18450 15934 18452 15986
rect 18396 15922 18452 15934
rect 18060 15250 18116 15260
rect 18620 15316 18676 15326
rect 18620 15222 18676 15260
rect 18396 15090 18452 15102
rect 18396 15038 18398 15090
rect 18450 15038 18452 15090
rect 18060 14532 18116 14542
rect 17948 13972 18004 13982
rect 17948 13878 18004 13916
rect 18060 13970 18116 14476
rect 18060 13918 18062 13970
rect 18114 13918 18116 13970
rect 18060 13906 18116 13918
rect 16828 13010 16884 13020
rect 17836 13746 17892 13758
rect 17836 13694 17838 13746
rect 17890 13694 17892 13746
rect 17836 12852 17892 13694
rect 18284 13636 18340 13646
rect 18284 13542 18340 13580
rect 17836 12786 17892 12796
rect 15932 12114 15988 12124
rect 18060 11844 18116 11854
rect 16604 4900 16660 4910
rect 16156 4898 16660 4900
rect 16156 4846 16606 4898
rect 16658 4846 16660 4898
rect 16156 4844 16660 4846
rect 16044 4564 16100 4574
rect 16044 4470 16100 4508
rect 15708 3554 15876 3556
rect 15708 3502 15710 3554
rect 15762 3502 15876 3554
rect 15708 3500 15876 3502
rect 16156 3554 16212 4844
rect 16604 4834 16660 4844
rect 16156 3502 16158 3554
rect 16210 3502 16212 3554
rect 15708 3490 15764 3500
rect 15484 3332 15652 3388
rect 15484 800 15540 3332
rect 16156 800 16212 3502
rect 16380 4676 16436 4686
rect 16380 3330 16436 4620
rect 16380 3278 16382 3330
rect 16434 3278 16436 3330
rect 16380 3266 16436 3278
rect 16828 4226 16884 4238
rect 16828 4174 16830 4226
rect 16882 4174 16884 4226
rect 16828 3556 16884 4174
rect 17612 4226 17668 4238
rect 17612 4174 17614 4226
rect 17666 4174 17668 4226
rect 17052 3556 17108 3566
rect 16828 3554 17108 3556
rect 16828 3502 17054 3554
rect 17106 3502 17108 3554
rect 16828 3500 17108 3502
rect 16828 800 16884 3500
rect 17052 3490 17108 3500
rect 17612 3556 17668 4174
rect 17724 3556 17780 3566
rect 17612 3554 17780 3556
rect 17612 3502 17726 3554
rect 17778 3502 17780 3554
rect 17612 3500 17780 3502
rect 17388 3444 17444 3482
rect 17612 3388 17668 3500
rect 17724 3490 17780 3500
rect 17388 3378 17444 3388
rect 17500 3332 17668 3388
rect 18060 3442 18116 11788
rect 18060 3390 18062 3442
rect 18114 3390 18116 3442
rect 18060 3378 18116 3390
rect 18172 4226 18228 4238
rect 18172 4174 18174 4226
rect 18226 4174 18228 4226
rect 18172 3556 18228 4174
rect 17500 800 17556 3332
rect 18172 800 18228 3500
rect 18396 3442 18452 15038
rect 18620 14980 18676 14990
rect 18508 13524 18564 13534
rect 18508 13430 18564 13468
rect 18620 4676 18676 14924
rect 18732 11844 18788 16044
rect 18844 16034 18900 16044
rect 18956 15876 19012 16268
rect 18956 15810 19012 15820
rect 19068 15538 19124 16380
rect 19404 16324 19460 16604
rect 19628 16594 19684 16604
rect 19068 15486 19070 15538
rect 19122 15486 19124 15538
rect 19068 15474 19124 15486
rect 19180 16268 19460 16324
rect 19516 16436 19572 16446
rect 19180 16098 19236 16268
rect 19180 16046 19182 16098
rect 19234 16046 19236 16098
rect 18844 15314 18900 15326
rect 18844 15262 18846 15314
rect 18898 15262 18900 15314
rect 18844 12180 18900 15262
rect 19180 15316 19236 16046
rect 19516 16098 19572 16380
rect 19516 16046 19518 16098
rect 19570 16046 19572 16098
rect 19516 16034 19572 16046
rect 19740 16100 19796 16110
rect 19180 15250 19236 15260
rect 19292 15874 19348 15886
rect 19292 15822 19294 15874
rect 19346 15822 19348 15874
rect 18956 15202 19012 15214
rect 18956 15150 18958 15202
rect 19010 15150 19012 15202
rect 18956 14420 19012 15150
rect 19292 14980 19348 15822
rect 19292 14914 19348 14924
rect 19404 15874 19460 15886
rect 19404 15822 19406 15874
rect 19458 15822 19460 15874
rect 19404 14868 19460 15822
rect 19516 15876 19572 15886
rect 19516 15428 19572 15820
rect 19516 15426 19684 15428
rect 19516 15374 19518 15426
rect 19570 15374 19684 15426
rect 19516 15372 19684 15374
rect 19516 15362 19572 15372
rect 19404 14802 19460 14812
rect 19516 14532 19572 14542
rect 19404 14530 19572 14532
rect 19404 14478 19518 14530
rect 19570 14478 19572 14530
rect 19404 14476 19572 14478
rect 19404 14420 19460 14476
rect 19516 14466 19572 14476
rect 18956 14364 19460 14420
rect 19628 14420 19684 15372
rect 19628 14354 19684 14364
rect 19740 13746 19796 16044
rect 19860 15708 20124 15718
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 19860 15642 20124 15652
rect 20076 15316 20132 15326
rect 20076 15222 20132 15260
rect 20188 15204 20244 15214
rect 20188 15110 20244 15148
rect 20188 14644 20244 14654
rect 19964 14420 20020 14430
rect 19964 14326 20020 14364
rect 19860 14140 20124 14150
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 19860 14074 20124 14084
rect 19740 13694 19742 13746
rect 19794 13694 19796 13746
rect 18956 13636 19012 13646
rect 18956 13542 19012 13580
rect 19292 13522 19348 13534
rect 19292 13470 19294 13522
rect 19346 13470 19348 13522
rect 19292 13188 19348 13470
rect 19292 13122 19348 13132
rect 19292 12964 19348 12974
rect 19292 12870 19348 12908
rect 19740 12962 19796 13694
rect 20076 13858 20132 13870
rect 20076 13806 20078 13858
rect 20130 13806 20132 13858
rect 20076 13076 20132 13806
rect 20188 13300 20244 14588
rect 20300 13524 20356 16828
rect 20412 14532 20468 17052
rect 20524 16996 20580 17006
rect 21084 16996 21140 18286
rect 21644 17668 21700 17678
rect 21756 17668 21812 19740
rect 21868 19572 21924 19582
rect 21868 19122 21924 19516
rect 22092 19572 22148 19852
rect 22652 19796 22708 19966
rect 22764 20020 22820 20030
rect 22764 19926 22820 19964
rect 23100 19796 23156 19806
rect 22092 19506 22148 19516
rect 22204 19794 23156 19796
rect 22204 19742 23102 19794
rect 23154 19742 23156 19794
rect 22204 19740 23156 19742
rect 21980 19236 22036 19246
rect 22204 19236 22260 19740
rect 23100 19730 23156 19740
rect 21980 19234 22260 19236
rect 21980 19182 21982 19234
rect 22034 19182 22260 19234
rect 21980 19180 22260 19182
rect 21980 19170 22036 19180
rect 21868 19070 21870 19122
rect 21922 19070 21924 19122
rect 21868 19058 21924 19070
rect 23212 18676 23268 20076
rect 23436 20018 23492 20030
rect 23436 19966 23438 20018
rect 23490 19966 23492 20018
rect 23324 19908 23380 19918
rect 23436 19908 23492 19966
rect 23772 20020 23828 20132
rect 23772 20018 23940 20020
rect 23772 19966 23774 20018
rect 23826 19966 23940 20018
rect 23772 19964 23940 19966
rect 23772 19954 23828 19964
rect 23380 19852 23492 19908
rect 23324 19842 23380 19852
rect 23548 19796 23604 19806
rect 23212 18610 23268 18620
rect 23436 19740 23548 19796
rect 21644 17666 21812 17668
rect 21644 17614 21646 17666
rect 21698 17614 21812 17666
rect 21644 17612 21812 17614
rect 22204 18562 22260 18574
rect 22204 18510 22206 18562
rect 22258 18510 22260 18562
rect 21644 17602 21700 17612
rect 21308 17442 21364 17454
rect 21308 17390 21310 17442
rect 21362 17390 21364 17442
rect 21308 17108 21364 17390
rect 22204 17444 22260 18510
rect 22540 18450 22596 18462
rect 22540 18398 22542 18450
rect 22594 18398 22596 18450
rect 22540 18340 22596 18398
rect 22876 18452 22932 18462
rect 22876 18358 22932 18396
rect 22540 18274 22596 18284
rect 22988 18340 23044 18350
rect 22988 18246 23044 18284
rect 22988 17666 23044 17678
rect 22988 17614 22990 17666
rect 23042 17614 23044 17666
rect 22204 17378 22260 17388
rect 22316 17442 22372 17454
rect 22316 17390 22318 17442
rect 22370 17390 22372 17442
rect 22092 17108 22148 17118
rect 22316 17108 22372 17390
rect 22652 17444 22708 17454
rect 22652 17350 22708 17388
rect 21308 17042 21364 17052
rect 21868 17052 22092 17108
rect 20524 16994 21140 16996
rect 20524 16942 20526 16994
rect 20578 16942 21140 16994
rect 20524 16940 21140 16942
rect 20524 16930 20580 16940
rect 21868 16882 21924 17052
rect 22092 17042 22148 17052
rect 22204 17052 22372 17108
rect 22988 17108 23044 17614
rect 23436 17666 23492 19740
rect 23548 19730 23604 19740
rect 23436 17614 23438 17666
rect 23490 17614 23492 17666
rect 23436 17602 23492 17614
rect 23884 17444 23940 19964
rect 23996 19908 24052 20132
rect 24220 20132 24276 21308
rect 24332 21298 24388 21308
rect 24522 21196 24786 21206
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24522 21130 24786 21140
rect 24332 21028 24388 21038
rect 24332 20802 24388 20972
rect 24332 20750 24334 20802
rect 24386 20750 24388 20802
rect 24332 20738 24388 20750
rect 24444 20804 24500 20814
rect 24220 20066 24276 20076
rect 24444 20018 24500 20748
rect 24892 20802 24948 20814
rect 24892 20750 24894 20802
rect 24946 20750 24948 20802
rect 24892 20468 24948 20750
rect 25004 20804 25060 21420
rect 25004 20738 25060 20748
rect 24892 20402 24948 20412
rect 25004 20578 25060 20590
rect 25004 20526 25006 20578
rect 25058 20526 25060 20578
rect 25004 20356 25060 20526
rect 25004 20290 25060 20300
rect 25228 20188 25284 21534
rect 25564 20804 25620 20814
rect 25564 20468 25620 20748
rect 25564 20402 25620 20412
rect 24444 19966 24446 20018
rect 24498 19966 24500 20018
rect 24444 19954 24500 19966
rect 24668 20132 25284 20188
rect 25340 20244 25396 20254
rect 24668 20130 24724 20132
rect 24668 20078 24670 20130
rect 24722 20078 24724 20130
rect 23996 19842 24052 19852
rect 24668 19796 24724 20078
rect 24668 19730 24724 19740
rect 24522 19628 24786 19638
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24522 19562 24786 19572
rect 25116 18564 25172 20132
rect 25228 19906 25284 19918
rect 25228 19854 25230 19906
rect 25282 19854 25284 19906
rect 25228 19796 25284 19854
rect 25228 19348 25284 19740
rect 25228 19282 25284 19292
rect 25340 19346 25396 20188
rect 25340 19294 25342 19346
rect 25394 19294 25396 19346
rect 25340 19282 25396 19294
rect 25676 19236 25732 24668
rect 25900 24658 25956 24668
rect 26460 24722 26516 25228
rect 26572 24836 26628 24846
rect 26572 24742 26628 24780
rect 26460 24670 26462 24722
rect 26514 24670 26516 24722
rect 26460 24658 26516 24670
rect 27020 24722 27076 24734
rect 27020 24670 27022 24722
rect 27074 24670 27076 24722
rect 26348 24500 26404 24510
rect 25788 23154 25844 23166
rect 26348 23156 26404 24444
rect 26460 23380 26516 23390
rect 26460 23286 26516 23324
rect 25788 23102 25790 23154
rect 25842 23102 25844 23154
rect 25788 22260 25844 23102
rect 25788 21586 25844 22204
rect 25788 21534 25790 21586
rect 25842 21534 25844 21586
rect 25788 21522 25844 21534
rect 26236 23154 26404 23156
rect 26236 23102 26350 23154
rect 26402 23102 26404 23154
rect 26236 23100 26404 23102
rect 26236 20802 26292 23100
rect 26348 23090 26404 23100
rect 27020 23268 27076 24670
rect 27804 24724 27860 24734
rect 27804 24630 27860 24668
rect 28700 24722 28756 28700
rect 29184 28252 29448 28262
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29184 28186 29448 28196
rect 37212 27746 37268 27758
rect 37212 27694 37214 27746
rect 37266 27694 37268 27746
rect 37212 27636 37268 27694
rect 37212 27570 37268 27580
rect 33846 27468 34110 27478
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 33846 27402 34110 27412
rect 37324 27188 37380 31052
rect 37884 31042 37940 31052
rect 38220 30994 38276 31006
rect 38220 30942 38222 30994
rect 38274 30942 38276 30994
rect 37660 30884 37716 30894
rect 38220 30884 38276 30942
rect 37660 30882 38276 30884
rect 37660 30830 37662 30882
rect 37714 30830 38276 30882
rect 37660 30828 38276 30830
rect 37660 30818 37716 30828
rect 38220 30324 38276 30828
rect 38220 30258 38276 30268
rect 37660 30100 37716 30110
rect 37660 30006 37716 30044
rect 38220 30100 38276 30110
rect 37884 29988 37940 29998
rect 37884 29894 37940 29932
rect 38220 29652 38276 30044
rect 38892 29988 38948 29998
rect 38508 29820 38772 29830
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38508 29754 38772 29764
rect 38220 29586 38276 29596
rect 37884 29540 37940 29550
rect 37212 27132 37380 27188
rect 37436 29538 37940 29540
rect 37436 29486 37886 29538
rect 37938 29486 37940 29538
rect 37436 29484 37940 29486
rect 37100 27076 37156 27086
rect 36988 26850 37044 26862
rect 36988 26798 36990 26850
rect 37042 26798 37044 26850
rect 29184 26684 29448 26694
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29184 26618 29448 26628
rect 33846 25900 34110 25910
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 33846 25834 34110 25844
rect 29184 25116 29448 25126
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29184 25050 29448 25060
rect 28700 24670 28702 24722
rect 28754 24670 28756 24722
rect 28700 24658 28756 24670
rect 36988 24724 37044 26798
rect 36988 24658 37044 24668
rect 33846 24332 34110 24342
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 33846 24266 34110 24276
rect 29184 23548 29448 23558
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29184 23482 29448 23492
rect 27020 23154 27076 23212
rect 27020 23102 27022 23154
rect 27074 23102 27076 23154
rect 27020 23090 27076 23102
rect 27692 23154 27748 23166
rect 27692 23102 27694 23154
rect 27746 23102 27748 23154
rect 27692 22932 27748 23102
rect 28476 23156 28532 23166
rect 28476 23062 28532 23100
rect 28812 23156 28868 23166
rect 27692 22866 27748 22876
rect 28812 22932 28868 23100
rect 28252 21028 28308 21038
rect 28252 20914 28308 20972
rect 28252 20862 28254 20914
rect 28306 20862 28308 20914
rect 28252 20850 28308 20862
rect 26236 20750 26238 20802
rect 26290 20750 26292 20802
rect 26236 20738 26292 20750
rect 27132 20804 27188 20814
rect 27132 20710 27188 20748
rect 27804 20692 27860 20702
rect 27804 20598 27860 20636
rect 25788 20468 25844 20478
rect 25788 20242 25844 20412
rect 25788 20190 25790 20242
rect 25842 20190 25844 20242
rect 25788 20178 25844 20190
rect 26908 20020 26964 20030
rect 26908 19926 26964 19964
rect 27468 20018 27524 20030
rect 27468 19966 27470 20018
rect 27522 19966 27524 20018
rect 26236 19906 26292 19918
rect 26236 19854 26238 19906
rect 26290 19854 26292 19906
rect 26236 19796 26292 19854
rect 26572 19908 26628 19918
rect 26572 19814 26628 19852
rect 26236 19730 26292 19740
rect 25788 19236 25844 19246
rect 25676 19234 25844 19236
rect 25676 19182 25790 19234
rect 25842 19182 25844 19234
rect 25676 19180 25844 19182
rect 25116 18508 25284 18564
rect 25228 18450 25284 18508
rect 25228 18398 25230 18450
rect 25282 18398 25284 18450
rect 25228 18386 25284 18398
rect 25788 18338 25844 19180
rect 26236 19236 26292 19246
rect 26236 19142 26292 19180
rect 26908 19234 26964 19246
rect 26908 19182 26910 19234
rect 26962 19182 26964 19234
rect 26348 19124 26404 19134
rect 26348 19030 26404 19068
rect 25788 18286 25790 18338
rect 25842 18286 25844 18338
rect 24522 18060 24786 18070
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24522 17994 24786 18004
rect 25788 17666 25844 18286
rect 25788 17614 25790 17666
rect 25842 17614 25844 17666
rect 25340 17556 25396 17566
rect 25340 17462 25396 17500
rect 23884 17350 23940 17388
rect 24220 17444 24276 17454
rect 25788 17444 25844 17614
rect 26236 17666 26292 17678
rect 26236 17614 26238 17666
rect 26290 17614 26292 17666
rect 25788 17388 26068 17444
rect 21868 16830 21870 16882
rect 21922 16830 21924 16882
rect 21420 16772 21476 16782
rect 21308 16770 21476 16772
rect 21308 16718 21422 16770
rect 21474 16718 21476 16770
rect 21308 16716 21476 16718
rect 21196 15428 21252 15438
rect 20636 15314 20692 15326
rect 20636 15262 20638 15314
rect 20690 15262 20692 15314
rect 20636 14756 20692 15262
rect 21196 15314 21252 15372
rect 21196 15262 21198 15314
rect 21250 15262 21252 15314
rect 21196 15250 21252 15262
rect 20972 15092 21028 15102
rect 21308 15092 21364 16716
rect 21420 16706 21476 16716
rect 21644 16324 21700 16334
rect 21644 15538 21700 16268
rect 21644 15486 21646 15538
rect 21698 15486 21700 15538
rect 21644 15474 21700 15486
rect 20636 14690 20692 14700
rect 20748 15090 21028 15092
rect 20748 15038 20974 15090
rect 21026 15038 21028 15090
rect 20748 15036 21028 15038
rect 20636 14532 20692 14542
rect 20468 14476 20580 14532
rect 20412 14466 20468 14476
rect 20412 14308 20468 14318
rect 20412 14214 20468 14252
rect 20524 13748 20580 14476
rect 20636 14438 20692 14476
rect 20748 14308 20804 15036
rect 20972 15026 21028 15036
rect 21196 15036 21364 15092
rect 21420 15314 21476 15326
rect 21420 15262 21422 15314
rect 21474 15262 21476 15314
rect 21196 14532 21252 15036
rect 20524 13682 20580 13692
rect 20636 14252 20804 14308
rect 20860 14476 21252 14532
rect 21308 14868 21364 14878
rect 21308 14530 21364 14812
rect 21420 14644 21476 15262
rect 21532 15316 21588 15326
rect 21532 15222 21588 15260
rect 21420 14578 21476 14588
rect 21308 14478 21310 14530
rect 21362 14478 21364 14530
rect 20356 13468 20580 13524
rect 20300 13458 20356 13468
rect 20188 13244 20356 13300
rect 20076 13010 20132 13020
rect 19740 12910 19742 12962
rect 19794 12910 19796 12962
rect 18956 12740 19012 12750
rect 18956 12646 19012 12684
rect 18956 12404 19012 12414
rect 18956 12310 19012 12348
rect 18844 12124 19124 12180
rect 18732 11778 18788 11788
rect 18620 4610 18676 4620
rect 18844 4226 18900 4238
rect 18844 4174 18846 4226
rect 18898 4174 18900 4226
rect 18620 3556 18676 3566
rect 18620 3462 18676 3500
rect 18396 3390 18398 3442
rect 18450 3390 18452 3442
rect 18396 3378 18452 3390
rect 18844 2548 18900 4174
rect 19068 3442 19124 12124
rect 19740 12178 19796 12910
rect 20076 12850 20132 12862
rect 20076 12798 20078 12850
rect 20130 12798 20132 12850
rect 20076 12740 20132 12798
rect 20076 12684 20244 12740
rect 19860 12572 20124 12582
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 19860 12506 20124 12516
rect 20188 12404 20244 12684
rect 20076 12348 20244 12404
rect 19740 12126 19742 12178
rect 19794 12126 19796 12178
rect 19740 12114 19796 12126
rect 19852 12290 19908 12302
rect 19852 12238 19854 12290
rect 19906 12238 19908 12290
rect 19292 11954 19348 11966
rect 19292 11902 19294 11954
rect 19346 11902 19348 11954
rect 19292 10164 19348 11902
rect 19852 11172 19908 12238
rect 19292 10098 19348 10108
rect 19740 11116 19908 11172
rect 20076 11172 20132 12348
rect 19516 3668 19572 3678
rect 19068 3390 19070 3442
rect 19122 3390 19124 3442
rect 19068 3378 19124 3390
rect 19292 3554 19348 3566
rect 19292 3502 19294 3554
rect 19346 3502 19348 3554
rect 19292 2548 19348 3502
rect 18844 2492 19348 2548
rect 18844 800 18900 2492
rect 19516 800 19572 3612
rect 19740 3444 19796 11116
rect 20076 11106 20132 11116
rect 19860 11004 20124 11014
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 19860 10938 20124 10948
rect 19860 9436 20124 9446
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 19860 9370 20124 9380
rect 19860 7868 20124 7878
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 19860 7802 20124 7812
rect 19860 6300 20124 6310
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 19860 6234 20124 6244
rect 19860 4732 20124 4742
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 19860 4666 20124 4676
rect 19964 4226 20020 4238
rect 19964 4174 19966 4226
rect 20018 4174 20020 4226
rect 19964 3556 20020 4174
rect 20076 3556 20132 3566
rect 19964 3554 20132 3556
rect 19964 3502 20078 3554
rect 20130 3502 20132 3554
rect 19964 3500 20132 3502
rect 19852 3444 19908 3454
rect 19740 3442 19908 3444
rect 19740 3390 19854 3442
rect 19906 3390 19908 3442
rect 19740 3388 19908 3390
rect 19852 3378 19908 3388
rect 20076 3388 20132 3500
rect 20300 3444 20356 13244
rect 20524 12178 20580 13468
rect 20524 12126 20526 12178
rect 20578 12126 20580 12178
rect 20524 12114 20580 12126
rect 20636 4564 20692 14252
rect 20748 12740 20804 12750
rect 20748 12178 20804 12684
rect 20748 12126 20750 12178
rect 20802 12126 20804 12178
rect 20748 12114 20804 12126
rect 20636 4498 20692 4508
rect 20860 4564 20916 14476
rect 21308 14466 21364 14478
rect 21532 14532 21588 14542
rect 21588 14476 21812 14532
rect 21532 14466 21588 14476
rect 21420 14420 21476 14430
rect 21420 14326 21476 14364
rect 21196 14308 21252 14318
rect 20972 13748 21028 13758
rect 20972 12740 21028 13692
rect 20972 12402 21028 12684
rect 20972 12350 20974 12402
rect 21026 12350 21028 12402
rect 20972 12338 21028 12350
rect 21084 13636 21140 13646
rect 21084 12402 21140 13580
rect 21084 12350 21086 12402
rect 21138 12350 21140 12402
rect 21084 12338 21140 12350
rect 21196 12402 21252 14252
rect 21420 13634 21476 13646
rect 21420 13582 21422 13634
rect 21474 13582 21476 13634
rect 21308 13524 21364 13534
rect 21308 13186 21364 13468
rect 21308 13134 21310 13186
rect 21362 13134 21364 13186
rect 21308 13122 21364 13134
rect 21196 12350 21198 12402
rect 21250 12350 21252 12402
rect 21196 12338 21252 12350
rect 20860 4498 20916 4508
rect 21084 11172 21140 11182
rect 21084 4562 21140 11116
rect 21420 4900 21476 13582
rect 21644 13076 21700 13086
rect 21756 13076 21812 14476
rect 21868 13746 21924 16830
rect 21980 16772 22036 16782
rect 22204 16772 22260 17052
rect 22428 16996 22484 17006
rect 22428 16902 22484 16940
rect 22036 16716 22260 16772
rect 22316 16882 22372 16894
rect 22316 16830 22318 16882
rect 22370 16830 22372 16882
rect 22316 16772 22372 16830
rect 21980 16706 22036 16716
rect 22092 13860 22148 16716
rect 22316 16706 22372 16716
rect 22988 15148 23044 17052
rect 23660 17108 23716 17118
rect 23100 16884 23156 16894
rect 23100 16790 23156 16828
rect 23660 16882 23716 17052
rect 23660 16830 23662 16882
rect 23714 16830 23716 16882
rect 23660 16818 23716 16830
rect 24220 16884 24276 17388
rect 24220 16818 24276 16828
rect 24556 16884 24612 16894
rect 26012 16884 26068 17388
rect 26236 17108 26292 17614
rect 26348 17668 26404 17678
rect 26348 17554 26404 17612
rect 26348 17502 26350 17554
rect 26402 17502 26404 17554
rect 26348 17490 26404 17502
rect 26908 17666 26964 19182
rect 27468 19012 27524 19966
rect 28812 20018 28868 22876
rect 33846 22764 34110 22774
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 33846 22698 34110 22708
rect 36540 22260 36596 22270
rect 36540 22166 36596 22204
rect 29184 21980 29448 21990
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29184 21914 29448 21924
rect 33846 21196 34110 21206
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 33846 21130 34110 21140
rect 37100 21028 37156 27020
rect 37212 26404 37268 27132
rect 37324 26964 37380 26974
rect 37324 26870 37380 26908
rect 37212 26348 37380 26404
rect 37212 26180 37268 26190
rect 37212 26086 37268 26124
rect 37324 23268 37380 26348
rect 37436 24612 37492 29484
rect 37884 29474 37940 29484
rect 38220 29426 38276 29438
rect 38220 29374 38222 29426
rect 38274 29374 38276 29426
rect 37660 29316 37716 29326
rect 38220 29316 38276 29374
rect 37660 29314 38276 29316
rect 37660 29262 37662 29314
rect 37714 29262 38276 29314
rect 37660 29260 38276 29262
rect 37660 29250 37716 29260
rect 38220 28980 38276 29260
rect 38220 28914 38276 28924
rect 37884 28756 37940 28766
rect 37660 28644 37716 28654
rect 37660 28550 37716 28588
rect 37884 28530 37940 28700
rect 38108 28644 38164 28654
rect 38108 28550 38164 28588
rect 37884 28478 37886 28530
rect 37938 28478 37940 28530
rect 37884 28466 37940 28478
rect 38508 28252 38772 28262
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38508 28186 38772 28196
rect 37884 27972 37940 27982
rect 37884 27970 38164 27972
rect 37884 27918 37886 27970
rect 37938 27918 38164 27970
rect 37884 27916 38164 27918
rect 37884 27906 37940 27916
rect 37660 27748 37716 27758
rect 37660 27746 37940 27748
rect 37660 27694 37662 27746
rect 37714 27694 37940 27746
rect 37660 27692 37940 27694
rect 37660 27682 37716 27692
rect 37660 27076 37716 27086
rect 37884 27076 37940 27692
rect 38108 27300 38164 27916
rect 38220 27858 38276 27870
rect 38220 27806 38222 27858
rect 38274 27806 38276 27858
rect 38220 27636 38276 27806
rect 38220 27570 38276 27580
rect 38108 27244 38388 27300
rect 38108 27076 38164 27086
rect 37884 27074 38164 27076
rect 37884 27022 38110 27074
rect 38162 27022 38164 27074
rect 37884 27020 38164 27022
rect 37660 26982 37716 27020
rect 37772 26964 37828 26974
rect 37660 26516 37716 26526
rect 37772 26516 37828 26908
rect 37660 26514 37828 26516
rect 37660 26462 37662 26514
rect 37714 26462 37828 26514
rect 37660 26460 37828 26462
rect 37660 26450 37716 26460
rect 37884 26404 37940 26414
rect 37884 26402 38052 26404
rect 37884 26350 37886 26402
rect 37938 26350 38052 26402
rect 37884 26348 38052 26350
rect 37884 26338 37940 26348
rect 37660 25396 37716 25406
rect 37660 25302 37716 25340
rect 37884 25284 37940 25294
rect 37884 25190 37940 25228
rect 37884 24836 37940 24846
rect 37436 24546 37492 24556
rect 37548 24834 37940 24836
rect 37548 24782 37886 24834
rect 37938 24782 37940 24834
rect 37548 24780 37940 24782
rect 37324 23202 37380 23212
rect 37548 23156 37604 24780
rect 37884 24770 37940 24780
rect 37996 24836 38052 26348
rect 38108 26292 38164 27020
rect 38108 26226 38164 26236
rect 38220 26290 38276 26302
rect 38220 26238 38222 26290
rect 38274 26238 38276 26290
rect 38220 26180 38276 26238
rect 38220 25620 38276 26124
rect 38220 25554 38276 25564
rect 38220 25396 38276 25406
rect 38220 24948 38276 25340
rect 38220 24882 38276 24892
rect 37996 24770 38052 24780
rect 38220 24722 38276 24734
rect 38220 24670 38222 24722
rect 38274 24670 38276 24722
rect 37660 24612 37716 24622
rect 38220 24612 38276 24670
rect 37660 24610 38276 24612
rect 37660 24558 37662 24610
rect 37714 24558 38276 24610
rect 37660 24556 38276 24558
rect 37660 24546 37716 24556
rect 38220 24276 38276 24556
rect 38220 24210 38276 24220
rect 38220 23826 38276 23838
rect 38220 23774 38222 23826
rect 38274 23774 38276 23826
rect 37660 23716 37716 23726
rect 37660 23622 37716 23660
rect 37884 23716 37940 23726
rect 38220 23716 38276 23774
rect 37884 23714 38052 23716
rect 37884 23662 37886 23714
rect 37938 23662 38052 23714
rect 37884 23660 38052 23662
rect 37884 23650 37940 23660
rect 37884 23268 37940 23278
rect 37548 23090 37604 23100
rect 37772 23266 37940 23268
rect 37772 23214 37886 23266
rect 37938 23214 37940 23266
rect 37772 23212 37940 23214
rect 37660 23042 37716 23054
rect 37660 22990 37662 23042
rect 37714 22990 37716 23042
rect 37660 22932 37716 22990
rect 37660 22866 37716 22876
rect 37772 22484 37828 23212
rect 37884 23202 37940 23212
rect 37436 22428 37828 22484
rect 37212 22148 37268 22158
rect 37212 22146 37380 22148
rect 37212 22094 37214 22146
rect 37266 22094 37380 22146
rect 37212 22092 37380 22094
rect 37212 22082 37268 22092
rect 37212 21476 37268 21486
rect 37212 21382 37268 21420
rect 37100 20962 37156 20972
rect 29932 20468 29988 20478
rect 29184 20412 29448 20422
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29184 20346 29448 20356
rect 29932 20244 29988 20412
rect 29932 20178 29988 20188
rect 36988 20132 37044 20142
rect 28812 19966 28814 20018
rect 28866 19966 28868 20018
rect 28812 19954 28868 19966
rect 29932 20020 29988 20030
rect 29932 19926 29988 19964
rect 27692 19906 27748 19918
rect 27692 19854 27694 19906
rect 27746 19854 27748 19906
rect 27692 19460 27748 19854
rect 28476 19796 28532 19806
rect 28476 19702 28532 19740
rect 33846 19628 34110 19638
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 33846 19562 34110 19572
rect 27692 19394 27748 19404
rect 27580 19236 27636 19246
rect 27580 19142 27636 19180
rect 28476 19234 28532 19246
rect 28476 19182 28478 19234
rect 28530 19182 28532 19234
rect 27468 18946 27524 18956
rect 28476 19012 28532 19182
rect 36988 19236 37044 20076
rect 37324 20020 37380 22092
rect 37436 20356 37492 22428
rect 37548 22258 37604 22270
rect 37548 22206 37550 22258
rect 37602 22206 37604 22258
rect 37548 21588 37604 22206
rect 37884 22148 37940 22158
rect 37548 21494 37604 21532
rect 37660 22146 37940 22148
rect 37660 22094 37886 22146
rect 37938 22094 37940 22146
rect 37660 22092 37940 22094
rect 37660 21140 37716 22092
rect 37884 22082 37940 22092
rect 37436 20290 37492 20300
rect 37548 21084 37716 21140
rect 37884 21698 37940 21710
rect 37884 21646 37886 21698
rect 37938 21646 37940 21698
rect 37324 19954 37380 19964
rect 37548 19908 37604 21084
rect 37884 20804 37940 21646
rect 37996 20916 38052 23660
rect 38220 23650 38276 23660
rect 38220 23154 38276 23166
rect 38220 23102 38222 23154
rect 38274 23102 38276 23154
rect 38220 22932 38276 23102
rect 38332 23044 38388 27244
rect 38508 26684 38772 26694
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38508 26618 38772 26628
rect 38508 25116 38772 25126
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38508 25050 38772 25060
rect 38508 23548 38772 23558
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38508 23482 38772 23492
rect 38332 22978 38388 22988
rect 38220 22866 38276 22876
rect 38220 22260 38276 22270
rect 38220 22166 38276 22204
rect 38508 21980 38772 21990
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38508 21914 38772 21924
rect 37996 20850 38052 20860
rect 38220 21586 38276 21598
rect 38220 21534 38222 21586
rect 38274 21534 38276 21586
rect 38220 21476 38276 21534
rect 38220 20916 38276 21420
rect 38220 20850 38276 20860
rect 37884 20738 37940 20748
rect 38220 20690 38276 20702
rect 38220 20638 38222 20690
rect 38274 20638 38276 20690
rect 37660 20578 37716 20590
rect 37660 20526 37662 20578
rect 37714 20526 37716 20578
rect 37660 20244 37716 20526
rect 37884 20580 37940 20590
rect 37884 20486 37940 20524
rect 37660 20178 37716 20188
rect 38220 20244 38276 20638
rect 38892 20692 38948 29932
rect 38892 20626 38948 20636
rect 38508 20412 38772 20422
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38508 20346 38772 20356
rect 38220 20178 38276 20188
rect 37884 20132 37940 20142
rect 37884 20038 37940 20076
rect 38220 20018 38276 20030
rect 38220 19966 38222 20018
rect 38274 19966 38276 20018
rect 37548 19842 37604 19852
rect 37660 19908 37716 19918
rect 38220 19908 38276 19966
rect 37660 19906 38276 19908
rect 37660 19854 37662 19906
rect 37714 19854 38276 19906
rect 37660 19852 38276 19854
rect 37660 19842 37716 19852
rect 38220 19572 38276 19852
rect 38220 19506 38276 19516
rect 36988 19170 37044 19180
rect 37884 19348 37940 19358
rect 37884 19122 37940 19292
rect 37884 19070 37886 19122
rect 37938 19070 37940 19122
rect 37884 19058 37940 19070
rect 38220 19122 38276 19134
rect 38220 19070 38222 19122
rect 38274 19070 38276 19122
rect 28476 18946 28532 18956
rect 37660 19012 37716 19022
rect 37660 18918 37716 18956
rect 38220 19012 38276 19070
rect 38220 18946 38276 18956
rect 37772 18900 37828 18910
rect 29184 18844 29448 18854
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29184 18778 29448 18788
rect 37772 18676 37828 18844
rect 38508 18844 38772 18854
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38508 18778 38772 18788
rect 37884 18676 37940 18686
rect 37772 18674 37940 18676
rect 37772 18622 37886 18674
rect 37938 18622 37940 18674
rect 37772 18620 37940 18622
rect 37884 18610 37940 18620
rect 38220 18450 38276 18462
rect 38220 18398 38222 18450
rect 38274 18398 38276 18450
rect 37660 18338 37716 18350
rect 37660 18286 37662 18338
rect 37714 18286 37716 18338
rect 37660 18228 37716 18286
rect 37660 18162 37716 18172
rect 37884 18340 37940 18350
rect 33846 18060 34110 18070
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 33846 17994 34110 18004
rect 26908 17614 26910 17666
rect 26962 17614 26964 17666
rect 26908 17444 26964 17614
rect 26908 17378 26964 17388
rect 27356 17666 27412 17678
rect 27356 17614 27358 17666
rect 27410 17614 27412 17666
rect 26908 17220 26964 17230
rect 26236 17052 26404 17108
rect 26236 16884 26292 16894
rect 24556 16882 24948 16884
rect 24556 16830 24558 16882
rect 24610 16830 24948 16882
rect 24556 16828 24948 16830
rect 26012 16882 26292 16884
rect 26012 16830 26238 16882
rect 26290 16830 26292 16882
rect 26012 16828 26292 16830
rect 24556 16818 24612 16828
rect 24522 16492 24786 16502
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24522 16426 24786 16436
rect 22988 15092 23268 15148
rect 22204 14530 22260 14542
rect 22204 14478 22206 14530
rect 22258 14478 22260 14530
rect 22204 13972 22260 14478
rect 23212 14530 23268 15092
rect 24522 14924 24786 14934
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24522 14858 24786 14868
rect 23212 14478 23214 14530
rect 23266 14478 23268 14530
rect 22764 14418 22820 14430
rect 22764 14366 22766 14418
rect 22818 14366 22820 14418
rect 22316 14308 22372 14318
rect 22316 14306 22708 14308
rect 22316 14254 22318 14306
rect 22370 14254 22708 14306
rect 22316 14252 22708 14254
rect 22316 14242 22372 14252
rect 22204 13906 22260 13916
rect 22428 13860 22484 13870
rect 22092 13794 22148 13804
rect 22316 13858 22484 13860
rect 22316 13806 22430 13858
rect 22482 13806 22484 13858
rect 22316 13804 22484 13806
rect 21868 13694 21870 13746
rect 21922 13694 21924 13746
rect 21868 13682 21924 13694
rect 22204 13748 22260 13758
rect 22204 13654 22260 13692
rect 22316 13300 22372 13804
rect 22428 13794 22484 13804
rect 21980 13244 22372 13300
rect 21868 13076 21924 13086
rect 21756 13074 21924 13076
rect 21756 13022 21870 13074
rect 21922 13022 21924 13074
rect 21756 13020 21924 13022
rect 21532 12962 21588 12974
rect 21532 12910 21534 12962
rect 21586 12910 21588 12962
rect 21532 12404 21588 12910
rect 21532 12338 21588 12348
rect 21420 4834 21476 4844
rect 21084 4510 21086 4562
rect 21138 4510 21140 4562
rect 21084 4498 21140 4510
rect 21644 4564 21700 13020
rect 21868 13010 21924 13020
rect 21980 12962 22036 13244
rect 21980 12910 21982 12962
rect 22034 12910 22036 12962
rect 21980 12898 22036 12910
rect 21756 12740 21812 12750
rect 21756 12646 21812 12684
rect 22652 8932 22708 14252
rect 22764 13076 22820 14366
rect 22876 13860 22932 13870
rect 22876 13766 22932 13804
rect 22764 13010 22820 13020
rect 23212 12962 23268 14478
rect 23660 14530 23716 14542
rect 23660 14478 23662 14530
rect 23714 14478 23716 14530
rect 23212 12910 23214 12962
rect 23266 12910 23268 12962
rect 23212 12898 23268 12910
rect 23548 13746 23604 13758
rect 23548 13694 23550 13746
rect 23602 13694 23604 13746
rect 22764 12852 22820 12862
rect 22764 12850 23044 12852
rect 22764 12798 22766 12850
rect 22818 12798 23044 12850
rect 22764 12796 23044 12798
rect 22764 12786 22820 12796
rect 22652 8876 22932 8932
rect 22204 4900 22260 4910
rect 22204 4898 22708 4900
rect 22204 4846 22206 4898
rect 22258 4846 22708 4898
rect 22204 4844 22708 4846
rect 21756 4564 21812 4574
rect 21644 4562 21812 4564
rect 21644 4510 21758 4562
rect 21810 4510 21812 4562
rect 21644 4508 21812 4510
rect 21756 4498 21812 4508
rect 20860 4340 20916 4350
rect 20860 4246 20916 4284
rect 21308 4338 21364 4350
rect 21308 4286 21310 4338
rect 21362 4286 21364 4338
rect 20076 3332 20244 3388
rect 20300 3378 20356 3388
rect 20412 4226 20468 4238
rect 20412 4174 20414 4226
rect 20466 4174 20468 4226
rect 19860 3164 20124 3174
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 19860 3098 20124 3108
rect 20188 800 20244 3332
rect 20412 2884 20468 4174
rect 20972 3668 21028 3678
rect 20972 3574 21028 3612
rect 21308 2884 21364 4286
rect 20412 2828 21364 2884
rect 21532 4340 21588 4350
rect 20860 800 20916 2828
rect 21532 800 21588 4284
rect 21980 4340 22036 4350
rect 21980 4246 22036 4284
rect 22204 800 22260 4844
rect 22428 4564 22484 4574
rect 22428 4470 22484 4508
rect 22652 4338 22708 4844
rect 22652 4286 22654 4338
rect 22706 4286 22708 4338
rect 22652 4274 22708 4286
rect 22876 3554 22932 8876
rect 22988 5012 23044 12796
rect 22988 4946 23044 4956
rect 22876 3502 22878 3554
rect 22930 3502 22932 3554
rect 22876 3490 22932 3502
rect 23436 4226 23492 4238
rect 23436 4174 23438 4226
rect 23490 4174 23492 4226
rect 22988 3444 23044 3454
rect 22876 3332 23044 3388
rect 23436 3444 23492 4174
rect 23548 3780 23604 13694
rect 23660 13188 23716 14478
rect 24220 14418 24276 14430
rect 24220 14366 24222 14418
rect 24274 14366 24276 14418
rect 23772 14308 23828 14318
rect 23772 14214 23828 14252
rect 24220 13860 24276 14366
rect 24892 13972 24948 16828
rect 26236 16818 26292 16828
rect 25900 16772 25956 16782
rect 25900 16770 26068 16772
rect 25900 16718 25902 16770
rect 25954 16718 26068 16770
rect 25900 16716 26068 16718
rect 25900 16706 25956 16716
rect 25004 14532 25060 14542
rect 25004 14438 25060 14476
rect 25900 14530 25956 14542
rect 25900 14478 25902 14530
rect 25954 14478 25956 14530
rect 24892 13906 24948 13916
rect 23660 13132 23828 13188
rect 23660 12962 23716 12974
rect 23660 12910 23662 12962
rect 23714 12910 23716 12962
rect 23660 10388 23716 12910
rect 23772 12964 23828 13132
rect 23772 12898 23828 12908
rect 24220 12962 24276 13804
rect 24556 13748 24612 13758
rect 25452 13748 25508 13758
rect 24556 13746 24948 13748
rect 24556 13694 24558 13746
rect 24610 13694 24948 13746
rect 24556 13692 24948 13694
rect 24556 13682 24612 13692
rect 24522 13356 24786 13366
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24522 13290 24786 13300
rect 24220 12910 24222 12962
rect 24274 12910 24276 12962
rect 24220 12898 24276 12910
rect 24332 13076 24388 13086
rect 23772 12740 23828 12750
rect 23772 12646 23828 12684
rect 23660 10322 23716 10332
rect 23548 3714 23604 3724
rect 23660 4900 23716 4910
rect 23436 3378 23492 3388
rect 23660 3442 23716 4844
rect 24332 4452 24388 13020
rect 24522 11788 24786 11798
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24522 11722 24786 11732
rect 24522 10220 24786 10230
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24522 10154 24786 10164
rect 24522 8652 24786 8662
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24522 8586 24786 8596
rect 24522 7084 24786 7094
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24522 7018 24786 7028
rect 24522 5516 24786 5526
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24522 5450 24786 5460
rect 24892 4564 24948 13692
rect 25452 13654 25508 13692
rect 25900 13188 25956 14478
rect 25900 13122 25956 13132
rect 24892 4498 24948 4508
rect 25004 12962 25060 12974
rect 25004 12910 25006 12962
rect 25058 12910 25060 12962
rect 24220 4396 24388 4452
rect 25004 4452 25060 12910
rect 25900 12962 25956 12974
rect 25900 12910 25902 12962
rect 25954 12910 25956 12962
rect 25788 10388 25844 10398
rect 23660 3390 23662 3442
rect 23714 3390 23716 3442
rect 23660 3378 23716 3390
rect 23884 3554 23940 3566
rect 23884 3502 23886 3554
rect 23938 3502 23940 3554
rect 23884 3444 23940 3502
rect 24220 3444 24276 4396
rect 25004 4386 25060 4396
rect 25228 5012 25284 5022
rect 24332 4226 24388 4238
rect 24332 4174 24334 4226
rect 24386 4174 24388 4226
rect 24332 3668 24388 4174
rect 24522 3948 24786 3958
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24522 3882 24786 3892
rect 24332 3612 24836 3668
rect 24780 3554 24836 3612
rect 24780 3502 24782 3554
rect 24834 3502 24836 3554
rect 24556 3444 24612 3454
rect 24220 3442 24612 3444
rect 24220 3390 24558 3442
rect 24610 3390 24612 3442
rect 24220 3388 24612 3390
rect 23884 3378 23940 3388
rect 24556 3378 24612 3388
rect 22876 800 22932 3332
rect 24780 2548 24836 3502
rect 23548 2492 24836 2548
rect 24892 3556 24948 3566
rect 23548 800 23604 2492
rect 24892 2324 24948 3500
rect 24220 2268 24948 2324
rect 25004 3444 25060 3454
rect 24220 800 24276 2268
rect 25004 2212 25060 3388
rect 25228 3442 25284 4956
rect 25452 4226 25508 4238
rect 25452 4174 25454 4226
rect 25506 4174 25508 4226
rect 25452 3556 25508 4174
rect 25452 3462 25508 3500
rect 25564 4114 25620 4126
rect 25564 4062 25566 4114
rect 25618 4062 25620 4114
rect 25228 3390 25230 3442
rect 25282 3390 25284 3442
rect 25228 3378 25284 3390
rect 24892 2156 25060 2212
rect 24892 800 24948 2156
rect 25564 800 25620 4062
rect 25788 3444 25844 10332
rect 25900 5012 25956 12910
rect 26012 12292 26068 16716
rect 26348 15428 26404 17052
rect 26908 17106 26964 17164
rect 26908 17054 26910 17106
rect 26962 17054 26964 17106
rect 26908 17042 26964 17054
rect 26796 16882 26852 16894
rect 26796 16830 26798 16882
rect 26850 16830 26852 16882
rect 26796 15876 26852 16830
rect 26796 15810 26852 15820
rect 26348 15362 26404 15372
rect 26012 12226 26068 12236
rect 26572 12964 26628 12974
rect 25900 4946 25956 4956
rect 25900 4226 25956 4238
rect 25900 4174 25902 4226
rect 25954 4174 25956 4226
rect 25900 3780 25956 4174
rect 26348 4226 26404 4238
rect 26348 4174 26350 4226
rect 26402 4174 26404 4226
rect 26348 4114 26404 4174
rect 26348 4062 26350 4114
rect 26402 4062 26404 4114
rect 26348 4050 26404 4062
rect 25900 3724 26292 3780
rect 26124 3556 26180 3566
rect 25900 3444 25956 3454
rect 25788 3442 25956 3444
rect 25788 3390 25902 3442
rect 25954 3390 25956 3442
rect 25788 3388 25956 3390
rect 25900 3378 25956 3388
rect 26124 3388 26180 3500
rect 26236 3556 26292 3724
rect 26236 3554 26404 3556
rect 26236 3502 26238 3554
rect 26290 3502 26404 3554
rect 26236 3500 26404 3502
rect 26236 3490 26292 3500
rect 26348 3444 26404 3500
rect 26124 3332 26292 3388
rect 26348 3378 26404 3388
rect 26572 3442 26628 12908
rect 27356 12852 27412 17614
rect 28476 17666 28532 17678
rect 28476 17614 28478 17666
rect 28530 17614 28532 17666
rect 27468 17444 27524 17454
rect 27468 16882 27524 17388
rect 27468 16830 27470 16882
rect 27522 16830 27524 16882
rect 27468 16818 27524 16830
rect 28140 16882 28196 16894
rect 28140 16830 28142 16882
rect 28194 16830 28196 16882
rect 28140 12964 28196 16830
rect 28140 12898 28196 12908
rect 28252 13188 28308 13198
rect 27356 12786 27412 12796
rect 27132 4564 27188 4574
rect 27132 4470 27188 4508
rect 27356 4338 27412 4350
rect 27356 4286 27358 4338
rect 27410 4286 27412 4338
rect 26908 4228 26964 4238
rect 27356 4228 27412 4286
rect 26908 4226 27412 4228
rect 26908 4174 26910 4226
rect 26962 4174 27412 4226
rect 26908 4172 27412 4174
rect 27916 4226 27972 4238
rect 27916 4174 27918 4226
rect 27970 4174 27972 4226
rect 26908 4162 26964 4172
rect 26796 4114 26852 4126
rect 26796 4062 26798 4114
rect 26850 4062 26852 4114
rect 26796 3554 26852 4062
rect 26796 3502 26798 3554
rect 26850 3502 26852 3554
rect 26796 3490 26852 3502
rect 26572 3390 26574 3442
rect 26626 3390 26628 3442
rect 26572 3378 26628 3390
rect 26236 800 26292 3332
rect 27020 2996 27076 4172
rect 27244 3780 27300 3790
rect 27244 3442 27300 3724
rect 27468 3556 27524 3566
rect 27468 3462 27524 3500
rect 27916 3556 27972 4174
rect 27916 3490 27972 3500
rect 28140 3556 28196 3566
rect 27244 3390 27246 3442
rect 27298 3390 27300 3442
rect 27244 3378 27300 3390
rect 27692 3444 27748 3454
rect 27692 3108 27748 3388
rect 26908 2940 27076 2996
rect 27580 3052 27748 3108
rect 28140 3108 28196 3500
rect 28252 3444 28308 13132
rect 28476 10724 28532 17614
rect 29260 17556 29316 17566
rect 29260 17462 29316 17500
rect 29596 17556 29652 17566
rect 29184 17276 29448 17286
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29184 17210 29448 17220
rect 29596 16996 29652 17500
rect 36540 17556 36596 17566
rect 36540 17462 36596 17500
rect 37548 17554 37604 17566
rect 37548 17502 37550 17554
rect 37602 17502 37604 17554
rect 37212 17442 37268 17454
rect 37212 17390 37214 17442
rect 37266 17390 37268 17442
rect 37212 17108 37268 17390
rect 37212 17042 37268 17052
rect 29596 16930 29652 16940
rect 37324 16996 37380 17006
rect 37548 16996 37604 17502
rect 37884 17554 37940 18284
rect 38220 18228 38276 18398
rect 38220 18162 38276 18172
rect 37884 17502 37886 17554
rect 37938 17502 37940 17554
rect 37884 17490 37940 17502
rect 38220 17556 38276 17566
rect 38220 17462 38276 17500
rect 38508 17276 38772 17286
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38508 17210 38772 17220
rect 37380 16940 37492 16996
rect 37324 16930 37380 16940
rect 29036 16882 29092 16894
rect 29036 16830 29038 16882
rect 29090 16830 29092 16882
rect 29036 14308 29092 16830
rect 37212 16884 37268 16894
rect 37212 16790 37268 16828
rect 33846 16492 34110 16502
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 33846 16426 34110 16436
rect 29184 15708 29448 15718
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29184 15642 29448 15652
rect 33846 14924 34110 14934
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 33846 14858 34110 14868
rect 29036 14242 29092 14252
rect 31052 14532 31108 14542
rect 29184 14140 29448 14150
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29184 14074 29448 14084
rect 30380 13636 30436 13646
rect 29184 12572 29448 12582
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29184 12506 29448 12516
rect 29184 11004 29448 11014
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29184 10938 29448 10948
rect 28476 10658 28532 10668
rect 29184 9436 29448 9446
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29184 9370 29448 9380
rect 29184 7868 29448 7878
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29184 7802 29448 7812
rect 29184 6300 29448 6310
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29184 6234 29448 6244
rect 29036 5012 29092 5022
rect 28476 4226 28532 4238
rect 28924 4228 28980 4238
rect 28476 4174 28478 4226
rect 28530 4174 28532 4226
rect 28476 3556 28532 4174
rect 28812 4226 28980 4228
rect 28812 4174 28926 4226
rect 28978 4174 28980 4226
rect 28812 4172 28980 4174
rect 28588 3556 28644 3566
rect 28476 3554 28644 3556
rect 28476 3502 28590 3554
rect 28642 3502 28644 3554
rect 28476 3500 28644 3502
rect 28364 3444 28420 3454
rect 28252 3442 28420 3444
rect 28252 3390 28366 3442
rect 28418 3390 28420 3442
rect 28252 3388 28420 3390
rect 28364 3378 28420 3388
rect 28588 3444 28644 3500
rect 28812 3556 28868 4172
rect 28924 4162 28980 4172
rect 28812 3490 28868 3500
rect 28588 3378 28644 3388
rect 29036 3330 29092 4956
rect 29184 4732 29448 4742
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29184 4666 29448 4676
rect 29596 4620 29988 4676
rect 29484 4564 29540 4574
rect 29596 4564 29652 4620
rect 29484 4562 29652 4564
rect 29484 4510 29486 4562
rect 29538 4510 29652 4562
rect 29484 4508 29652 4510
rect 29484 4498 29540 4508
rect 29708 4452 29764 4462
rect 29372 3444 29428 3454
rect 29372 3350 29428 3388
rect 29596 3444 29652 3454
rect 29036 3278 29038 3330
rect 29090 3278 29092 3330
rect 29036 3266 29092 3278
rect 29184 3164 29448 3174
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 28140 3052 28308 3108
rect 29184 3098 29448 3108
rect 26908 800 26964 2940
rect 27580 800 27636 3052
rect 28252 800 28308 3052
rect 28924 2882 28980 2894
rect 28924 2830 28926 2882
rect 28978 2830 28980 2882
rect 28924 800 28980 2830
rect 29596 800 29652 3388
rect 29708 3442 29764 4396
rect 29708 3390 29710 3442
rect 29762 3390 29764 3442
rect 29708 3378 29764 3390
rect 29932 3554 29988 4620
rect 29932 3502 29934 3554
rect 29986 3502 29988 3554
rect 29932 2882 29988 3502
rect 30156 4226 30212 4238
rect 30156 4174 30158 4226
rect 30210 4174 30212 4226
rect 30156 3444 30212 4174
rect 30156 3378 30212 3388
rect 30380 3442 30436 13580
rect 30828 4226 30884 4238
rect 30828 4174 30830 4226
rect 30882 4174 30884 4226
rect 30380 3390 30382 3442
rect 30434 3390 30436 3442
rect 30380 3378 30436 3390
rect 30604 3554 30660 3566
rect 30604 3502 30606 3554
rect 30658 3502 30660 3554
rect 30604 3444 30660 3502
rect 30604 3378 30660 3388
rect 30828 3220 30884 4174
rect 31052 3442 31108 14476
rect 33846 13356 34110 13366
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 33846 13290 34110 13300
rect 37212 12852 37268 12862
rect 37212 12758 37268 12796
rect 36540 12740 36596 12750
rect 36540 12646 36596 12684
rect 37212 12068 37268 12078
rect 37212 11974 37268 12012
rect 37436 11956 37492 16940
rect 37548 16902 37604 16940
rect 37884 16994 37940 17006
rect 37884 16942 37886 16994
rect 37938 16942 37940 16994
rect 37884 16772 37940 16942
rect 37884 16706 37940 16716
rect 38220 16884 38276 16894
rect 38220 16212 38276 16828
rect 38220 16146 38276 16156
rect 38220 15986 38276 15998
rect 38220 15934 38222 15986
rect 38274 15934 38276 15986
rect 37660 15874 37716 15886
rect 37660 15822 37662 15874
rect 37714 15822 37716 15874
rect 37660 15540 37716 15822
rect 37884 15876 37940 15886
rect 37884 15782 37940 15820
rect 37660 15474 37716 15484
rect 38220 15540 38276 15934
rect 38508 15708 38772 15718
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38508 15642 38772 15652
rect 38220 15474 38276 15484
rect 37884 15428 37940 15438
rect 37884 15334 37940 15372
rect 38220 15314 38276 15326
rect 38220 15262 38222 15314
rect 38274 15262 38276 15314
rect 37660 15204 37716 15214
rect 38220 15204 38276 15262
rect 37660 15202 38276 15204
rect 37660 15150 37662 15202
rect 37714 15150 38276 15202
rect 37660 15148 38276 15150
rect 37660 15138 37716 15148
rect 38220 14868 38276 15148
rect 38220 14802 38276 14812
rect 37660 14420 37716 14430
rect 37660 14326 37716 14364
rect 38220 14418 38276 14430
rect 38220 14366 38222 14418
rect 38274 14366 38276 14418
rect 37884 14308 37940 14318
rect 37884 14214 37940 14252
rect 38220 14308 38276 14366
rect 38220 14242 38276 14252
rect 38508 14140 38772 14150
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38508 14074 38772 14084
rect 37884 13972 37940 13982
rect 37884 13878 37940 13916
rect 38220 13746 38276 13758
rect 38220 13694 38222 13746
rect 38274 13694 38276 13746
rect 37660 13634 37716 13646
rect 37660 13582 37662 13634
rect 37714 13582 37716 13634
rect 37660 13524 37716 13582
rect 37660 13458 37716 13468
rect 38220 13524 38276 13694
rect 38220 13458 38276 13468
rect 37884 12964 37940 12974
rect 37548 12850 37604 12862
rect 37548 12798 37550 12850
rect 37602 12798 37604 12850
rect 37548 12180 37604 12798
rect 37884 12850 37940 12908
rect 37884 12798 37886 12850
rect 37938 12798 37940 12850
rect 37884 12786 37940 12798
rect 38220 12852 38276 12862
rect 38220 12758 38276 12796
rect 38508 12572 38772 12582
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38508 12506 38772 12516
rect 37884 12292 37940 12302
rect 37884 12198 37940 12236
rect 37548 12086 37604 12124
rect 38220 12178 38276 12190
rect 38220 12126 38222 12178
rect 38274 12126 38276 12178
rect 38220 12068 38276 12126
rect 37436 11900 37940 11956
rect 33846 11788 34110 11798
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 33846 11722 34110 11732
rect 37884 11282 37940 11900
rect 38220 11508 38276 12012
rect 38220 11442 38276 11452
rect 37884 11230 37886 11282
rect 37938 11230 37940 11282
rect 37884 11218 37940 11230
rect 38220 11282 38276 11294
rect 38220 11230 38222 11282
rect 38274 11230 38276 11282
rect 37660 11170 37716 11182
rect 37660 11118 37662 11170
rect 37714 11118 37716 11170
rect 37660 10836 37716 11118
rect 37660 10770 37716 10780
rect 38220 10836 38276 11230
rect 38508 11004 38772 11014
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38508 10938 38772 10948
rect 38220 10770 38276 10780
rect 37884 10724 37940 10734
rect 37884 10630 37940 10668
rect 37660 10612 37716 10622
rect 37660 10518 37716 10556
rect 38220 10612 38276 10622
rect 33846 10220 34110 10230
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 33846 10154 34110 10164
rect 38220 10164 38276 10556
rect 38220 10098 38276 10108
rect 38508 9436 38772 9446
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38508 9370 38772 9380
rect 33846 8652 34110 8662
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 33846 8586 34110 8596
rect 38508 7868 38772 7878
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38508 7802 38772 7812
rect 33846 7084 34110 7094
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 33846 7018 34110 7028
rect 38508 6300 38772 6310
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38508 6234 38772 6244
rect 33846 5516 34110 5526
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 33846 5450 34110 5460
rect 38508 4732 38772 4742
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38508 4666 38772 4676
rect 33846 3948 34110 3958
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 33846 3882 34110 3892
rect 31052 3390 31054 3442
rect 31106 3390 31108 3442
rect 31052 3378 31108 3390
rect 31276 3554 31332 3566
rect 31276 3502 31278 3554
rect 31330 3502 31332 3554
rect 31276 3220 31332 3502
rect 30828 3164 31332 3220
rect 29932 2830 29934 2882
rect 29986 2830 29988 2882
rect 29932 2818 29988 2830
rect 30268 924 30660 980
rect 30268 800 30324 924
rect 12096 0 12208 800
rect 12768 0 12880 800
rect 13440 0 13552 800
rect 14112 0 14224 800
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 22176 0 22288 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
rect 25536 0 25648 800
rect 26208 0 26320 800
rect 26880 0 26992 800
rect 27552 0 27664 800
rect 28224 0 28336 800
rect 28896 0 29008 800
rect 29568 0 29680 800
rect 30240 0 30352 800
rect 30604 756 30660 924
rect 31276 756 31332 3164
rect 38508 3164 38772 3174
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38508 3098 38772 3108
rect 30604 700 31332 756
<< via2 >>
rect 5874 36874 5930 36876
rect 5874 36822 5876 36874
rect 5876 36822 5928 36874
rect 5928 36822 5930 36874
rect 5874 36820 5930 36822
rect 5978 36874 6034 36876
rect 5978 36822 5980 36874
rect 5980 36822 6032 36874
rect 6032 36822 6034 36874
rect 5978 36820 6034 36822
rect 6082 36874 6138 36876
rect 6082 36822 6084 36874
rect 6084 36822 6136 36874
rect 6136 36822 6138 36874
rect 10780 36876 10836 36932
rect 6082 36820 6138 36822
rect 11452 36876 11508 36932
rect 10668 36370 10724 36372
rect 10668 36318 10670 36370
rect 10670 36318 10722 36370
rect 10722 36318 10724 36370
rect 10668 36316 10724 36318
rect 10536 36090 10592 36092
rect 10536 36038 10538 36090
rect 10538 36038 10590 36090
rect 10590 36038 10592 36090
rect 10536 36036 10592 36038
rect 10640 36090 10696 36092
rect 10640 36038 10642 36090
rect 10642 36038 10694 36090
rect 10694 36038 10696 36090
rect 10640 36036 10696 36038
rect 10744 36090 10800 36092
rect 10744 36038 10746 36090
rect 10746 36038 10798 36090
rect 10798 36038 10800 36090
rect 10744 36036 10800 36038
rect 5874 35306 5930 35308
rect 5874 35254 5876 35306
rect 5876 35254 5928 35306
rect 5928 35254 5930 35306
rect 5874 35252 5930 35254
rect 5978 35306 6034 35308
rect 5978 35254 5980 35306
rect 5980 35254 6032 35306
rect 6032 35254 6034 35306
rect 5978 35252 6034 35254
rect 6082 35306 6138 35308
rect 6082 35254 6084 35306
rect 6084 35254 6136 35306
rect 6136 35254 6138 35306
rect 6082 35252 6138 35254
rect 10536 34522 10592 34524
rect 10536 34470 10538 34522
rect 10538 34470 10590 34522
rect 10590 34470 10592 34522
rect 10536 34468 10592 34470
rect 10640 34522 10696 34524
rect 10640 34470 10642 34522
rect 10642 34470 10694 34522
rect 10694 34470 10696 34522
rect 10640 34468 10696 34470
rect 10744 34522 10800 34524
rect 10744 34470 10746 34522
rect 10746 34470 10798 34522
rect 10798 34470 10800 34522
rect 10744 34468 10800 34470
rect 5874 33738 5930 33740
rect 5874 33686 5876 33738
rect 5876 33686 5928 33738
rect 5928 33686 5930 33738
rect 5874 33684 5930 33686
rect 5978 33738 6034 33740
rect 5978 33686 5980 33738
rect 5980 33686 6032 33738
rect 6032 33686 6034 33738
rect 5978 33684 6034 33686
rect 6082 33738 6138 33740
rect 6082 33686 6084 33738
rect 6084 33686 6136 33738
rect 6136 33686 6138 33738
rect 6082 33684 6138 33686
rect 10536 32954 10592 32956
rect 10536 32902 10538 32954
rect 10538 32902 10590 32954
rect 10590 32902 10592 32954
rect 10536 32900 10592 32902
rect 10640 32954 10696 32956
rect 10640 32902 10642 32954
rect 10642 32902 10694 32954
rect 10694 32902 10696 32954
rect 10640 32900 10696 32902
rect 10744 32954 10800 32956
rect 10744 32902 10746 32954
rect 10746 32902 10798 32954
rect 10798 32902 10800 32954
rect 10744 32900 10800 32902
rect 5874 32170 5930 32172
rect 5874 32118 5876 32170
rect 5876 32118 5928 32170
rect 5928 32118 5930 32170
rect 5874 32116 5930 32118
rect 5978 32170 6034 32172
rect 5978 32118 5980 32170
rect 5980 32118 6032 32170
rect 6032 32118 6034 32170
rect 5978 32116 6034 32118
rect 6082 32170 6138 32172
rect 6082 32118 6084 32170
rect 6084 32118 6136 32170
rect 6136 32118 6138 32170
rect 6082 32116 6138 32118
rect 11676 36316 11732 36372
rect 11900 36258 11956 36260
rect 11900 36206 11902 36258
rect 11902 36206 11954 36258
rect 11954 36206 11956 36258
rect 11900 36204 11956 36206
rect 10536 31386 10592 31388
rect 10536 31334 10538 31386
rect 10538 31334 10590 31386
rect 10590 31334 10592 31386
rect 10536 31332 10592 31334
rect 10640 31386 10696 31388
rect 10640 31334 10642 31386
rect 10642 31334 10694 31386
rect 10694 31334 10696 31386
rect 10640 31332 10696 31334
rect 10744 31386 10800 31388
rect 10744 31334 10746 31386
rect 10746 31334 10798 31386
rect 10798 31334 10800 31386
rect 10744 31332 10800 31334
rect 5874 30602 5930 30604
rect 5874 30550 5876 30602
rect 5876 30550 5928 30602
rect 5928 30550 5930 30602
rect 5874 30548 5930 30550
rect 5978 30602 6034 30604
rect 5978 30550 5980 30602
rect 5980 30550 6032 30602
rect 6032 30550 6034 30602
rect 5978 30548 6034 30550
rect 6082 30602 6138 30604
rect 6082 30550 6084 30602
rect 6084 30550 6136 30602
rect 6136 30550 6138 30602
rect 6082 30548 6138 30550
rect 10536 29818 10592 29820
rect 10536 29766 10538 29818
rect 10538 29766 10590 29818
rect 10590 29766 10592 29818
rect 10536 29764 10592 29766
rect 10640 29818 10696 29820
rect 10640 29766 10642 29818
rect 10642 29766 10694 29818
rect 10694 29766 10696 29818
rect 10640 29764 10696 29766
rect 10744 29818 10800 29820
rect 10744 29766 10746 29818
rect 10746 29766 10798 29818
rect 10798 29766 10800 29818
rect 10744 29764 10800 29766
rect 4284 29426 4340 29428
rect 4284 29374 4286 29426
rect 4286 29374 4338 29426
rect 4338 29374 4340 29426
rect 4284 29372 4340 29374
rect 1932 29202 1988 29204
rect 1932 29150 1934 29202
rect 1934 29150 1986 29202
rect 1986 29150 1988 29202
rect 1932 29148 1988 29150
rect 5874 29034 5930 29036
rect 5874 28982 5876 29034
rect 5876 28982 5928 29034
rect 5928 28982 5930 29034
rect 5874 28980 5930 28982
rect 5978 29034 6034 29036
rect 5978 28982 5980 29034
rect 5980 28982 6032 29034
rect 6032 28982 6034 29034
rect 5978 28980 6034 28982
rect 6082 29034 6138 29036
rect 6082 28982 6084 29034
rect 6084 28982 6136 29034
rect 6136 28982 6138 29034
rect 6082 28980 6138 28982
rect 1708 28252 1764 28308
rect 2492 28252 2548 28308
rect 10536 28250 10592 28252
rect 10536 28198 10538 28250
rect 10538 28198 10590 28250
rect 10590 28198 10592 28250
rect 10536 28196 10592 28198
rect 10640 28250 10696 28252
rect 10640 28198 10642 28250
rect 10642 28198 10694 28250
rect 10694 28198 10696 28250
rect 10640 28196 10696 28198
rect 10744 28250 10800 28252
rect 10744 28198 10746 28250
rect 10746 28198 10798 28250
rect 10798 28198 10800 28250
rect 10744 28196 10800 28198
rect 1708 27580 1764 27636
rect 2044 27244 2100 27300
rect 2380 26962 2436 26964
rect 2380 26910 2382 26962
rect 2382 26910 2434 26962
rect 2434 26910 2436 26962
rect 2380 26908 2436 26910
rect 2044 26402 2100 26404
rect 2044 26350 2046 26402
rect 2046 26350 2098 26402
rect 2098 26350 2100 26402
rect 2044 26348 2100 26350
rect 1820 26236 1876 26292
rect 1708 26124 1764 26180
rect 2492 26178 2548 26180
rect 2492 26126 2494 26178
rect 2494 26126 2546 26178
rect 2546 26126 2548 26178
rect 2492 26124 2548 26126
rect 1708 25564 1764 25620
rect 2044 25282 2100 25284
rect 2044 25230 2046 25282
rect 2046 25230 2098 25282
rect 2098 25230 2100 25282
rect 2044 25228 2100 25230
rect 1708 24892 1764 24948
rect 2492 24892 2548 24948
rect 1708 24220 1764 24276
rect 2044 23714 2100 23716
rect 2044 23662 2046 23714
rect 2046 23662 2098 23714
rect 2098 23662 2100 23714
rect 2044 23660 2100 23662
rect 1708 23548 1764 23604
rect 2044 23266 2100 23268
rect 2044 23214 2046 23266
rect 2046 23214 2098 23266
rect 2098 23214 2100 23266
rect 2044 23212 2100 23214
rect 1708 22876 1764 22932
rect 2044 22316 2100 22372
rect 1708 22258 1764 22260
rect 1708 22206 1710 22258
rect 1710 22206 1762 22258
rect 1762 22206 1764 22258
rect 1708 22204 1764 22206
rect 2044 21698 2100 21700
rect 2044 21646 2046 21698
rect 2046 21646 2098 21698
rect 2098 21646 2100 21698
rect 2044 21644 2100 21646
rect 1708 21420 1764 21476
rect 1708 20860 1764 20916
rect 2492 24220 2548 24276
rect 2492 23548 2548 23604
rect 2492 22876 2548 22932
rect 2492 22204 2548 22260
rect 2380 21532 2436 21588
rect 2716 23996 2772 24052
rect 2604 21308 2660 21364
rect 1708 20188 1764 20244
rect 2044 20130 2100 20132
rect 2044 20078 2046 20130
rect 2046 20078 2098 20130
rect 2098 20078 2100 20130
rect 2044 20076 2100 20078
rect 2268 20524 2324 20580
rect 2492 20188 2548 20244
rect 2156 19740 2212 19796
rect 1708 19516 1764 19572
rect 2492 19516 2548 19572
rect 2940 27580 2996 27636
rect 5874 27466 5930 27468
rect 5874 27414 5876 27466
rect 5876 27414 5928 27466
rect 5928 27414 5930 27466
rect 5874 27412 5930 27414
rect 5978 27466 6034 27468
rect 5978 27414 5980 27466
rect 5980 27414 6032 27466
rect 6032 27414 6034 27466
rect 5978 27412 6034 27414
rect 6082 27466 6138 27468
rect 6082 27414 6084 27466
rect 6084 27414 6136 27466
rect 6136 27414 6138 27466
rect 6082 27412 6138 27414
rect 3164 26962 3220 26964
rect 3164 26910 3166 26962
rect 3166 26910 3218 26962
rect 3218 26910 3220 26962
rect 3164 26908 3220 26910
rect 10536 26682 10592 26684
rect 10536 26630 10538 26682
rect 10538 26630 10590 26682
rect 10590 26630 10592 26682
rect 10536 26628 10592 26630
rect 10640 26682 10696 26684
rect 10640 26630 10642 26682
rect 10642 26630 10694 26682
rect 10694 26630 10696 26682
rect 10640 26628 10696 26630
rect 10744 26682 10800 26684
rect 10744 26630 10746 26682
rect 10746 26630 10798 26682
rect 10798 26630 10800 26682
rect 10744 26628 10800 26630
rect 15198 36874 15254 36876
rect 15198 36822 15200 36874
rect 15200 36822 15252 36874
rect 15252 36822 15254 36874
rect 15198 36820 15254 36822
rect 15302 36874 15358 36876
rect 15302 36822 15304 36874
rect 15304 36822 15356 36874
rect 15356 36822 15358 36874
rect 15302 36820 15358 36822
rect 15406 36874 15462 36876
rect 15406 36822 15408 36874
rect 15408 36822 15460 36874
rect 15460 36822 15462 36874
rect 15406 36820 15462 36822
rect 16156 36652 16212 36708
rect 12572 27132 12628 27188
rect 11228 26460 11284 26516
rect 12572 26908 12628 26964
rect 5874 25898 5930 25900
rect 5874 25846 5876 25898
rect 5876 25846 5928 25898
rect 5928 25846 5930 25898
rect 5874 25844 5930 25846
rect 5978 25898 6034 25900
rect 5978 25846 5980 25898
rect 5980 25846 6032 25898
rect 6032 25846 6034 25898
rect 5978 25844 6034 25846
rect 6082 25898 6138 25900
rect 6082 25846 6084 25898
rect 6084 25846 6136 25898
rect 6136 25846 6138 25898
rect 6082 25844 6138 25846
rect 12348 25228 12404 25284
rect 10536 25114 10592 25116
rect 10536 25062 10538 25114
rect 10538 25062 10590 25114
rect 10590 25062 10592 25114
rect 10536 25060 10592 25062
rect 10640 25114 10696 25116
rect 10640 25062 10642 25114
rect 10642 25062 10694 25114
rect 10694 25062 10696 25114
rect 10640 25060 10696 25062
rect 10744 25114 10800 25116
rect 10744 25062 10746 25114
rect 10746 25062 10798 25114
rect 10798 25062 10800 25114
rect 10744 25060 10800 25062
rect 12460 24444 12516 24500
rect 5874 24330 5930 24332
rect 5874 24278 5876 24330
rect 5876 24278 5928 24330
rect 5928 24278 5930 24330
rect 5874 24276 5930 24278
rect 5978 24330 6034 24332
rect 5978 24278 5980 24330
rect 5980 24278 6032 24330
rect 6032 24278 6034 24330
rect 5978 24276 6034 24278
rect 6082 24330 6138 24332
rect 6082 24278 6084 24330
rect 6084 24278 6136 24330
rect 6136 24278 6138 24330
rect 6082 24276 6138 24278
rect 10536 23546 10592 23548
rect 10536 23494 10538 23546
rect 10538 23494 10590 23546
rect 10590 23494 10592 23546
rect 10536 23492 10592 23494
rect 10640 23546 10696 23548
rect 10640 23494 10642 23546
rect 10642 23494 10694 23546
rect 10694 23494 10696 23546
rect 10640 23492 10696 23494
rect 10744 23546 10800 23548
rect 10744 23494 10746 23546
rect 10746 23494 10798 23546
rect 10798 23494 10800 23546
rect 10744 23492 10800 23494
rect 12348 23548 12404 23604
rect 5874 22762 5930 22764
rect 5874 22710 5876 22762
rect 5876 22710 5928 22762
rect 5928 22710 5930 22762
rect 5874 22708 5930 22710
rect 5978 22762 6034 22764
rect 5978 22710 5980 22762
rect 5980 22710 6032 22762
rect 6032 22710 6034 22762
rect 5978 22708 6034 22710
rect 6082 22762 6138 22764
rect 6082 22710 6084 22762
rect 6084 22710 6136 22762
rect 6136 22710 6138 22762
rect 6082 22708 6138 22710
rect 10536 21978 10592 21980
rect 10536 21926 10538 21978
rect 10538 21926 10590 21978
rect 10590 21926 10592 21978
rect 10536 21924 10592 21926
rect 10640 21978 10696 21980
rect 10640 21926 10642 21978
rect 10642 21926 10694 21978
rect 10694 21926 10696 21978
rect 10640 21924 10696 21926
rect 10744 21978 10800 21980
rect 10744 21926 10746 21978
rect 10746 21926 10798 21978
rect 10798 21926 10800 21978
rect 10744 21924 10800 21926
rect 3164 21532 3220 21588
rect 12236 21644 12292 21700
rect 2940 21474 2996 21476
rect 2940 21422 2942 21474
rect 2942 21422 2994 21474
rect 2994 21422 2996 21474
rect 2940 21420 2996 21422
rect 12124 21308 12180 21364
rect 5874 21194 5930 21196
rect 5874 21142 5876 21194
rect 5876 21142 5928 21194
rect 5928 21142 5930 21194
rect 5874 21140 5930 21142
rect 5978 21194 6034 21196
rect 5978 21142 5980 21194
rect 5980 21142 6032 21194
rect 6032 21142 6034 21194
rect 5978 21140 6034 21142
rect 6082 21194 6138 21196
rect 6082 21142 6084 21194
rect 6084 21142 6136 21194
rect 6136 21142 6138 21194
rect 6082 21140 6138 21142
rect 2828 20860 2884 20916
rect 11340 20802 11396 20804
rect 11340 20750 11342 20802
rect 11342 20750 11394 20802
rect 11394 20750 11396 20802
rect 11340 20748 11396 20750
rect 11788 20690 11844 20692
rect 11788 20638 11790 20690
rect 11790 20638 11842 20690
rect 11842 20638 11844 20690
rect 11788 20636 11844 20638
rect 10536 20410 10592 20412
rect 10536 20358 10538 20410
rect 10538 20358 10590 20410
rect 10590 20358 10592 20410
rect 10536 20356 10592 20358
rect 10640 20410 10696 20412
rect 10640 20358 10642 20410
rect 10642 20358 10694 20410
rect 10694 20358 10696 20410
rect 10640 20356 10696 20358
rect 10744 20410 10800 20412
rect 10744 20358 10746 20410
rect 10746 20358 10798 20410
rect 10798 20358 10800 20410
rect 10744 20356 10800 20358
rect 12236 20076 12292 20132
rect 5874 19626 5930 19628
rect 5874 19574 5876 19626
rect 5876 19574 5928 19626
rect 5928 19574 5930 19626
rect 5874 19572 5930 19574
rect 5978 19626 6034 19628
rect 5978 19574 5980 19626
rect 5980 19574 6032 19626
rect 6032 19574 6034 19626
rect 5978 19572 6034 19574
rect 6082 19626 6138 19628
rect 6082 19574 6084 19626
rect 6084 19574 6136 19626
rect 6136 19574 6138 19626
rect 6082 19572 6138 19574
rect 2716 19292 2772 19348
rect 12460 20914 12516 20916
rect 12460 20862 12462 20914
rect 12462 20862 12514 20914
rect 12514 20862 12516 20914
rect 12460 20860 12516 20862
rect 4284 19234 4340 19236
rect 4284 19182 4286 19234
rect 4286 19182 4338 19234
rect 4338 19182 4340 19234
rect 4284 19180 4340 19182
rect 12908 25340 12964 25396
rect 13132 24722 13188 24724
rect 13132 24670 13134 24722
rect 13134 24670 13186 24722
rect 13186 24670 13188 24722
rect 13132 24668 13188 24670
rect 13580 27244 13636 27300
rect 13692 25340 13748 25396
rect 14364 29148 14420 29204
rect 15198 35306 15254 35308
rect 15198 35254 15200 35306
rect 15200 35254 15252 35306
rect 15252 35254 15254 35306
rect 15198 35252 15254 35254
rect 15302 35306 15358 35308
rect 15302 35254 15304 35306
rect 15304 35254 15356 35306
rect 15356 35254 15358 35306
rect 15302 35252 15358 35254
rect 15406 35306 15462 35308
rect 15406 35254 15408 35306
rect 15408 35254 15460 35306
rect 15460 35254 15462 35306
rect 15406 35252 15462 35254
rect 15198 33738 15254 33740
rect 15198 33686 15200 33738
rect 15200 33686 15252 33738
rect 15252 33686 15254 33738
rect 15198 33684 15254 33686
rect 15302 33738 15358 33740
rect 15302 33686 15304 33738
rect 15304 33686 15356 33738
rect 15356 33686 15358 33738
rect 15302 33684 15358 33686
rect 15406 33738 15462 33740
rect 15406 33686 15408 33738
rect 15408 33686 15460 33738
rect 15460 33686 15462 33738
rect 15406 33684 15462 33686
rect 15198 32170 15254 32172
rect 15198 32118 15200 32170
rect 15200 32118 15252 32170
rect 15252 32118 15254 32170
rect 15198 32116 15254 32118
rect 15302 32170 15358 32172
rect 15302 32118 15304 32170
rect 15304 32118 15356 32170
rect 15356 32118 15358 32170
rect 15302 32116 15358 32118
rect 15406 32170 15462 32172
rect 15406 32118 15408 32170
rect 15408 32118 15460 32170
rect 15460 32118 15462 32170
rect 15406 32116 15462 32118
rect 15198 30602 15254 30604
rect 15198 30550 15200 30602
rect 15200 30550 15252 30602
rect 15252 30550 15254 30602
rect 15198 30548 15254 30550
rect 15302 30602 15358 30604
rect 15302 30550 15304 30602
rect 15304 30550 15356 30602
rect 15356 30550 15358 30602
rect 15302 30548 15358 30550
rect 15406 30602 15462 30604
rect 15406 30550 15408 30602
rect 15408 30550 15460 30602
rect 15460 30550 15462 30602
rect 15406 30548 15462 30550
rect 16156 36482 16212 36484
rect 16156 36430 16158 36482
rect 16158 36430 16210 36482
rect 16210 36430 16212 36482
rect 16156 36428 16212 36430
rect 16492 36428 16548 36484
rect 15820 29148 15876 29204
rect 15198 29034 15254 29036
rect 15198 28982 15200 29034
rect 15200 28982 15252 29034
rect 15252 28982 15254 29034
rect 15198 28980 15254 28982
rect 15302 29034 15358 29036
rect 15302 28982 15304 29034
rect 15304 28982 15356 29034
rect 15356 28982 15358 29034
rect 15302 28980 15358 28982
rect 15406 29034 15462 29036
rect 15406 28982 15408 29034
rect 15408 28982 15460 29034
rect 15460 28982 15462 29034
rect 15406 28980 15462 28982
rect 15036 28812 15092 28868
rect 15708 28812 15764 28868
rect 15036 27804 15092 27860
rect 15198 27466 15254 27468
rect 15198 27414 15200 27466
rect 15200 27414 15252 27466
rect 15252 27414 15254 27466
rect 15198 27412 15254 27414
rect 15302 27466 15358 27468
rect 15302 27414 15304 27466
rect 15304 27414 15356 27466
rect 15356 27414 15358 27466
rect 15302 27412 15358 27414
rect 15406 27466 15462 27468
rect 15406 27414 15408 27466
rect 15408 27414 15460 27466
rect 15460 27414 15462 27466
rect 15406 27412 15462 27414
rect 14364 26348 14420 26404
rect 14812 26236 14868 26292
rect 15198 25898 15254 25900
rect 15198 25846 15200 25898
rect 15200 25846 15252 25898
rect 15252 25846 15254 25898
rect 15198 25844 15254 25846
rect 15302 25898 15358 25900
rect 15302 25846 15304 25898
rect 15304 25846 15356 25898
rect 15356 25846 15358 25898
rect 15302 25844 15358 25846
rect 15406 25898 15462 25900
rect 15406 25846 15408 25898
rect 15408 25846 15460 25898
rect 15460 25846 15462 25898
rect 15406 25844 15462 25846
rect 13804 24892 13860 24948
rect 15932 29036 15988 29092
rect 14700 24722 14756 24724
rect 14700 24670 14702 24722
rect 14702 24670 14754 24722
rect 14754 24670 14756 24722
rect 14700 24668 14756 24670
rect 13356 24108 13412 24164
rect 14700 24444 14756 24500
rect 14364 23996 14420 24052
rect 15596 24444 15652 24500
rect 15198 24330 15254 24332
rect 15198 24278 15200 24330
rect 15200 24278 15252 24330
rect 15252 24278 15254 24330
rect 15198 24276 15254 24278
rect 15302 24330 15358 24332
rect 15302 24278 15304 24330
rect 15304 24278 15356 24330
rect 15356 24278 15358 24330
rect 15302 24276 15358 24278
rect 15406 24330 15462 24332
rect 15406 24278 15408 24330
rect 15408 24278 15460 24330
rect 15460 24278 15462 24330
rect 15406 24276 15462 24278
rect 13132 23100 13188 23156
rect 13804 23100 13860 23156
rect 13580 22092 13636 22148
rect 14476 21644 14532 21700
rect 12908 20972 12964 21028
rect 15596 23436 15652 23492
rect 15596 23154 15652 23156
rect 15596 23102 15598 23154
rect 15598 23102 15650 23154
rect 15650 23102 15652 23154
rect 15596 23100 15652 23102
rect 15198 22762 15254 22764
rect 15198 22710 15200 22762
rect 15200 22710 15252 22762
rect 15252 22710 15254 22762
rect 15198 22708 15254 22710
rect 15302 22762 15358 22764
rect 15302 22710 15304 22762
rect 15304 22710 15356 22762
rect 15356 22710 15358 22762
rect 15302 22708 15358 22710
rect 15406 22762 15462 22764
rect 15406 22710 15408 22762
rect 15408 22710 15460 22762
rect 15460 22710 15462 22762
rect 15406 22708 15462 22710
rect 15036 22428 15092 22484
rect 13580 20860 13636 20916
rect 13468 20802 13524 20804
rect 13468 20750 13470 20802
rect 13470 20750 13522 20802
rect 13522 20750 13524 20802
rect 13468 20748 13524 20750
rect 12908 19404 12964 19460
rect 1932 18844 1988 18900
rect 10536 18842 10592 18844
rect 10536 18790 10538 18842
rect 10538 18790 10590 18842
rect 10590 18790 10592 18842
rect 10536 18788 10592 18790
rect 10640 18842 10696 18844
rect 10640 18790 10642 18842
rect 10642 18790 10694 18842
rect 10694 18790 10696 18842
rect 10640 18788 10696 18790
rect 10744 18842 10800 18844
rect 10744 18790 10746 18842
rect 10746 18790 10798 18842
rect 10798 18790 10800 18842
rect 10744 18788 10800 18790
rect 2044 18396 2100 18452
rect 1708 18172 1764 18228
rect 2492 18172 2548 18228
rect 13468 19234 13524 19236
rect 13468 19182 13470 19234
rect 13470 19182 13522 19234
rect 13522 19182 13524 19234
rect 13468 19180 13524 19182
rect 15372 21308 15428 21364
rect 17164 36706 17220 36708
rect 17164 36654 17166 36706
rect 17166 36654 17218 36706
rect 17218 36654 17220 36706
rect 17164 36652 17220 36654
rect 16828 36428 16884 36484
rect 18060 35810 18116 35812
rect 18060 35758 18062 35810
rect 18062 35758 18114 35810
rect 18114 35758 18116 35810
rect 18060 35756 18116 35758
rect 17500 27186 17556 27188
rect 17500 27134 17502 27186
rect 17502 27134 17554 27186
rect 17554 27134 17556 27186
rect 17500 27132 17556 27134
rect 16492 27074 16548 27076
rect 16492 27022 16494 27074
rect 16494 27022 16546 27074
rect 16546 27022 16548 27074
rect 16492 27020 16548 27022
rect 17612 27074 17668 27076
rect 17612 27022 17614 27074
rect 17614 27022 17666 27074
rect 17666 27022 17668 27074
rect 17612 27020 17668 27022
rect 20188 36876 20244 36932
rect 20860 36652 20916 36708
rect 21420 36876 21476 36932
rect 16604 26290 16660 26292
rect 16604 26238 16606 26290
rect 16606 26238 16658 26290
rect 16658 26238 16660 26290
rect 16604 26236 16660 26238
rect 16268 24834 16324 24836
rect 16268 24782 16270 24834
rect 16270 24782 16322 24834
rect 16322 24782 16324 24834
rect 16268 24780 16324 24782
rect 16492 25452 16548 25508
rect 16380 23884 16436 23940
rect 15932 22370 15988 22372
rect 15932 22318 15934 22370
rect 15934 22318 15986 22370
rect 15986 22318 15988 22370
rect 15932 22316 15988 22318
rect 15820 21644 15876 21700
rect 15198 21194 15254 21196
rect 15198 21142 15200 21194
rect 15200 21142 15252 21194
rect 15252 21142 15254 21194
rect 15198 21140 15254 21142
rect 15302 21194 15358 21196
rect 15302 21142 15304 21194
rect 15304 21142 15356 21194
rect 15356 21142 15358 21194
rect 15302 21140 15358 21142
rect 15406 21194 15462 21196
rect 15406 21142 15408 21194
rect 15408 21142 15460 21194
rect 15460 21142 15462 21194
rect 15406 21140 15462 21142
rect 17724 26514 17780 26516
rect 17724 26462 17726 26514
rect 17726 26462 17778 26514
rect 17778 26462 17780 26514
rect 17724 26460 17780 26462
rect 17388 25506 17444 25508
rect 17388 25454 17390 25506
rect 17390 25454 17442 25506
rect 17442 25454 17444 25506
rect 17388 25452 17444 25454
rect 17052 25228 17108 25284
rect 18620 25228 18676 25284
rect 17948 24892 18004 24948
rect 16716 24556 16772 24612
rect 17836 24162 17892 24164
rect 17836 24110 17838 24162
rect 17838 24110 17890 24162
rect 17890 24110 17892 24162
rect 17836 24108 17892 24110
rect 16716 24050 16772 24052
rect 16716 23998 16718 24050
rect 16718 23998 16770 24050
rect 16770 23998 16772 24050
rect 16716 23996 16772 23998
rect 17500 23938 17556 23940
rect 17500 23886 17502 23938
rect 17502 23886 17554 23938
rect 17554 23886 17556 23938
rect 17500 23884 17556 23886
rect 19628 36204 19684 36260
rect 19292 35756 19348 35812
rect 18732 23996 18788 24052
rect 16492 23436 16548 23492
rect 17388 23436 17444 23492
rect 16716 23266 16772 23268
rect 16716 23214 16718 23266
rect 16718 23214 16770 23266
rect 16770 23214 16772 23266
rect 16716 23212 16772 23214
rect 17612 22876 17668 22932
rect 16828 22428 16884 22484
rect 17388 22428 17444 22484
rect 16268 20972 16324 21028
rect 15820 20860 15876 20916
rect 15372 20018 15428 20020
rect 15372 19966 15374 20018
rect 15374 19966 15426 20018
rect 15426 19966 15428 20018
rect 15372 19964 15428 19966
rect 16940 20914 16996 20916
rect 16940 20862 16942 20914
rect 16942 20862 16994 20914
rect 16994 20862 16996 20914
rect 16940 20860 16996 20862
rect 16828 20636 16884 20692
rect 15198 19626 15254 19628
rect 15198 19574 15200 19626
rect 15200 19574 15252 19626
rect 15252 19574 15254 19626
rect 15198 19572 15254 19574
rect 15302 19626 15358 19628
rect 15302 19574 15304 19626
rect 15304 19574 15356 19626
rect 15356 19574 15358 19626
rect 15302 19572 15358 19574
rect 15406 19626 15462 19628
rect 15406 19574 15408 19626
rect 15408 19574 15460 19626
rect 15460 19574 15462 19626
rect 15406 19572 15462 19574
rect 14924 18620 14980 18676
rect 12572 18172 12628 18228
rect 13020 18284 13076 18340
rect 5874 18058 5930 18060
rect 5874 18006 5876 18058
rect 5876 18006 5928 18058
rect 5928 18006 5930 18058
rect 5874 18004 5930 18006
rect 5978 18058 6034 18060
rect 5978 18006 5980 18058
rect 5980 18006 6032 18058
rect 6032 18006 6034 18058
rect 5978 18004 6034 18006
rect 6082 18058 6138 18060
rect 6082 18006 6084 18058
rect 6084 18006 6136 18058
rect 6136 18006 6138 18058
rect 6082 18004 6138 18006
rect 12796 17890 12852 17892
rect 12796 17838 12798 17890
rect 12798 17838 12850 17890
rect 12850 17838 12852 17890
rect 12796 17836 12852 17838
rect 1932 17778 1988 17780
rect 1932 17726 1934 17778
rect 1934 17726 1986 17778
rect 1986 17726 1988 17778
rect 1932 17724 1988 17726
rect 2156 17724 2212 17780
rect 2716 17612 2772 17668
rect 1708 16882 1764 16884
rect 1708 16830 1710 16882
rect 1710 16830 1762 16882
rect 1762 16830 1764 16882
rect 1708 16828 1764 16830
rect 1708 15484 1764 15540
rect 1708 14812 1764 14868
rect 2380 16716 2436 16772
rect 2044 16268 2100 16324
rect 2268 16604 2324 16660
rect 2044 15874 2100 15876
rect 2044 15822 2046 15874
rect 2046 15822 2098 15874
rect 2098 15822 2100 15874
rect 2044 15820 2100 15822
rect 2044 15426 2100 15428
rect 2044 15374 2046 15426
rect 2046 15374 2098 15426
rect 2098 15374 2100 15426
rect 2044 15372 2100 15374
rect 1708 14140 1764 14196
rect 2380 16156 2436 16212
rect 2492 16828 2548 16884
rect 3164 16716 3220 16772
rect 11788 17612 11844 17668
rect 12236 17666 12292 17668
rect 12236 17614 12238 17666
rect 12238 17614 12290 17666
rect 12290 17614 12292 17666
rect 12236 17612 12292 17614
rect 13468 17836 13524 17892
rect 13804 17724 13860 17780
rect 14028 17666 14084 17668
rect 14028 17614 14030 17666
rect 14030 17614 14082 17666
rect 14082 17614 14084 17666
rect 14028 17612 14084 17614
rect 10536 17274 10592 17276
rect 10536 17222 10538 17274
rect 10538 17222 10590 17274
rect 10590 17222 10592 17274
rect 10536 17220 10592 17222
rect 10640 17274 10696 17276
rect 10640 17222 10642 17274
rect 10642 17222 10694 17274
rect 10694 17222 10696 17274
rect 10640 17220 10696 17222
rect 10744 17274 10800 17276
rect 10744 17222 10746 17274
rect 10746 17222 10798 17274
rect 10798 17222 10800 17274
rect 10744 17220 10800 17222
rect 12460 16770 12516 16772
rect 12460 16718 12462 16770
rect 12462 16718 12514 16770
rect 12514 16718 12516 16770
rect 12460 16716 12516 16718
rect 4284 16604 4340 16660
rect 5874 16490 5930 16492
rect 5874 16438 5876 16490
rect 5876 16438 5928 16490
rect 5928 16438 5930 16490
rect 5874 16436 5930 16438
rect 5978 16490 6034 16492
rect 5978 16438 5980 16490
rect 5980 16438 6032 16490
rect 6032 16438 6034 16490
rect 5978 16436 6034 16438
rect 6082 16490 6138 16492
rect 6082 16438 6084 16490
rect 6084 16438 6136 16490
rect 6136 16438 6138 16490
rect 6082 16436 6138 16438
rect 13132 16882 13188 16884
rect 13132 16830 13134 16882
rect 13134 16830 13186 16882
rect 13186 16830 13188 16882
rect 13132 16828 13188 16830
rect 13916 16658 13972 16660
rect 13916 16606 13918 16658
rect 13918 16606 13970 16658
rect 13970 16606 13972 16658
rect 13916 16604 13972 16606
rect 12796 16380 12852 16436
rect 14140 16380 14196 16436
rect 13804 16210 13860 16212
rect 13804 16158 13806 16210
rect 13806 16158 13858 16210
rect 13858 16158 13860 16210
rect 13804 16156 13860 16158
rect 10536 15706 10592 15708
rect 10536 15654 10538 15706
rect 10538 15654 10590 15706
rect 10590 15654 10592 15706
rect 10536 15652 10592 15654
rect 10640 15706 10696 15708
rect 10640 15654 10642 15706
rect 10642 15654 10694 15706
rect 10694 15654 10696 15706
rect 10640 15652 10696 15654
rect 10744 15706 10800 15708
rect 10744 15654 10746 15706
rect 10746 15654 10798 15706
rect 10798 15654 10800 15706
rect 10744 15652 10800 15654
rect 2940 15484 2996 15540
rect 14140 15372 14196 15428
rect 14924 18284 14980 18340
rect 15198 18058 15254 18060
rect 15198 18006 15200 18058
rect 15200 18006 15252 18058
rect 15252 18006 15254 18058
rect 15198 18004 15254 18006
rect 15302 18058 15358 18060
rect 15302 18006 15304 18058
rect 15304 18006 15356 18058
rect 15356 18006 15358 18058
rect 15302 18004 15358 18006
rect 15406 18058 15462 18060
rect 15406 18006 15408 18058
rect 15408 18006 15460 18058
rect 15460 18006 15462 18058
rect 15406 18004 15462 18006
rect 14700 16882 14756 16884
rect 14700 16830 14702 16882
rect 14702 16830 14754 16882
rect 14754 16830 14756 16882
rect 14700 16828 14756 16830
rect 14252 16044 14308 16100
rect 14028 15314 14084 15316
rect 14028 15262 14030 15314
rect 14030 15262 14082 15314
rect 14082 15262 14084 15314
rect 14028 15260 14084 15262
rect 15198 16490 15254 16492
rect 15198 16438 15200 16490
rect 15200 16438 15252 16490
rect 15252 16438 15254 16490
rect 15198 16436 15254 16438
rect 15302 16490 15358 16492
rect 15302 16438 15304 16490
rect 15304 16438 15356 16490
rect 15356 16438 15358 16490
rect 15302 16436 15358 16438
rect 15406 16490 15462 16492
rect 15406 16438 15408 16490
rect 15408 16438 15460 16490
rect 15460 16438 15462 16490
rect 15406 16436 15462 16438
rect 15820 18284 15876 18340
rect 15148 16098 15204 16100
rect 15148 16046 15150 16098
rect 15150 16046 15202 16098
rect 15202 16046 15204 16098
rect 15148 16044 15204 16046
rect 15372 15820 15428 15876
rect 2492 14812 2548 14868
rect 5874 14922 5930 14924
rect 5874 14870 5876 14922
rect 5876 14870 5928 14922
rect 5928 14870 5930 14922
rect 5874 14868 5930 14870
rect 5978 14922 6034 14924
rect 5978 14870 5980 14922
rect 5980 14870 6032 14922
rect 6032 14870 6034 14922
rect 5978 14868 6034 14870
rect 6082 14922 6138 14924
rect 6082 14870 6084 14922
rect 6084 14870 6136 14922
rect 6136 14870 6138 14922
rect 6082 14868 6138 14870
rect 15198 14922 15254 14924
rect 15198 14870 15200 14922
rect 15200 14870 15252 14922
rect 15252 14870 15254 14922
rect 15198 14868 15254 14870
rect 15302 14922 15358 14924
rect 15302 14870 15304 14922
rect 15304 14870 15356 14922
rect 15356 14870 15358 14922
rect 15302 14868 15358 14870
rect 15406 14922 15462 14924
rect 15406 14870 15408 14922
rect 15408 14870 15460 14922
rect 15460 14870 15462 14922
rect 15406 14868 15462 14870
rect 2492 14140 2548 14196
rect 10536 14138 10592 14140
rect 10536 14086 10538 14138
rect 10538 14086 10590 14138
rect 10590 14086 10592 14138
rect 10536 14084 10592 14086
rect 10640 14138 10696 14140
rect 10640 14086 10642 14138
rect 10642 14086 10694 14138
rect 10694 14086 10696 14138
rect 10640 14084 10696 14086
rect 10744 14138 10800 14140
rect 10744 14086 10746 14138
rect 10746 14086 10798 14138
rect 10798 14086 10800 14138
rect 10744 14084 10800 14086
rect 2716 13858 2772 13860
rect 2716 13806 2718 13858
rect 2718 13806 2770 13858
rect 2770 13806 2772 13858
rect 2716 13804 2772 13806
rect 15708 13804 15764 13860
rect 15820 14252 15876 14308
rect 1708 13468 1764 13524
rect 2380 13356 2436 13412
rect 3612 13468 3668 13524
rect 3164 13356 3220 13412
rect 5874 13354 5930 13356
rect 5874 13302 5876 13354
rect 5876 13302 5928 13354
rect 5928 13302 5930 13354
rect 5874 13300 5930 13302
rect 5978 13354 6034 13356
rect 5978 13302 5980 13354
rect 5980 13302 6032 13354
rect 6032 13302 6034 13354
rect 5978 13300 6034 13302
rect 6082 13354 6138 13356
rect 6082 13302 6084 13354
rect 6084 13302 6136 13354
rect 6136 13302 6138 13354
rect 6082 13300 6138 13302
rect 15198 13354 15254 13356
rect 15198 13302 15200 13354
rect 15200 13302 15252 13354
rect 15252 13302 15254 13354
rect 15198 13300 15254 13302
rect 15302 13354 15358 13356
rect 15302 13302 15304 13354
rect 15304 13302 15356 13354
rect 15356 13302 15358 13354
rect 15302 13300 15358 13302
rect 15406 13354 15462 13356
rect 15406 13302 15408 13354
rect 15408 13302 15460 13354
rect 15460 13302 15462 13354
rect 15406 13300 15462 13302
rect 14700 13132 14756 13188
rect 4284 13020 4340 13076
rect 12684 12908 12740 12964
rect 2380 12796 2436 12852
rect 10536 12570 10592 12572
rect 10536 12518 10538 12570
rect 10538 12518 10590 12570
rect 10590 12518 10592 12570
rect 10536 12516 10592 12518
rect 10640 12570 10696 12572
rect 10640 12518 10642 12570
rect 10642 12518 10694 12570
rect 10694 12518 10696 12570
rect 10640 12516 10696 12518
rect 10744 12570 10800 12572
rect 10744 12518 10746 12570
rect 10746 12518 10798 12570
rect 10798 12518 10800 12570
rect 10744 12516 10800 12518
rect 1932 12124 1988 12180
rect 4284 12178 4340 12180
rect 4284 12126 4286 12178
rect 4286 12126 4338 12178
rect 4338 12126 4340 12178
rect 4284 12124 4340 12126
rect 5874 11786 5930 11788
rect 5874 11734 5876 11786
rect 5876 11734 5928 11786
rect 5928 11734 5930 11786
rect 5874 11732 5930 11734
rect 5978 11786 6034 11788
rect 5978 11734 5980 11786
rect 5980 11734 6032 11786
rect 6032 11734 6034 11786
rect 5978 11732 6034 11734
rect 6082 11786 6138 11788
rect 6082 11734 6084 11786
rect 6084 11734 6136 11786
rect 6136 11734 6138 11786
rect 6082 11732 6138 11734
rect 1932 11452 1988 11508
rect 10536 11002 10592 11004
rect 10536 10950 10538 11002
rect 10538 10950 10590 11002
rect 10590 10950 10592 11002
rect 10536 10948 10592 10950
rect 10640 11002 10696 11004
rect 10640 10950 10642 11002
rect 10642 10950 10694 11002
rect 10694 10950 10696 11002
rect 10640 10948 10696 10950
rect 10744 11002 10800 11004
rect 10744 10950 10746 11002
rect 10746 10950 10798 11002
rect 10798 10950 10800 11002
rect 10744 10948 10800 10950
rect 5874 10218 5930 10220
rect 5874 10166 5876 10218
rect 5876 10166 5928 10218
rect 5928 10166 5930 10218
rect 5874 10164 5930 10166
rect 5978 10218 6034 10220
rect 5978 10166 5980 10218
rect 5980 10166 6032 10218
rect 6032 10166 6034 10218
rect 5978 10164 6034 10166
rect 6082 10218 6138 10220
rect 6082 10166 6084 10218
rect 6084 10166 6136 10218
rect 6136 10166 6138 10218
rect 6082 10164 6138 10166
rect 10536 9434 10592 9436
rect 10536 9382 10538 9434
rect 10538 9382 10590 9434
rect 10590 9382 10592 9434
rect 10536 9380 10592 9382
rect 10640 9434 10696 9436
rect 10640 9382 10642 9434
rect 10642 9382 10694 9434
rect 10694 9382 10696 9434
rect 10640 9380 10696 9382
rect 10744 9434 10800 9436
rect 10744 9382 10746 9434
rect 10746 9382 10798 9434
rect 10798 9382 10800 9434
rect 10744 9380 10800 9382
rect 5874 8650 5930 8652
rect 5874 8598 5876 8650
rect 5876 8598 5928 8650
rect 5928 8598 5930 8650
rect 5874 8596 5930 8598
rect 5978 8650 6034 8652
rect 5978 8598 5980 8650
rect 5980 8598 6032 8650
rect 6032 8598 6034 8650
rect 5978 8596 6034 8598
rect 6082 8650 6138 8652
rect 6082 8598 6084 8650
rect 6084 8598 6136 8650
rect 6136 8598 6138 8650
rect 6082 8596 6138 8598
rect 10536 7866 10592 7868
rect 10536 7814 10538 7866
rect 10538 7814 10590 7866
rect 10590 7814 10592 7866
rect 10536 7812 10592 7814
rect 10640 7866 10696 7868
rect 10640 7814 10642 7866
rect 10642 7814 10694 7866
rect 10694 7814 10696 7866
rect 10640 7812 10696 7814
rect 10744 7866 10800 7868
rect 10744 7814 10746 7866
rect 10746 7814 10798 7866
rect 10798 7814 10800 7866
rect 10744 7812 10800 7814
rect 5874 7082 5930 7084
rect 5874 7030 5876 7082
rect 5876 7030 5928 7082
rect 5928 7030 5930 7082
rect 5874 7028 5930 7030
rect 5978 7082 6034 7084
rect 5978 7030 5980 7082
rect 5980 7030 6032 7082
rect 6032 7030 6034 7082
rect 5978 7028 6034 7030
rect 6082 7082 6138 7084
rect 6082 7030 6084 7082
rect 6084 7030 6136 7082
rect 6136 7030 6138 7082
rect 6082 7028 6138 7030
rect 10536 6298 10592 6300
rect 10536 6246 10538 6298
rect 10538 6246 10590 6298
rect 10590 6246 10592 6298
rect 10536 6244 10592 6246
rect 10640 6298 10696 6300
rect 10640 6246 10642 6298
rect 10642 6246 10694 6298
rect 10694 6246 10696 6298
rect 10640 6244 10696 6246
rect 10744 6298 10800 6300
rect 10744 6246 10746 6298
rect 10746 6246 10798 6298
rect 10798 6246 10800 6298
rect 10744 6244 10800 6246
rect 5874 5514 5930 5516
rect 5874 5462 5876 5514
rect 5876 5462 5928 5514
rect 5928 5462 5930 5514
rect 5874 5460 5930 5462
rect 5978 5514 6034 5516
rect 5978 5462 5980 5514
rect 5980 5462 6032 5514
rect 6032 5462 6034 5514
rect 5978 5460 6034 5462
rect 6082 5514 6138 5516
rect 6082 5462 6084 5514
rect 6084 5462 6136 5514
rect 6136 5462 6138 5514
rect 6082 5460 6138 5462
rect 10536 4730 10592 4732
rect 10536 4678 10538 4730
rect 10538 4678 10590 4730
rect 10590 4678 10592 4730
rect 10536 4676 10592 4678
rect 10640 4730 10696 4732
rect 10640 4678 10642 4730
rect 10642 4678 10694 4730
rect 10694 4678 10696 4730
rect 10640 4676 10696 4678
rect 10744 4730 10800 4732
rect 10744 4678 10746 4730
rect 10746 4678 10798 4730
rect 10798 4678 10800 4730
rect 10744 4676 10800 4678
rect 5874 3946 5930 3948
rect 5874 3894 5876 3946
rect 5876 3894 5928 3946
rect 5928 3894 5930 3946
rect 5874 3892 5930 3894
rect 5978 3946 6034 3948
rect 5978 3894 5980 3946
rect 5980 3894 6032 3946
rect 6032 3894 6034 3946
rect 5978 3892 6034 3894
rect 6082 3946 6138 3948
rect 6082 3894 6084 3946
rect 6084 3894 6136 3946
rect 6136 3894 6138 3946
rect 6082 3892 6138 3894
rect 12348 3388 12404 3444
rect 10536 3162 10592 3164
rect 10536 3110 10538 3162
rect 10538 3110 10590 3162
rect 10590 3110 10592 3162
rect 10536 3108 10592 3110
rect 10640 3162 10696 3164
rect 10640 3110 10642 3162
rect 10642 3110 10694 3162
rect 10694 3110 10696 3162
rect 10640 3108 10696 3110
rect 10744 3162 10800 3164
rect 10744 3110 10746 3162
rect 10746 3110 10798 3162
rect 10798 3110 10800 3162
rect 10744 3108 10800 3110
rect 14140 4898 14196 4900
rect 14140 4846 14142 4898
rect 14142 4846 14194 4898
rect 14194 4846 14196 4898
rect 14140 4844 14196 4846
rect 15198 11786 15254 11788
rect 15198 11734 15200 11786
rect 15200 11734 15252 11786
rect 15252 11734 15254 11786
rect 15198 11732 15254 11734
rect 15302 11786 15358 11788
rect 15302 11734 15304 11786
rect 15304 11734 15356 11786
rect 15356 11734 15358 11786
rect 15302 11732 15358 11734
rect 15406 11786 15462 11788
rect 15406 11734 15408 11786
rect 15408 11734 15460 11786
rect 15460 11734 15462 11786
rect 15406 11732 15462 11734
rect 15198 10218 15254 10220
rect 15198 10166 15200 10218
rect 15200 10166 15252 10218
rect 15252 10166 15254 10218
rect 15198 10164 15254 10166
rect 15302 10218 15358 10220
rect 15302 10166 15304 10218
rect 15304 10166 15356 10218
rect 15356 10166 15358 10218
rect 15302 10164 15358 10166
rect 15406 10218 15462 10220
rect 15406 10166 15408 10218
rect 15408 10166 15460 10218
rect 15460 10166 15462 10218
rect 15406 10164 15462 10166
rect 15596 10108 15652 10164
rect 15198 8650 15254 8652
rect 15198 8598 15200 8650
rect 15200 8598 15252 8650
rect 15252 8598 15254 8650
rect 15198 8596 15254 8598
rect 15302 8650 15358 8652
rect 15302 8598 15304 8650
rect 15304 8598 15356 8650
rect 15356 8598 15358 8650
rect 15302 8596 15358 8598
rect 15406 8650 15462 8652
rect 15406 8598 15408 8650
rect 15408 8598 15460 8650
rect 15460 8598 15462 8650
rect 15406 8596 15462 8598
rect 15198 7082 15254 7084
rect 15198 7030 15200 7082
rect 15200 7030 15252 7082
rect 15252 7030 15254 7082
rect 15198 7028 15254 7030
rect 15302 7082 15358 7084
rect 15302 7030 15304 7082
rect 15304 7030 15356 7082
rect 15356 7030 15358 7082
rect 15302 7028 15358 7030
rect 15406 7082 15462 7084
rect 15406 7030 15408 7082
rect 15408 7030 15460 7082
rect 15460 7030 15462 7082
rect 15406 7028 15462 7030
rect 15198 5514 15254 5516
rect 15198 5462 15200 5514
rect 15200 5462 15252 5514
rect 15252 5462 15254 5514
rect 15198 5460 15254 5462
rect 15302 5514 15358 5516
rect 15302 5462 15304 5514
rect 15304 5462 15356 5514
rect 15356 5462 15358 5514
rect 15302 5460 15358 5462
rect 15406 5514 15462 5516
rect 15406 5462 15408 5514
rect 15408 5462 15460 5514
rect 15460 5462 15462 5514
rect 15406 5460 15462 5462
rect 14812 5068 14868 5124
rect 13468 3388 13524 3444
rect 14924 4338 14980 4340
rect 14924 4286 14926 4338
rect 14926 4286 14978 4338
rect 14978 4286 14980 4338
rect 14924 4284 14980 4286
rect 15198 3946 15254 3948
rect 15198 3894 15200 3946
rect 15200 3894 15252 3946
rect 15252 3894 15254 3946
rect 15198 3892 15254 3894
rect 15302 3946 15358 3948
rect 15302 3894 15304 3946
rect 15304 3894 15356 3946
rect 15356 3894 15358 3946
rect 15302 3892 15358 3894
rect 15406 3946 15462 3948
rect 15406 3894 15408 3946
rect 15408 3894 15460 3946
rect 15460 3894 15462 3946
rect 15406 3892 15462 3894
rect 16828 18396 16884 18452
rect 17388 18338 17444 18340
rect 17388 18286 17390 18338
rect 17390 18286 17442 18338
rect 17442 18286 17444 18338
rect 17388 18284 17444 18286
rect 16268 17836 16324 17892
rect 16268 17388 16324 17444
rect 16044 15314 16100 15316
rect 16044 15262 16046 15314
rect 16046 15262 16098 15314
rect 16098 15262 16100 15314
rect 16044 15260 16100 15262
rect 19404 35308 19460 35364
rect 19516 27858 19572 27860
rect 19516 27806 19518 27858
rect 19518 27806 19570 27858
rect 19570 27806 19572 27858
rect 19516 27804 19572 27806
rect 19860 36090 19916 36092
rect 19860 36038 19862 36090
rect 19862 36038 19914 36090
rect 19914 36038 19916 36090
rect 19860 36036 19916 36038
rect 19964 36090 20020 36092
rect 19964 36038 19966 36090
rect 19966 36038 20018 36090
rect 20018 36038 20020 36090
rect 19964 36036 20020 36038
rect 20068 36090 20124 36092
rect 20068 36038 20070 36090
rect 20070 36038 20122 36090
rect 20122 36038 20124 36090
rect 20068 36036 20124 36038
rect 19860 34522 19916 34524
rect 19860 34470 19862 34522
rect 19862 34470 19914 34522
rect 19914 34470 19916 34522
rect 19860 34468 19916 34470
rect 19964 34522 20020 34524
rect 19964 34470 19966 34522
rect 19966 34470 20018 34522
rect 20018 34470 20020 34522
rect 19964 34468 20020 34470
rect 20068 34522 20124 34524
rect 20068 34470 20070 34522
rect 20070 34470 20122 34522
rect 20122 34470 20124 34522
rect 20068 34468 20124 34470
rect 19860 32954 19916 32956
rect 19860 32902 19862 32954
rect 19862 32902 19914 32954
rect 19914 32902 19916 32954
rect 19860 32900 19916 32902
rect 19964 32954 20020 32956
rect 19964 32902 19966 32954
rect 19966 32902 20018 32954
rect 20018 32902 20020 32954
rect 19964 32900 20020 32902
rect 20068 32954 20124 32956
rect 20068 32902 20070 32954
rect 20070 32902 20122 32954
rect 20122 32902 20124 32954
rect 20068 32900 20124 32902
rect 19860 31386 19916 31388
rect 19860 31334 19862 31386
rect 19862 31334 19914 31386
rect 19914 31334 19916 31386
rect 19860 31332 19916 31334
rect 19964 31386 20020 31388
rect 19964 31334 19966 31386
rect 19966 31334 20018 31386
rect 20018 31334 20020 31386
rect 19964 31332 20020 31334
rect 20068 31386 20124 31388
rect 20068 31334 20070 31386
rect 20070 31334 20122 31386
rect 20122 31334 20124 31386
rect 20068 31332 20124 31334
rect 19860 29818 19916 29820
rect 19860 29766 19862 29818
rect 19862 29766 19914 29818
rect 19914 29766 19916 29818
rect 19860 29764 19916 29766
rect 19964 29818 20020 29820
rect 19964 29766 19966 29818
rect 19966 29766 20018 29818
rect 20018 29766 20020 29818
rect 19964 29764 20020 29766
rect 20068 29818 20124 29820
rect 20068 29766 20070 29818
rect 20070 29766 20122 29818
rect 20122 29766 20124 29818
rect 20068 29764 20124 29766
rect 19860 28250 19916 28252
rect 19860 28198 19862 28250
rect 19862 28198 19914 28250
rect 19914 28198 19916 28250
rect 19860 28196 19916 28198
rect 19964 28250 20020 28252
rect 19964 28198 19966 28250
rect 19966 28198 20018 28250
rect 20018 28198 20020 28250
rect 19964 28196 20020 28198
rect 20068 28250 20124 28252
rect 20068 28198 20070 28250
rect 20070 28198 20122 28250
rect 20122 28198 20124 28250
rect 20068 28196 20124 28198
rect 20636 31948 20692 32004
rect 20412 27244 20468 27300
rect 20300 26908 20356 26964
rect 19860 26682 19916 26684
rect 19860 26630 19862 26682
rect 19862 26630 19914 26682
rect 19914 26630 19916 26682
rect 19860 26628 19916 26630
rect 19964 26682 20020 26684
rect 19964 26630 19966 26682
rect 19966 26630 20018 26682
rect 20018 26630 20020 26682
rect 19964 26628 20020 26630
rect 20068 26682 20124 26684
rect 20068 26630 20070 26682
rect 20070 26630 20122 26682
rect 20122 26630 20124 26682
rect 20068 26628 20124 26630
rect 20188 25228 20244 25284
rect 19860 25114 19916 25116
rect 19860 25062 19862 25114
rect 19862 25062 19914 25114
rect 19914 25062 19916 25114
rect 19860 25060 19916 25062
rect 19964 25114 20020 25116
rect 19964 25062 19966 25114
rect 19966 25062 20018 25114
rect 20018 25062 20020 25114
rect 19964 25060 20020 25062
rect 20068 25114 20124 25116
rect 20068 25062 20070 25114
rect 20070 25062 20122 25114
rect 20122 25062 20124 25114
rect 20068 25060 20124 25062
rect 19740 24668 19796 24724
rect 20300 24722 20356 24724
rect 20300 24670 20302 24722
rect 20302 24670 20354 24722
rect 20354 24670 20356 24722
rect 20300 24668 20356 24670
rect 19860 23546 19916 23548
rect 19860 23494 19862 23546
rect 19862 23494 19914 23546
rect 19914 23494 19916 23546
rect 19860 23492 19916 23494
rect 19964 23546 20020 23548
rect 19964 23494 19966 23546
rect 19966 23494 20018 23546
rect 20018 23494 20020 23546
rect 19964 23492 20020 23494
rect 20068 23546 20124 23548
rect 20068 23494 20070 23546
rect 20070 23494 20122 23546
rect 20122 23494 20124 23546
rect 20068 23492 20124 23494
rect 20188 23212 20244 23268
rect 19068 22428 19124 22484
rect 18508 21644 18564 21700
rect 17948 21474 18004 21476
rect 17948 21422 17950 21474
rect 17950 21422 18002 21474
rect 18002 21422 18004 21474
rect 17948 21420 18004 21422
rect 18508 20972 18564 21028
rect 18956 21420 19012 21476
rect 18284 20690 18340 20692
rect 18284 20638 18286 20690
rect 18286 20638 18338 20690
rect 18338 20638 18340 20690
rect 18284 20636 18340 20638
rect 18620 20578 18676 20580
rect 18620 20526 18622 20578
rect 18622 20526 18674 20578
rect 18674 20526 18676 20578
rect 18620 20524 18676 20526
rect 18508 19122 18564 19124
rect 18508 19070 18510 19122
rect 18510 19070 18562 19122
rect 18562 19070 18564 19122
rect 18508 19068 18564 19070
rect 18732 19180 18788 19236
rect 17948 16716 18004 16772
rect 18060 17052 18116 17108
rect 17388 16098 17444 16100
rect 17388 16046 17390 16098
rect 17390 16046 17442 16098
rect 17442 16046 17444 16098
rect 17388 16044 17444 16046
rect 17948 16098 18004 16100
rect 17948 16046 17950 16098
rect 17950 16046 18002 16098
rect 18002 16046 18004 16098
rect 17948 16044 18004 16046
rect 18284 16044 18340 16100
rect 18508 17500 18564 17556
rect 18620 18508 18676 18564
rect 18508 16940 18564 16996
rect 18732 16380 18788 16436
rect 19628 22428 19684 22484
rect 19516 22092 19572 22148
rect 19860 21978 19916 21980
rect 19860 21926 19862 21978
rect 19862 21926 19914 21978
rect 19914 21926 19916 21978
rect 19860 21924 19916 21926
rect 19964 21978 20020 21980
rect 19964 21926 19966 21978
rect 19966 21926 20018 21978
rect 20018 21926 20020 21978
rect 19964 21924 20020 21926
rect 20068 21978 20124 21980
rect 20068 21926 20070 21978
rect 20070 21926 20122 21978
rect 20122 21926 20124 21978
rect 20068 21924 20124 21926
rect 20076 21420 20132 21476
rect 20412 21698 20468 21700
rect 20412 21646 20414 21698
rect 20414 21646 20466 21698
rect 20466 21646 20468 21698
rect 20412 21644 20468 21646
rect 20636 26124 20692 26180
rect 20636 22146 20692 22148
rect 20636 22094 20638 22146
rect 20638 22094 20690 22146
rect 20690 22094 20692 22146
rect 20636 22092 20692 22094
rect 20300 21474 20356 21476
rect 20300 21422 20302 21474
rect 20302 21422 20354 21474
rect 20354 21422 20356 21474
rect 20300 21420 20356 21422
rect 20188 20802 20244 20804
rect 20188 20750 20190 20802
rect 20190 20750 20242 20802
rect 20242 20750 20244 20802
rect 20188 20748 20244 20750
rect 20860 35308 20916 35364
rect 22092 36706 22148 36708
rect 22092 36654 22094 36706
rect 22094 36654 22146 36706
rect 22146 36654 22148 36706
rect 22092 36652 22148 36654
rect 24220 36764 24276 36820
rect 24522 36874 24578 36876
rect 24522 36822 24524 36874
rect 24524 36822 24576 36874
rect 24576 36822 24578 36874
rect 24522 36820 24578 36822
rect 24626 36874 24682 36876
rect 24626 36822 24628 36874
rect 24628 36822 24680 36874
rect 24680 36822 24682 36874
rect 24626 36820 24682 36822
rect 24730 36874 24786 36876
rect 24730 36822 24732 36874
rect 24732 36822 24784 36874
rect 24784 36822 24786 36874
rect 24730 36820 24786 36822
rect 26236 36876 26292 36932
rect 27468 36876 27524 36932
rect 22876 36428 22932 36484
rect 22204 35756 22260 35812
rect 23100 35756 23156 35812
rect 22764 35644 22820 35700
rect 22652 34860 22708 34916
rect 21868 32284 21924 32340
rect 21084 27244 21140 27300
rect 20972 26290 21028 26292
rect 20972 26238 20974 26290
rect 20974 26238 21026 26290
rect 21026 26238 21028 26290
rect 20972 26236 21028 26238
rect 20972 24722 21028 24724
rect 20972 24670 20974 24722
rect 20974 24670 21026 24722
rect 21026 24670 21028 24722
rect 20972 24668 21028 24670
rect 21308 26962 21364 26964
rect 21308 26910 21310 26962
rect 21310 26910 21362 26962
rect 21362 26910 21364 26962
rect 21308 26908 21364 26910
rect 21420 26178 21476 26180
rect 21420 26126 21422 26178
rect 21422 26126 21474 26178
rect 21474 26126 21476 26178
rect 21420 26124 21476 26126
rect 21196 25282 21252 25284
rect 21196 25230 21198 25282
rect 21198 25230 21250 25282
rect 21250 25230 21252 25282
rect 21196 25228 21252 25230
rect 21532 25394 21588 25396
rect 21532 25342 21534 25394
rect 21534 25342 21586 25394
rect 21586 25342 21588 25394
rect 21532 25340 21588 25342
rect 21644 25228 21700 25284
rect 21756 26124 21812 26180
rect 21308 24892 21364 24948
rect 22092 31948 22148 32004
rect 22204 31500 22260 31556
rect 21532 23324 21588 23380
rect 21756 23212 21812 23268
rect 20860 22092 20916 22148
rect 19860 20410 19916 20412
rect 19860 20358 19862 20410
rect 19862 20358 19914 20410
rect 19914 20358 19916 20410
rect 19860 20356 19916 20358
rect 19964 20410 20020 20412
rect 19964 20358 19966 20410
rect 19966 20358 20018 20410
rect 20018 20358 20020 20410
rect 19964 20356 20020 20358
rect 20068 20410 20124 20412
rect 20068 20358 20070 20410
rect 20070 20358 20122 20410
rect 20122 20358 20124 20410
rect 20068 20356 20124 20358
rect 19292 19404 19348 19460
rect 19740 20076 19796 20132
rect 19964 20188 20020 20244
rect 19628 19234 19684 19236
rect 19628 19182 19630 19234
rect 19630 19182 19682 19234
rect 19682 19182 19684 19234
rect 19628 19180 19684 19182
rect 20300 20076 20356 20132
rect 20412 19292 20468 19348
rect 19180 18620 19236 18676
rect 19860 18842 19916 18844
rect 19860 18790 19862 18842
rect 19862 18790 19914 18842
rect 19914 18790 19916 18842
rect 19860 18788 19916 18790
rect 19964 18842 20020 18844
rect 19964 18790 19966 18842
rect 19966 18790 20018 18842
rect 20018 18790 20020 18842
rect 19964 18788 20020 18790
rect 20068 18842 20124 18844
rect 20068 18790 20070 18842
rect 20070 18790 20122 18842
rect 20122 18790 20124 18842
rect 20068 18788 20124 18790
rect 18956 18450 19012 18452
rect 18956 18398 18958 18450
rect 18958 18398 19010 18450
rect 19010 18398 19012 18450
rect 18956 18396 19012 18398
rect 19292 18172 19348 18228
rect 19740 18508 19796 18564
rect 21196 20748 21252 20804
rect 21532 22092 21588 22148
rect 20972 20188 21028 20244
rect 21420 20636 21476 20692
rect 20860 19292 20916 19348
rect 20412 18450 20468 18452
rect 20412 18398 20414 18450
rect 20414 18398 20466 18450
rect 20466 18398 20468 18450
rect 20412 18396 20468 18398
rect 21084 19180 21140 19236
rect 21756 20132 21812 20188
rect 21532 19740 21588 19796
rect 21644 20018 21700 20020
rect 21644 19966 21646 20018
rect 21646 19966 21698 20018
rect 21698 19966 21700 20018
rect 21644 19964 21700 19966
rect 22540 25228 22596 25284
rect 22652 24834 22708 24836
rect 22652 24782 22654 24834
rect 22654 24782 22706 24834
rect 22706 24782 22708 24834
rect 22652 24780 22708 24782
rect 23548 35756 23604 35812
rect 23996 35810 24052 35812
rect 23996 35758 23998 35810
rect 23998 35758 24050 35810
rect 24050 35758 24052 35810
rect 23996 35756 24052 35758
rect 24892 36540 24948 36596
rect 25452 36652 25508 36708
rect 24780 36482 24836 36484
rect 24780 36430 24782 36482
rect 24782 36430 24834 36482
rect 24834 36430 24836 36482
rect 24780 36428 24836 36430
rect 24220 35420 24276 35476
rect 23324 31500 23380 31556
rect 23996 33404 24052 33460
rect 22876 25394 22932 25396
rect 22876 25342 22878 25394
rect 22878 25342 22930 25394
rect 22930 25342 22932 25394
rect 22876 25340 22932 25342
rect 22876 24946 22932 24948
rect 22876 24894 22878 24946
rect 22878 24894 22930 24946
rect 22930 24894 22932 24946
rect 22876 24892 22932 24894
rect 22988 24834 23044 24836
rect 22988 24782 22990 24834
rect 22990 24782 23042 24834
rect 23042 24782 23044 24834
rect 22988 24780 23044 24782
rect 25004 36204 25060 36260
rect 24522 35306 24578 35308
rect 24522 35254 24524 35306
rect 24524 35254 24576 35306
rect 24576 35254 24578 35306
rect 24522 35252 24578 35254
rect 24626 35306 24682 35308
rect 24626 35254 24628 35306
rect 24628 35254 24680 35306
rect 24680 35254 24682 35306
rect 24626 35252 24682 35254
rect 24730 35306 24786 35308
rect 24730 35254 24732 35306
rect 24732 35254 24784 35306
rect 24784 35254 24786 35306
rect 24730 35252 24786 35254
rect 24332 34860 24388 34916
rect 24522 33738 24578 33740
rect 24522 33686 24524 33738
rect 24524 33686 24576 33738
rect 24576 33686 24578 33738
rect 24522 33684 24578 33686
rect 24626 33738 24682 33740
rect 24626 33686 24628 33738
rect 24628 33686 24680 33738
rect 24680 33686 24682 33738
rect 24626 33684 24682 33686
rect 24730 33738 24786 33740
rect 24730 33686 24732 33738
rect 24732 33686 24784 33738
rect 24784 33686 24786 33738
rect 24730 33684 24786 33686
rect 24892 33516 24948 33572
rect 24522 32170 24578 32172
rect 24522 32118 24524 32170
rect 24524 32118 24576 32170
rect 24576 32118 24578 32170
rect 24522 32116 24578 32118
rect 24626 32170 24682 32172
rect 24626 32118 24628 32170
rect 24628 32118 24680 32170
rect 24680 32118 24682 32170
rect 24626 32116 24682 32118
rect 24730 32170 24786 32172
rect 24730 32118 24732 32170
rect 24732 32118 24784 32170
rect 24784 32118 24786 32170
rect 24730 32116 24786 32118
rect 24522 30602 24578 30604
rect 24522 30550 24524 30602
rect 24524 30550 24576 30602
rect 24576 30550 24578 30602
rect 24522 30548 24578 30550
rect 24626 30602 24682 30604
rect 24626 30550 24628 30602
rect 24628 30550 24680 30602
rect 24680 30550 24682 30602
rect 24626 30548 24682 30550
rect 24730 30602 24786 30604
rect 24730 30550 24732 30602
rect 24732 30550 24784 30602
rect 24784 30550 24786 30602
rect 24730 30548 24786 30550
rect 24522 29034 24578 29036
rect 24522 28982 24524 29034
rect 24524 28982 24576 29034
rect 24576 28982 24578 29034
rect 24522 28980 24578 28982
rect 24626 29034 24682 29036
rect 24626 28982 24628 29034
rect 24628 28982 24680 29034
rect 24680 28982 24682 29034
rect 24626 28980 24682 28982
rect 24730 29034 24786 29036
rect 24730 28982 24732 29034
rect 24732 28982 24784 29034
rect 24784 28982 24786 29034
rect 24730 28980 24786 28982
rect 24522 27466 24578 27468
rect 24522 27414 24524 27466
rect 24524 27414 24576 27466
rect 24576 27414 24578 27466
rect 24522 27412 24578 27414
rect 24626 27466 24682 27468
rect 24626 27414 24628 27466
rect 24628 27414 24680 27466
rect 24680 27414 24682 27466
rect 24626 27412 24682 27414
rect 24730 27466 24786 27468
rect 24730 27414 24732 27466
rect 24732 27414 24784 27466
rect 24784 27414 24786 27466
rect 24730 27412 24786 27414
rect 24522 25898 24578 25900
rect 24522 25846 24524 25898
rect 24524 25846 24576 25898
rect 24576 25846 24578 25898
rect 24522 25844 24578 25846
rect 24626 25898 24682 25900
rect 24626 25846 24628 25898
rect 24628 25846 24680 25898
rect 24680 25846 24682 25898
rect 24626 25844 24682 25846
rect 24730 25898 24786 25900
rect 24730 25846 24732 25898
rect 24732 25846 24784 25898
rect 24784 25846 24786 25898
rect 24730 25844 24786 25846
rect 24522 24330 24578 24332
rect 24522 24278 24524 24330
rect 24524 24278 24576 24330
rect 24576 24278 24578 24330
rect 24522 24276 24578 24278
rect 24626 24330 24682 24332
rect 24626 24278 24628 24330
rect 24628 24278 24680 24330
rect 24680 24278 24682 24330
rect 24626 24276 24682 24278
rect 24730 24330 24786 24332
rect 24730 24278 24732 24330
rect 24732 24278 24784 24330
rect 24784 24278 24786 24330
rect 24730 24276 24786 24278
rect 26236 36482 26292 36484
rect 26236 36430 26238 36482
rect 26238 36430 26290 36482
rect 26290 36430 26292 36482
rect 26236 36428 26292 36430
rect 25228 35420 25284 35476
rect 26572 36258 26628 36260
rect 26572 36206 26574 36258
rect 26574 36206 26626 36258
rect 26626 36206 26628 36258
rect 26572 36204 26628 36206
rect 28476 36876 28532 36932
rect 33846 36874 33902 36876
rect 33846 36822 33848 36874
rect 33848 36822 33900 36874
rect 33900 36822 33902 36874
rect 33846 36820 33902 36822
rect 33950 36874 34006 36876
rect 33950 36822 33952 36874
rect 33952 36822 34004 36874
rect 34004 36822 34006 36874
rect 33950 36820 34006 36822
rect 34054 36874 34110 36876
rect 34054 36822 34056 36874
rect 34056 36822 34108 36874
rect 34108 36822 34110 36874
rect 34054 36820 34110 36822
rect 29184 36090 29240 36092
rect 29184 36038 29186 36090
rect 29186 36038 29238 36090
rect 29238 36038 29240 36090
rect 29184 36036 29240 36038
rect 29288 36090 29344 36092
rect 29288 36038 29290 36090
rect 29290 36038 29342 36090
rect 29342 36038 29344 36090
rect 29288 36036 29344 36038
rect 29392 36090 29448 36092
rect 29392 36038 29394 36090
rect 29394 36038 29446 36090
rect 29446 36038 29448 36090
rect 29392 36036 29448 36038
rect 38508 36090 38564 36092
rect 38508 36038 38510 36090
rect 38510 36038 38562 36090
rect 38562 36038 38564 36090
rect 38508 36036 38564 36038
rect 38612 36090 38668 36092
rect 38612 36038 38614 36090
rect 38614 36038 38666 36090
rect 38666 36038 38668 36090
rect 38612 36036 38668 36038
rect 38716 36090 38772 36092
rect 38716 36038 38718 36090
rect 38718 36038 38770 36090
rect 38770 36038 38772 36090
rect 38716 36036 38772 36038
rect 33846 35306 33902 35308
rect 33846 35254 33848 35306
rect 33848 35254 33900 35306
rect 33900 35254 33902 35306
rect 33846 35252 33902 35254
rect 33950 35306 34006 35308
rect 33950 35254 33952 35306
rect 33952 35254 34004 35306
rect 34004 35254 34006 35306
rect 33950 35252 34006 35254
rect 34054 35306 34110 35308
rect 34054 35254 34056 35306
rect 34056 35254 34108 35306
rect 34108 35254 34110 35306
rect 34054 35252 34110 35254
rect 29184 34522 29240 34524
rect 29184 34470 29186 34522
rect 29186 34470 29238 34522
rect 29238 34470 29240 34522
rect 29184 34468 29240 34470
rect 29288 34522 29344 34524
rect 29288 34470 29290 34522
rect 29290 34470 29342 34522
rect 29342 34470 29344 34522
rect 29288 34468 29344 34470
rect 29392 34522 29448 34524
rect 29392 34470 29394 34522
rect 29394 34470 29446 34522
rect 29446 34470 29448 34522
rect 29392 34468 29448 34470
rect 38508 34522 38564 34524
rect 38508 34470 38510 34522
rect 38510 34470 38562 34522
rect 38562 34470 38564 34522
rect 38508 34468 38564 34470
rect 38612 34522 38668 34524
rect 38612 34470 38614 34522
rect 38614 34470 38666 34522
rect 38666 34470 38668 34522
rect 38612 34468 38668 34470
rect 38716 34522 38772 34524
rect 38716 34470 38718 34522
rect 38718 34470 38770 34522
rect 38770 34470 38772 34522
rect 38716 34468 38772 34470
rect 33846 33738 33902 33740
rect 33846 33686 33848 33738
rect 33848 33686 33900 33738
rect 33900 33686 33902 33738
rect 33846 33684 33902 33686
rect 33950 33738 34006 33740
rect 33950 33686 33952 33738
rect 33952 33686 34004 33738
rect 34004 33686 34006 33738
rect 33950 33684 34006 33686
rect 34054 33738 34110 33740
rect 34054 33686 34056 33738
rect 34056 33686 34108 33738
rect 34108 33686 34110 33738
rect 34054 33684 34110 33686
rect 27468 33516 27524 33572
rect 27132 33404 27188 33460
rect 29184 32954 29240 32956
rect 29184 32902 29186 32954
rect 29186 32902 29238 32954
rect 29238 32902 29240 32954
rect 29184 32900 29240 32902
rect 29288 32954 29344 32956
rect 29288 32902 29290 32954
rect 29290 32902 29342 32954
rect 29342 32902 29344 32954
rect 29288 32900 29344 32902
rect 29392 32954 29448 32956
rect 29392 32902 29394 32954
rect 29394 32902 29446 32954
rect 29446 32902 29448 32954
rect 29392 32900 29448 32902
rect 38508 32954 38564 32956
rect 38508 32902 38510 32954
rect 38510 32902 38562 32954
rect 38562 32902 38564 32954
rect 38508 32900 38564 32902
rect 38612 32954 38668 32956
rect 38612 32902 38614 32954
rect 38614 32902 38666 32954
rect 38666 32902 38668 32954
rect 38612 32900 38668 32902
rect 38716 32954 38772 32956
rect 38716 32902 38718 32954
rect 38718 32902 38770 32954
rect 38770 32902 38772 32954
rect 38716 32900 38772 32902
rect 25788 32284 25844 32340
rect 33846 32170 33902 32172
rect 33846 32118 33848 32170
rect 33848 32118 33900 32170
rect 33900 32118 33902 32170
rect 33846 32116 33902 32118
rect 33950 32170 34006 32172
rect 33950 32118 33952 32170
rect 33952 32118 34004 32170
rect 34004 32118 34006 32170
rect 33950 32116 34006 32118
rect 34054 32170 34110 32172
rect 34054 32118 34056 32170
rect 34056 32118 34108 32170
rect 34108 32118 34110 32170
rect 34054 32116 34110 32118
rect 29184 31386 29240 31388
rect 29184 31334 29186 31386
rect 29186 31334 29238 31386
rect 29238 31334 29240 31386
rect 29184 31332 29240 31334
rect 29288 31386 29344 31388
rect 29288 31334 29290 31386
rect 29290 31334 29342 31386
rect 29342 31334 29344 31386
rect 29288 31332 29344 31334
rect 29392 31386 29448 31388
rect 29392 31334 29394 31386
rect 29394 31334 29446 31386
rect 29446 31334 29448 31386
rect 29392 31332 29448 31334
rect 38508 31386 38564 31388
rect 38508 31334 38510 31386
rect 38510 31334 38562 31386
rect 38562 31334 38564 31386
rect 38508 31332 38564 31334
rect 38612 31386 38668 31388
rect 38612 31334 38614 31386
rect 38614 31334 38666 31386
rect 38666 31334 38668 31386
rect 38612 31332 38668 31334
rect 38716 31386 38772 31388
rect 38716 31334 38718 31386
rect 38718 31334 38770 31386
rect 38770 31334 38772 31386
rect 38716 31332 38772 31334
rect 33846 30602 33902 30604
rect 33846 30550 33848 30602
rect 33848 30550 33900 30602
rect 33900 30550 33902 30602
rect 33846 30548 33902 30550
rect 33950 30602 34006 30604
rect 33950 30550 33952 30602
rect 33952 30550 34004 30602
rect 34004 30550 34006 30602
rect 33950 30548 34006 30550
rect 34054 30602 34110 30604
rect 34054 30550 34056 30602
rect 34056 30550 34108 30602
rect 34108 30550 34110 30602
rect 34054 30548 34110 30550
rect 29184 29818 29240 29820
rect 29184 29766 29186 29818
rect 29186 29766 29238 29818
rect 29238 29766 29240 29818
rect 29184 29764 29240 29766
rect 29288 29818 29344 29820
rect 29288 29766 29290 29818
rect 29290 29766 29342 29818
rect 29342 29766 29344 29818
rect 29288 29764 29344 29766
rect 29392 29818 29448 29820
rect 29392 29766 29394 29818
rect 29394 29766 29446 29818
rect 29446 29766 29448 29818
rect 29392 29764 29448 29766
rect 33846 29034 33902 29036
rect 33846 28982 33848 29034
rect 33848 28982 33900 29034
rect 33900 28982 33902 29034
rect 33846 28980 33902 28982
rect 33950 29034 34006 29036
rect 33950 28982 33952 29034
rect 33952 28982 34004 29034
rect 34004 28982 34006 29034
rect 33950 28980 34006 28982
rect 34054 29034 34110 29036
rect 34054 28982 34056 29034
rect 34056 28982 34108 29034
rect 34108 28982 34110 29034
rect 34054 28980 34110 28982
rect 28700 28700 28756 28756
rect 26460 25228 26516 25284
rect 25564 24610 25620 24612
rect 25564 24558 25566 24610
rect 25566 24558 25618 24610
rect 25618 24558 25620 24610
rect 25564 24556 25620 24558
rect 23548 23266 23604 23268
rect 23548 23214 23550 23266
rect 23550 23214 23602 23266
rect 23602 23214 23604 23266
rect 23548 23212 23604 23214
rect 21980 22258 22036 22260
rect 21980 22206 21982 22258
rect 21982 22206 22034 22258
rect 22034 22206 22036 22258
rect 21980 22204 22036 22206
rect 22204 22146 22260 22148
rect 22204 22094 22206 22146
rect 22206 22094 22258 22146
rect 22258 22094 22260 22146
rect 22204 22092 22260 22094
rect 21868 19852 21924 19908
rect 22764 20300 22820 20356
rect 23212 21474 23268 21476
rect 23212 21422 23214 21474
rect 23214 21422 23266 21474
rect 23266 21422 23268 21474
rect 23212 21420 23268 21422
rect 23100 20690 23156 20692
rect 23100 20638 23102 20690
rect 23102 20638 23154 20690
rect 23154 20638 23156 20690
rect 23100 20636 23156 20638
rect 25452 23042 25508 23044
rect 25452 22990 25454 23042
rect 25454 22990 25506 23042
rect 25506 22990 25508 23042
rect 25452 22988 25508 22990
rect 24522 22762 24578 22764
rect 24522 22710 24524 22762
rect 24524 22710 24576 22762
rect 24576 22710 24578 22762
rect 24522 22708 24578 22710
rect 24626 22762 24682 22764
rect 24626 22710 24628 22762
rect 24628 22710 24680 22762
rect 24680 22710 24682 22762
rect 24626 22708 24682 22710
rect 24730 22762 24786 22764
rect 24730 22710 24732 22762
rect 24732 22710 24784 22762
rect 24784 22710 24786 22762
rect 24730 22708 24786 22710
rect 23436 21420 23492 21476
rect 23772 21420 23828 21476
rect 23772 20972 23828 21028
rect 23436 20636 23492 20692
rect 24444 21474 24500 21476
rect 24444 21422 24446 21474
rect 24446 21422 24498 21474
rect 24498 21422 24500 21474
rect 24444 21420 24500 21422
rect 25004 21420 25060 21476
rect 23996 20524 24052 20580
rect 22876 20076 22932 20132
rect 23212 20130 23268 20132
rect 23212 20078 23214 20130
rect 23214 20078 23266 20130
rect 23266 20078 23268 20130
rect 23212 20076 23268 20078
rect 21644 19516 21700 19572
rect 21532 18450 21588 18452
rect 21532 18398 21534 18450
rect 21534 18398 21586 18450
rect 21586 18398 21588 18450
rect 21532 18396 21588 18398
rect 19068 17554 19124 17556
rect 19068 17502 19070 17554
rect 19070 17502 19122 17554
rect 19122 17502 19124 17554
rect 19068 17500 19124 17502
rect 19628 17836 19684 17892
rect 19964 17666 20020 17668
rect 19964 17614 19966 17666
rect 19966 17614 20018 17666
rect 20018 17614 20020 17666
rect 19964 17612 20020 17614
rect 19852 17554 19908 17556
rect 19852 17502 19854 17554
rect 19854 17502 19906 17554
rect 19906 17502 19908 17554
rect 19852 17500 19908 17502
rect 20412 17554 20468 17556
rect 20412 17502 20414 17554
rect 20414 17502 20466 17554
rect 20466 17502 20468 17554
rect 20412 17500 20468 17502
rect 20188 17442 20244 17444
rect 20188 17390 20190 17442
rect 20190 17390 20242 17442
rect 20242 17390 20244 17442
rect 20188 17388 20244 17390
rect 19860 17274 19916 17276
rect 19860 17222 19862 17274
rect 19862 17222 19914 17274
rect 19914 17222 19916 17274
rect 19860 17220 19916 17222
rect 19964 17274 20020 17276
rect 19964 17222 19966 17274
rect 19966 17222 20018 17274
rect 20018 17222 20020 17274
rect 19964 17220 20020 17222
rect 20068 17274 20124 17276
rect 20068 17222 20070 17274
rect 20070 17222 20122 17274
rect 20122 17222 20124 17274
rect 20068 17220 20124 17222
rect 20524 17164 20580 17220
rect 19740 17106 19796 17108
rect 19740 17054 19742 17106
rect 19742 17054 19794 17106
rect 19794 17054 19796 17106
rect 19740 17052 19796 17054
rect 20412 17106 20468 17108
rect 20412 17054 20414 17106
rect 20414 17054 20466 17106
rect 20466 17054 20468 17106
rect 20412 17052 20468 17054
rect 19180 16828 19236 16884
rect 19964 16882 20020 16884
rect 19964 16830 19966 16882
rect 19966 16830 20018 16882
rect 20018 16830 20020 16882
rect 19964 16828 20020 16830
rect 18956 16770 19012 16772
rect 18956 16718 18958 16770
rect 18958 16718 19010 16770
rect 19010 16718 19012 16770
rect 18956 16716 19012 16718
rect 19292 16770 19348 16772
rect 19292 16718 19294 16770
rect 19294 16718 19346 16770
rect 19346 16718 19348 16770
rect 19292 16716 19348 16718
rect 19068 16380 19124 16436
rect 18060 15260 18116 15316
rect 18620 15314 18676 15316
rect 18620 15262 18622 15314
rect 18622 15262 18674 15314
rect 18674 15262 18676 15314
rect 18620 15260 18676 15262
rect 18060 14476 18116 14532
rect 17948 13970 18004 13972
rect 17948 13918 17950 13970
rect 17950 13918 18002 13970
rect 18002 13918 18004 13970
rect 17948 13916 18004 13918
rect 16828 13020 16884 13076
rect 18284 13634 18340 13636
rect 18284 13582 18286 13634
rect 18286 13582 18338 13634
rect 18338 13582 18340 13634
rect 18284 13580 18340 13582
rect 17836 12796 17892 12852
rect 15932 12124 15988 12180
rect 18060 11788 18116 11844
rect 16044 4562 16100 4564
rect 16044 4510 16046 4562
rect 16046 4510 16098 4562
rect 16098 4510 16100 4562
rect 16044 4508 16100 4510
rect 16380 4620 16436 4676
rect 17388 3442 17444 3444
rect 17388 3390 17390 3442
rect 17390 3390 17442 3442
rect 17442 3390 17444 3442
rect 17388 3388 17444 3390
rect 18172 3500 18228 3556
rect 18620 14924 18676 14980
rect 18508 13522 18564 13524
rect 18508 13470 18510 13522
rect 18510 13470 18562 13522
rect 18562 13470 18564 13522
rect 18508 13468 18564 13470
rect 18956 15820 19012 15876
rect 19516 16380 19572 16436
rect 19740 16044 19796 16100
rect 19180 15260 19236 15316
rect 19292 14924 19348 14980
rect 19516 15820 19572 15876
rect 19404 14812 19460 14868
rect 19628 14364 19684 14420
rect 19860 15706 19916 15708
rect 19860 15654 19862 15706
rect 19862 15654 19914 15706
rect 19914 15654 19916 15706
rect 19860 15652 19916 15654
rect 19964 15706 20020 15708
rect 19964 15654 19966 15706
rect 19966 15654 20018 15706
rect 20018 15654 20020 15706
rect 19964 15652 20020 15654
rect 20068 15706 20124 15708
rect 20068 15654 20070 15706
rect 20070 15654 20122 15706
rect 20122 15654 20124 15706
rect 20068 15652 20124 15654
rect 20076 15314 20132 15316
rect 20076 15262 20078 15314
rect 20078 15262 20130 15314
rect 20130 15262 20132 15314
rect 20076 15260 20132 15262
rect 20188 15202 20244 15204
rect 20188 15150 20190 15202
rect 20190 15150 20242 15202
rect 20242 15150 20244 15202
rect 20188 15148 20244 15150
rect 20188 14588 20244 14644
rect 19964 14418 20020 14420
rect 19964 14366 19966 14418
rect 19966 14366 20018 14418
rect 20018 14366 20020 14418
rect 19964 14364 20020 14366
rect 19860 14138 19916 14140
rect 19860 14086 19862 14138
rect 19862 14086 19914 14138
rect 19914 14086 19916 14138
rect 19860 14084 19916 14086
rect 19964 14138 20020 14140
rect 19964 14086 19966 14138
rect 19966 14086 20018 14138
rect 20018 14086 20020 14138
rect 19964 14084 20020 14086
rect 20068 14138 20124 14140
rect 20068 14086 20070 14138
rect 20070 14086 20122 14138
rect 20122 14086 20124 14138
rect 20068 14084 20124 14086
rect 18956 13634 19012 13636
rect 18956 13582 18958 13634
rect 18958 13582 19010 13634
rect 19010 13582 19012 13634
rect 18956 13580 19012 13582
rect 19292 13132 19348 13188
rect 19292 12962 19348 12964
rect 19292 12910 19294 12962
rect 19294 12910 19346 12962
rect 19346 12910 19348 12962
rect 19292 12908 19348 12910
rect 21868 19516 21924 19572
rect 22764 20018 22820 20020
rect 22764 19966 22766 20018
rect 22766 19966 22818 20018
rect 22818 19966 22820 20018
rect 22764 19964 22820 19966
rect 22092 19516 22148 19572
rect 23324 19852 23380 19908
rect 23212 18620 23268 18676
rect 23548 19740 23604 19796
rect 22876 18450 22932 18452
rect 22876 18398 22878 18450
rect 22878 18398 22930 18450
rect 22930 18398 22932 18450
rect 22876 18396 22932 18398
rect 22540 18284 22596 18340
rect 22988 18338 23044 18340
rect 22988 18286 22990 18338
rect 22990 18286 23042 18338
rect 23042 18286 23044 18338
rect 22988 18284 23044 18286
rect 22204 17388 22260 17444
rect 22652 17442 22708 17444
rect 22652 17390 22654 17442
rect 22654 17390 22706 17442
rect 22706 17390 22708 17442
rect 22652 17388 22708 17390
rect 21308 17052 21364 17108
rect 22092 17052 22148 17108
rect 24522 21194 24578 21196
rect 24522 21142 24524 21194
rect 24524 21142 24576 21194
rect 24576 21142 24578 21194
rect 24522 21140 24578 21142
rect 24626 21194 24682 21196
rect 24626 21142 24628 21194
rect 24628 21142 24680 21194
rect 24680 21142 24682 21194
rect 24626 21140 24682 21142
rect 24730 21194 24786 21196
rect 24730 21142 24732 21194
rect 24732 21142 24784 21194
rect 24784 21142 24786 21194
rect 24730 21140 24786 21142
rect 24332 20972 24388 21028
rect 24444 20748 24500 20804
rect 24220 20076 24276 20132
rect 25004 20748 25060 20804
rect 24892 20412 24948 20468
rect 25004 20300 25060 20356
rect 25564 20802 25620 20804
rect 25564 20750 25566 20802
rect 25566 20750 25618 20802
rect 25618 20750 25620 20802
rect 25564 20748 25620 20750
rect 25564 20412 25620 20468
rect 25340 20188 25396 20244
rect 23996 19852 24052 19908
rect 24668 19740 24724 19796
rect 24522 19626 24578 19628
rect 24522 19574 24524 19626
rect 24524 19574 24576 19626
rect 24576 19574 24578 19626
rect 24522 19572 24578 19574
rect 24626 19626 24682 19628
rect 24626 19574 24628 19626
rect 24628 19574 24680 19626
rect 24680 19574 24682 19626
rect 24626 19572 24682 19574
rect 24730 19626 24786 19628
rect 24730 19574 24732 19626
rect 24732 19574 24784 19626
rect 24784 19574 24786 19626
rect 24730 19572 24786 19574
rect 25228 19740 25284 19796
rect 25228 19292 25284 19348
rect 26572 24834 26628 24836
rect 26572 24782 26574 24834
rect 26574 24782 26626 24834
rect 26626 24782 26628 24834
rect 26572 24780 26628 24782
rect 26348 24444 26404 24500
rect 26460 23378 26516 23380
rect 26460 23326 26462 23378
rect 26462 23326 26514 23378
rect 26514 23326 26516 23378
rect 26460 23324 26516 23326
rect 25788 22204 25844 22260
rect 27804 24722 27860 24724
rect 27804 24670 27806 24722
rect 27806 24670 27858 24722
rect 27858 24670 27860 24722
rect 27804 24668 27860 24670
rect 29184 28250 29240 28252
rect 29184 28198 29186 28250
rect 29186 28198 29238 28250
rect 29238 28198 29240 28250
rect 29184 28196 29240 28198
rect 29288 28250 29344 28252
rect 29288 28198 29290 28250
rect 29290 28198 29342 28250
rect 29342 28198 29344 28250
rect 29288 28196 29344 28198
rect 29392 28250 29448 28252
rect 29392 28198 29394 28250
rect 29394 28198 29446 28250
rect 29446 28198 29448 28250
rect 29392 28196 29448 28198
rect 37212 27580 37268 27636
rect 33846 27466 33902 27468
rect 33846 27414 33848 27466
rect 33848 27414 33900 27466
rect 33900 27414 33902 27466
rect 33846 27412 33902 27414
rect 33950 27466 34006 27468
rect 33950 27414 33952 27466
rect 33952 27414 34004 27466
rect 34004 27414 34006 27466
rect 33950 27412 34006 27414
rect 34054 27466 34110 27468
rect 34054 27414 34056 27466
rect 34056 27414 34108 27466
rect 34108 27414 34110 27466
rect 34054 27412 34110 27414
rect 38220 30268 38276 30324
rect 37660 30098 37716 30100
rect 37660 30046 37662 30098
rect 37662 30046 37714 30098
rect 37714 30046 37716 30098
rect 37660 30044 37716 30046
rect 38220 30098 38276 30100
rect 38220 30046 38222 30098
rect 38222 30046 38274 30098
rect 38274 30046 38276 30098
rect 38220 30044 38276 30046
rect 37884 29986 37940 29988
rect 37884 29934 37886 29986
rect 37886 29934 37938 29986
rect 37938 29934 37940 29986
rect 37884 29932 37940 29934
rect 38892 29932 38948 29988
rect 38508 29818 38564 29820
rect 38508 29766 38510 29818
rect 38510 29766 38562 29818
rect 38562 29766 38564 29818
rect 38508 29764 38564 29766
rect 38612 29818 38668 29820
rect 38612 29766 38614 29818
rect 38614 29766 38666 29818
rect 38666 29766 38668 29818
rect 38612 29764 38668 29766
rect 38716 29818 38772 29820
rect 38716 29766 38718 29818
rect 38718 29766 38770 29818
rect 38770 29766 38772 29818
rect 38716 29764 38772 29766
rect 38220 29596 38276 29652
rect 37100 27020 37156 27076
rect 29184 26682 29240 26684
rect 29184 26630 29186 26682
rect 29186 26630 29238 26682
rect 29238 26630 29240 26682
rect 29184 26628 29240 26630
rect 29288 26682 29344 26684
rect 29288 26630 29290 26682
rect 29290 26630 29342 26682
rect 29342 26630 29344 26682
rect 29288 26628 29344 26630
rect 29392 26682 29448 26684
rect 29392 26630 29394 26682
rect 29394 26630 29446 26682
rect 29446 26630 29448 26682
rect 29392 26628 29448 26630
rect 33846 25898 33902 25900
rect 33846 25846 33848 25898
rect 33848 25846 33900 25898
rect 33900 25846 33902 25898
rect 33846 25844 33902 25846
rect 33950 25898 34006 25900
rect 33950 25846 33952 25898
rect 33952 25846 34004 25898
rect 34004 25846 34006 25898
rect 33950 25844 34006 25846
rect 34054 25898 34110 25900
rect 34054 25846 34056 25898
rect 34056 25846 34108 25898
rect 34108 25846 34110 25898
rect 34054 25844 34110 25846
rect 29184 25114 29240 25116
rect 29184 25062 29186 25114
rect 29186 25062 29238 25114
rect 29238 25062 29240 25114
rect 29184 25060 29240 25062
rect 29288 25114 29344 25116
rect 29288 25062 29290 25114
rect 29290 25062 29342 25114
rect 29342 25062 29344 25114
rect 29288 25060 29344 25062
rect 29392 25114 29448 25116
rect 29392 25062 29394 25114
rect 29394 25062 29446 25114
rect 29446 25062 29448 25114
rect 29392 25060 29448 25062
rect 36988 24668 37044 24724
rect 33846 24330 33902 24332
rect 33846 24278 33848 24330
rect 33848 24278 33900 24330
rect 33900 24278 33902 24330
rect 33846 24276 33902 24278
rect 33950 24330 34006 24332
rect 33950 24278 33952 24330
rect 33952 24278 34004 24330
rect 34004 24278 34006 24330
rect 33950 24276 34006 24278
rect 34054 24330 34110 24332
rect 34054 24278 34056 24330
rect 34056 24278 34108 24330
rect 34108 24278 34110 24330
rect 34054 24276 34110 24278
rect 29184 23546 29240 23548
rect 29184 23494 29186 23546
rect 29186 23494 29238 23546
rect 29238 23494 29240 23546
rect 29184 23492 29240 23494
rect 29288 23546 29344 23548
rect 29288 23494 29290 23546
rect 29290 23494 29342 23546
rect 29342 23494 29344 23546
rect 29288 23492 29344 23494
rect 29392 23546 29448 23548
rect 29392 23494 29394 23546
rect 29394 23494 29446 23546
rect 29446 23494 29448 23546
rect 29392 23492 29448 23494
rect 27020 23212 27076 23268
rect 28476 23154 28532 23156
rect 28476 23102 28478 23154
rect 28478 23102 28530 23154
rect 28530 23102 28532 23154
rect 28476 23100 28532 23102
rect 28812 23100 28868 23156
rect 27692 22876 27748 22932
rect 28812 22876 28868 22932
rect 28252 20972 28308 21028
rect 27132 20802 27188 20804
rect 27132 20750 27134 20802
rect 27134 20750 27186 20802
rect 27186 20750 27188 20802
rect 27132 20748 27188 20750
rect 27804 20690 27860 20692
rect 27804 20638 27806 20690
rect 27806 20638 27858 20690
rect 27858 20638 27860 20690
rect 27804 20636 27860 20638
rect 25788 20412 25844 20468
rect 26908 20018 26964 20020
rect 26908 19966 26910 20018
rect 26910 19966 26962 20018
rect 26962 19966 26964 20018
rect 26908 19964 26964 19966
rect 26572 19906 26628 19908
rect 26572 19854 26574 19906
rect 26574 19854 26626 19906
rect 26626 19854 26628 19906
rect 26572 19852 26628 19854
rect 26236 19740 26292 19796
rect 26236 19234 26292 19236
rect 26236 19182 26238 19234
rect 26238 19182 26290 19234
rect 26290 19182 26292 19234
rect 26236 19180 26292 19182
rect 26348 19122 26404 19124
rect 26348 19070 26350 19122
rect 26350 19070 26402 19122
rect 26402 19070 26404 19122
rect 26348 19068 26404 19070
rect 24522 18058 24578 18060
rect 24522 18006 24524 18058
rect 24524 18006 24576 18058
rect 24576 18006 24578 18058
rect 24522 18004 24578 18006
rect 24626 18058 24682 18060
rect 24626 18006 24628 18058
rect 24628 18006 24680 18058
rect 24680 18006 24682 18058
rect 24626 18004 24682 18006
rect 24730 18058 24786 18060
rect 24730 18006 24732 18058
rect 24732 18006 24784 18058
rect 24784 18006 24786 18058
rect 24730 18004 24786 18006
rect 25340 17554 25396 17556
rect 25340 17502 25342 17554
rect 25342 17502 25394 17554
rect 25394 17502 25396 17554
rect 25340 17500 25396 17502
rect 23884 17442 23940 17444
rect 23884 17390 23886 17442
rect 23886 17390 23938 17442
rect 23938 17390 23940 17442
rect 23884 17388 23940 17390
rect 24220 17442 24276 17444
rect 24220 17390 24222 17442
rect 24222 17390 24274 17442
rect 24274 17390 24276 17442
rect 24220 17388 24276 17390
rect 22988 17052 23044 17108
rect 21196 15372 21252 15428
rect 21644 16268 21700 16324
rect 20636 14700 20692 14756
rect 20412 14476 20468 14532
rect 20412 14306 20468 14308
rect 20412 14254 20414 14306
rect 20414 14254 20466 14306
rect 20466 14254 20468 14306
rect 20412 14252 20468 14254
rect 20636 14530 20692 14532
rect 20636 14478 20638 14530
rect 20638 14478 20690 14530
rect 20690 14478 20692 14530
rect 20636 14476 20692 14478
rect 20524 13692 20580 13748
rect 21308 14812 21364 14868
rect 21532 15314 21588 15316
rect 21532 15262 21534 15314
rect 21534 15262 21586 15314
rect 21586 15262 21588 15314
rect 21532 15260 21588 15262
rect 21420 14588 21476 14644
rect 20300 13468 20356 13524
rect 20076 13020 20132 13076
rect 18956 12738 19012 12740
rect 18956 12686 18958 12738
rect 18958 12686 19010 12738
rect 19010 12686 19012 12738
rect 18956 12684 19012 12686
rect 18956 12402 19012 12404
rect 18956 12350 18958 12402
rect 18958 12350 19010 12402
rect 19010 12350 19012 12402
rect 18956 12348 19012 12350
rect 18732 11788 18788 11844
rect 18620 4620 18676 4676
rect 18620 3554 18676 3556
rect 18620 3502 18622 3554
rect 18622 3502 18674 3554
rect 18674 3502 18676 3554
rect 18620 3500 18676 3502
rect 19860 12570 19916 12572
rect 19860 12518 19862 12570
rect 19862 12518 19914 12570
rect 19914 12518 19916 12570
rect 19860 12516 19916 12518
rect 19964 12570 20020 12572
rect 19964 12518 19966 12570
rect 19966 12518 20018 12570
rect 20018 12518 20020 12570
rect 19964 12516 20020 12518
rect 20068 12570 20124 12572
rect 20068 12518 20070 12570
rect 20070 12518 20122 12570
rect 20122 12518 20124 12570
rect 20068 12516 20124 12518
rect 19292 10108 19348 10164
rect 20076 11116 20132 11172
rect 19516 3612 19572 3668
rect 19860 11002 19916 11004
rect 19860 10950 19862 11002
rect 19862 10950 19914 11002
rect 19914 10950 19916 11002
rect 19860 10948 19916 10950
rect 19964 11002 20020 11004
rect 19964 10950 19966 11002
rect 19966 10950 20018 11002
rect 20018 10950 20020 11002
rect 19964 10948 20020 10950
rect 20068 11002 20124 11004
rect 20068 10950 20070 11002
rect 20070 10950 20122 11002
rect 20122 10950 20124 11002
rect 20068 10948 20124 10950
rect 19860 9434 19916 9436
rect 19860 9382 19862 9434
rect 19862 9382 19914 9434
rect 19914 9382 19916 9434
rect 19860 9380 19916 9382
rect 19964 9434 20020 9436
rect 19964 9382 19966 9434
rect 19966 9382 20018 9434
rect 20018 9382 20020 9434
rect 19964 9380 20020 9382
rect 20068 9434 20124 9436
rect 20068 9382 20070 9434
rect 20070 9382 20122 9434
rect 20122 9382 20124 9434
rect 20068 9380 20124 9382
rect 19860 7866 19916 7868
rect 19860 7814 19862 7866
rect 19862 7814 19914 7866
rect 19914 7814 19916 7866
rect 19860 7812 19916 7814
rect 19964 7866 20020 7868
rect 19964 7814 19966 7866
rect 19966 7814 20018 7866
rect 20018 7814 20020 7866
rect 19964 7812 20020 7814
rect 20068 7866 20124 7868
rect 20068 7814 20070 7866
rect 20070 7814 20122 7866
rect 20122 7814 20124 7866
rect 20068 7812 20124 7814
rect 19860 6298 19916 6300
rect 19860 6246 19862 6298
rect 19862 6246 19914 6298
rect 19914 6246 19916 6298
rect 19860 6244 19916 6246
rect 19964 6298 20020 6300
rect 19964 6246 19966 6298
rect 19966 6246 20018 6298
rect 20018 6246 20020 6298
rect 19964 6244 20020 6246
rect 20068 6298 20124 6300
rect 20068 6246 20070 6298
rect 20070 6246 20122 6298
rect 20122 6246 20124 6298
rect 20068 6244 20124 6246
rect 19860 4730 19916 4732
rect 19860 4678 19862 4730
rect 19862 4678 19914 4730
rect 19914 4678 19916 4730
rect 19860 4676 19916 4678
rect 19964 4730 20020 4732
rect 19964 4678 19966 4730
rect 19966 4678 20018 4730
rect 20018 4678 20020 4730
rect 19964 4676 20020 4678
rect 20068 4730 20124 4732
rect 20068 4678 20070 4730
rect 20070 4678 20122 4730
rect 20122 4678 20124 4730
rect 20068 4676 20124 4678
rect 20748 12684 20804 12740
rect 20636 4508 20692 4564
rect 21532 14476 21588 14532
rect 21420 14418 21476 14420
rect 21420 14366 21422 14418
rect 21422 14366 21474 14418
rect 21474 14366 21476 14418
rect 21420 14364 21476 14366
rect 21196 14252 21252 14308
rect 20972 13692 21028 13748
rect 20972 12684 21028 12740
rect 21084 13580 21140 13636
rect 21308 13468 21364 13524
rect 20860 4508 20916 4564
rect 21084 11116 21140 11172
rect 21644 13020 21700 13076
rect 22428 16994 22484 16996
rect 22428 16942 22430 16994
rect 22430 16942 22482 16994
rect 22482 16942 22484 16994
rect 22428 16940 22484 16942
rect 21980 16716 22036 16772
rect 22316 16716 22372 16772
rect 23660 17052 23716 17108
rect 23100 16882 23156 16884
rect 23100 16830 23102 16882
rect 23102 16830 23154 16882
rect 23154 16830 23156 16882
rect 23100 16828 23156 16830
rect 24220 16828 24276 16884
rect 26348 17612 26404 17668
rect 33846 22762 33902 22764
rect 33846 22710 33848 22762
rect 33848 22710 33900 22762
rect 33900 22710 33902 22762
rect 33846 22708 33902 22710
rect 33950 22762 34006 22764
rect 33950 22710 33952 22762
rect 33952 22710 34004 22762
rect 34004 22710 34006 22762
rect 33950 22708 34006 22710
rect 34054 22762 34110 22764
rect 34054 22710 34056 22762
rect 34056 22710 34108 22762
rect 34108 22710 34110 22762
rect 34054 22708 34110 22710
rect 36540 22258 36596 22260
rect 36540 22206 36542 22258
rect 36542 22206 36594 22258
rect 36594 22206 36596 22258
rect 36540 22204 36596 22206
rect 29184 21978 29240 21980
rect 29184 21926 29186 21978
rect 29186 21926 29238 21978
rect 29238 21926 29240 21978
rect 29184 21924 29240 21926
rect 29288 21978 29344 21980
rect 29288 21926 29290 21978
rect 29290 21926 29342 21978
rect 29342 21926 29344 21978
rect 29288 21924 29344 21926
rect 29392 21978 29448 21980
rect 29392 21926 29394 21978
rect 29394 21926 29446 21978
rect 29446 21926 29448 21978
rect 29392 21924 29448 21926
rect 33846 21194 33902 21196
rect 33846 21142 33848 21194
rect 33848 21142 33900 21194
rect 33900 21142 33902 21194
rect 33846 21140 33902 21142
rect 33950 21194 34006 21196
rect 33950 21142 33952 21194
rect 33952 21142 34004 21194
rect 34004 21142 34006 21194
rect 33950 21140 34006 21142
rect 34054 21194 34110 21196
rect 34054 21142 34056 21194
rect 34056 21142 34108 21194
rect 34108 21142 34110 21194
rect 34054 21140 34110 21142
rect 37324 26962 37380 26964
rect 37324 26910 37326 26962
rect 37326 26910 37378 26962
rect 37378 26910 37380 26962
rect 37324 26908 37380 26910
rect 37212 26178 37268 26180
rect 37212 26126 37214 26178
rect 37214 26126 37266 26178
rect 37266 26126 37268 26178
rect 37212 26124 37268 26126
rect 38220 28924 38276 28980
rect 37884 28700 37940 28756
rect 37660 28642 37716 28644
rect 37660 28590 37662 28642
rect 37662 28590 37714 28642
rect 37714 28590 37716 28642
rect 37660 28588 37716 28590
rect 38108 28642 38164 28644
rect 38108 28590 38110 28642
rect 38110 28590 38162 28642
rect 38162 28590 38164 28642
rect 38108 28588 38164 28590
rect 38508 28250 38564 28252
rect 38508 28198 38510 28250
rect 38510 28198 38562 28250
rect 38562 28198 38564 28250
rect 38508 28196 38564 28198
rect 38612 28250 38668 28252
rect 38612 28198 38614 28250
rect 38614 28198 38666 28250
rect 38666 28198 38668 28250
rect 38612 28196 38668 28198
rect 38716 28250 38772 28252
rect 38716 28198 38718 28250
rect 38718 28198 38770 28250
rect 38770 28198 38772 28250
rect 38716 28196 38772 28198
rect 37660 27074 37716 27076
rect 37660 27022 37662 27074
rect 37662 27022 37714 27074
rect 37714 27022 37716 27074
rect 37660 27020 37716 27022
rect 38220 27580 38276 27636
rect 37772 26908 37828 26964
rect 37660 25394 37716 25396
rect 37660 25342 37662 25394
rect 37662 25342 37714 25394
rect 37714 25342 37716 25394
rect 37660 25340 37716 25342
rect 37884 25282 37940 25284
rect 37884 25230 37886 25282
rect 37886 25230 37938 25282
rect 37938 25230 37940 25282
rect 37884 25228 37940 25230
rect 37436 24556 37492 24612
rect 37324 23212 37380 23268
rect 38108 26236 38164 26292
rect 38220 26124 38276 26180
rect 38220 25564 38276 25620
rect 38220 25394 38276 25396
rect 38220 25342 38222 25394
rect 38222 25342 38274 25394
rect 38274 25342 38276 25394
rect 38220 25340 38276 25342
rect 38220 24892 38276 24948
rect 37996 24780 38052 24836
rect 38220 24220 38276 24276
rect 37660 23714 37716 23716
rect 37660 23662 37662 23714
rect 37662 23662 37714 23714
rect 37714 23662 37716 23714
rect 37660 23660 37716 23662
rect 37548 23100 37604 23156
rect 37660 22876 37716 22932
rect 37212 21474 37268 21476
rect 37212 21422 37214 21474
rect 37214 21422 37266 21474
rect 37266 21422 37268 21474
rect 37212 21420 37268 21422
rect 37100 20972 37156 21028
rect 29184 20410 29240 20412
rect 29184 20358 29186 20410
rect 29186 20358 29238 20410
rect 29238 20358 29240 20410
rect 29184 20356 29240 20358
rect 29288 20410 29344 20412
rect 29288 20358 29290 20410
rect 29290 20358 29342 20410
rect 29342 20358 29344 20410
rect 29288 20356 29344 20358
rect 29392 20410 29448 20412
rect 29392 20358 29394 20410
rect 29394 20358 29446 20410
rect 29446 20358 29448 20410
rect 29392 20356 29448 20358
rect 29932 20412 29988 20468
rect 29932 20188 29988 20244
rect 36988 20076 37044 20132
rect 29932 20018 29988 20020
rect 29932 19966 29934 20018
rect 29934 19966 29986 20018
rect 29986 19966 29988 20018
rect 29932 19964 29988 19966
rect 28476 19794 28532 19796
rect 28476 19742 28478 19794
rect 28478 19742 28530 19794
rect 28530 19742 28532 19794
rect 28476 19740 28532 19742
rect 33846 19626 33902 19628
rect 33846 19574 33848 19626
rect 33848 19574 33900 19626
rect 33900 19574 33902 19626
rect 33846 19572 33902 19574
rect 33950 19626 34006 19628
rect 33950 19574 33952 19626
rect 33952 19574 34004 19626
rect 34004 19574 34006 19626
rect 33950 19572 34006 19574
rect 34054 19626 34110 19628
rect 34054 19574 34056 19626
rect 34056 19574 34108 19626
rect 34108 19574 34110 19626
rect 34054 19572 34110 19574
rect 27692 19404 27748 19460
rect 27580 19234 27636 19236
rect 27580 19182 27582 19234
rect 27582 19182 27634 19234
rect 27634 19182 27636 19234
rect 27580 19180 27636 19182
rect 27468 18956 27524 19012
rect 37548 21586 37604 21588
rect 37548 21534 37550 21586
rect 37550 21534 37602 21586
rect 37602 21534 37604 21586
rect 37548 21532 37604 21534
rect 37436 20300 37492 20356
rect 37324 19964 37380 20020
rect 38220 23660 38276 23716
rect 38508 26682 38564 26684
rect 38508 26630 38510 26682
rect 38510 26630 38562 26682
rect 38562 26630 38564 26682
rect 38508 26628 38564 26630
rect 38612 26682 38668 26684
rect 38612 26630 38614 26682
rect 38614 26630 38666 26682
rect 38666 26630 38668 26682
rect 38612 26628 38668 26630
rect 38716 26682 38772 26684
rect 38716 26630 38718 26682
rect 38718 26630 38770 26682
rect 38770 26630 38772 26682
rect 38716 26628 38772 26630
rect 38508 25114 38564 25116
rect 38508 25062 38510 25114
rect 38510 25062 38562 25114
rect 38562 25062 38564 25114
rect 38508 25060 38564 25062
rect 38612 25114 38668 25116
rect 38612 25062 38614 25114
rect 38614 25062 38666 25114
rect 38666 25062 38668 25114
rect 38612 25060 38668 25062
rect 38716 25114 38772 25116
rect 38716 25062 38718 25114
rect 38718 25062 38770 25114
rect 38770 25062 38772 25114
rect 38716 25060 38772 25062
rect 38508 23546 38564 23548
rect 38508 23494 38510 23546
rect 38510 23494 38562 23546
rect 38562 23494 38564 23546
rect 38508 23492 38564 23494
rect 38612 23546 38668 23548
rect 38612 23494 38614 23546
rect 38614 23494 38666 23546
rect 38666 23494 38668 23546
rect 38612 23492 38668 23494
rect 38716 23546 38772 23548
rect 38716 23494 38718 23546
rect 38718 23494 38770 23546
rect 38770 23494 38772 23546
rect 38716 23492 38772 23494
rect 38332 22988 38388 23044
rect 38220 22876 38276 22932
rect 38220 22258 38276 22260
rect 38220 22206 38222 22258
rect 38222 22206 38274 22258
rect 38274 22206 38276 22258
rect 38220 22204 38276 22206
rect 38508 21978 38564 21980
rect 38508 21926 38510 21978
rect 38510 21926 38562 21978
rect 38562 21926 38564 21978
rect 38508 21924 38564 21926
rect 38612 21978 38668 21980
rect 38612 21926 38614 21978
rect 38614 21926 38666 21978
rect 38666 21926 38668 21978
rect 38612 21924 38668 21926
rect 38716 21978 38772 21980
rect 38716 21926 38718 21978
rect 38718 21926 38770 21978
rect 38770 21926 38772 21978
rect 38716 21924 38772 21926
rect 37996 20860 38052 20916
rect 38220 21420 38276 21476
rect 38220 20860 38276 20916
rect 37884 20748 37940 20804
rect 37884 20578 37940 20580
rect 37884 20526 37886 20578
rect 37886 20526 37938 20578
rect 37938 20526 37940 20578
rect 37884 20524 37940 20526
rect 37660 20188 37716 20244
rect 38892 20636 38948 20692
rect 38508 20410 38564 20412
rect 38508 20358 38510 20410
rect 38510 20358 38562 20410
rect 38562 20358 38564 20410
rect 38508 20356 38564 20358
rect 38612 20410 38668 20412
rect 38612 20358 38614 20410
rect 38614 20358 38666 20410
rect 38666 20358 38668 20410
rect 38612 20356 38668 20358
rect 38716 20410 38772 20412
rect 38716 20358 38718 20410
rect 38718 20358 38770 20410
rect 38770 20358 38772 20410
rect 38716 20356 38772 20358
rect 38220 20188 38276 20244
rect 37884 20130 37940 20132
rect 37884 20078 37886 20130
rect 37886 20078 37938 20130
rect 37938 20078 37940 20130
rect 37884 20076 37940 20078
rect 37548 19852 37604 19908
rect 38220 19516 38276 19572
rect 36988 19180 37044 19236
rect 37884 19292 37940 19348
rect 28476 18956 28532 19012
rect 37660 19010 37716 19012
rect 37660 18958 37662 19010
rect 37662 18958 37714 19010
rect 37714 18958 37716 19010
rect 37660 18956 37716 18958
rect 38220 18956 38276 19012
rect 29184 18842 29240 18844
rect 29184 18790 29186 18842
rect 29186 18790 29238 18842
rect 29238 18790 29240 18842
rect 29184 18788 29240 18790
rect 29288 18842 29344 18844
rect 29288 18790 29290 18842
rect 29290 18790 29342 18842
rect 29342 18790 29344 18842
rect 29288 18788 29344 18790
rect 29392 18842 29448 18844
rect 29392 18790 29394 18842
rect 29394 18790 29446 18842
rect 29446 18790 29448 18842
rect 29392 18788 29448 18790
rect 37772 18844 37828 18900
rect 38508 18842 38564 18844
rect 38508 18790 38510 18842
rect 38510 18790 38562 18842
rect 38562 18790 38564 18842
rect 38508 18788 38564 18790
rect 38612 18842 38668 18844
rect 38612 18790 38614 18842
rect 38614 18790 38666 18842
rect 38666 18790 38668 18842
rect 38612 18788 38668 18790
rect 38716 18842 38772 18844
rect 38716 18790 38718 18842
rect 38718 18790 38770 18842
rect 38770 18790 38772 18842
rect 38716 18788 38772 18790
rect 37660 18172 37716 18228
rect 37884 18284 37940 18340
rect 33846 18058 33902 18060
rect 33846 18006 33848 18058
rect 33848 18006 33900 18058
rect 33900 18006 33902 18058
rect 33846 18004 33902 18006
rect 33950 18058 34006 18060
rect 33950 18006 33952 18058
rect 33952 18006 34004 18058
rect 34004 18006 34006 18058
rect 33950 18004 34006 18006
rect 34054 18058 34110 18060
rect 34054 18006 34056 18058
rect 34056 18006 34108 18058
rect 34108 18006 34110 18058
rect 34054 18004 34110 18006
rect 26908 17388 26964 17444
rect 26908 17164 26964 17220
rect 24522 16490 24578 16492
rect 24522 16438 24524 16490
rect 24524 16438 24576 16490
rect 24576 16438 24578 16490
rect 24522 16436 24578 16438
rect 24626 16490 24682 16492
rect 24626 16438 24628 16490
rect 24628 16438 24680 16490
rect 24680 16438 24682 16490
rect 24626 16436 24682 16438
rect 24730 16490 24786 16492
rect 24730 16438 24732 16490
rect 24732 16438 24784 16490
rect 24784 16438 24786 16490
rect 24730 16436 24786 16438
rect 24522 14922 24578 14924
rect 24522 14870 24524 14922
rect 24524 14870 24576 14922
rect 24576 14870 24578 14922
rect 24522 14868 24578 14870
rect 24626 14922 24682 14924
rect 24626 14870 24628 14922
rect 24628 14870 24680 14922
rect 24680 14870 24682 14922
rect 24626 14868 24682 14870
rect 24730 14922 24786 14924
rect 24730 14870 24732 14922
rect 24732 14870 24784 14922
rect 24784 14870 24786 14922
rect 24730 14868 24786 14870
rect 22204 13916 22260 13972
rect 22092 13804 22148 13860
rect 22204 13746 22260 13748
rect 22204 13694 22206 13746
rect 22206 13694 22258 13746
rect 22258 13694 22260 13746
rect 22204 13692 22260 13694
rect 21532 12348 21588 12404
rect 21420 4844 21476 4900
rect 21756 12738 21812 12740
rect 21756 12686 21758 12738
rect 21758 12686 21810 12738
rect 21810 12686 21812 12738
rect 21756 12684 21812 12686
rect 22876 13858 22932 13860
rect 22876 13806 22878 13858
rect 22878 13806 22930 13858
rect 22930 13806 22932 13858
rect 22876 13804 22932 13806
rect 22764 13020 22820 13076
rect 20860 4338 20916 4340
rect 20860 4286 20862 4338
rect 20862 4286 20914 4338
rect 20914 4286 20916 4338
rect 20860 4284 20916 4286
rect 20300 3388 20356 3444
rect 19860 3162 19916 3164
rect 19860 3110 19862 3162
rect 19862 3110 19914 3162
rect 19914 3110 19916 3162
rect 19860 3108 19916 3110
rect 19964 3162 20020 3164
rect 19964 3110 19966 3162
rect 19966 3110 20018 3162
rect 20018 3110 20020 3162
rect 19964 3108 20020 3110
rect 20068 3162 20124 3164
rect 20068 3110 20070 3162
rect 20070 3110 20122 3162
rect 20122 3110 20124 3162
rect 20068 3108 20124 3110
rect 20972 3666 21028 3668
rect 20972 3614 20974 3666
rect 20974 3614 21026 3666
rect 21026 3614 21028 3666
rect 20972 3612 21028 3614
rect 21532 4284 21588 4340
rect 21980 4338 22036 4340
rect 21980 4286 21982 4338
rect 21982 4286 22034 4338
rect 22034 4286 22036 4338
rect 21980 4284 22036 4286
rect 22428 4562 22484 4564
rect 22428 4510 22430 4562
rect 22430 4510 22482 4562
rect 22482 4510 22484 4562
rect 22428 4508 22484 4510
rect 22988 4956 23044 5012
rect 22988 3388 23044 3444
rect 23772 14306 23828 14308
rect 23772 14254 23774 14306
rect 23774 14254 23826 14306
rect 23826 14254 23828 14306
rect 23772 14252 23828 14254
rect 25004 14530 25060 14532
rect 25004 14478 25006 14530
rect 25006 14478 25058 14530
rect 25058 14478 25060 14530
rect 25004 14476 25060 14478
rect 24892 13916 24948 13972
rect 24220 13804 24276 13860
rect 23772 12908 23828 12964
rect 24522 13354 24578 13356
rect 24522 13302 24524 13354
rect 24524 13302 24576 13354
rect 24576 13302 24578 13354
rect 24522 13300 24578 13302
rect 24626 13354 24682 13356
rect 24626 13302 24628 13354
rect 24628 13302 24680 13354
rect 24680 13302 24682 13354
rect 24626 13300 24682 13302
rect 24730 13354 24786 13356
rect 24730 13302 24732 13354
rect 24732 13302 24784 13354
rect 24784 13302 24786 13354
rect 24730 13300 24786 13302
rect 24332 13020 24388 13076
rect 23772 12738 23828 12740
rect 23772 12686 23774 12738
rect 23774 12686 23826 12738
rect 23826 12686 23828 12738
rect 23772 12684 23828 12686
rect 23660 10332 23716 10388
rect 23548 3724 23604 3780
rect 23660 4844 23716 4900
rect 23436 3388 23492 3444
rect 24522 11786 24578 11788
rect 24522 11734 24524 11786
rect 24524 11734 24576 11786
rect 24576 11734 24578 11786
rect 24522 11732 24578 11734
rect 24626 11786 24682 11788
rect 24626 11734 24628 11786
rect 24628 11734 24680 11786
rect 24680 11734 24682 11786
rect 24626 11732 24682 11734
rect 24730 11786 24786 11788
rect 24730 11734 24732 11786
rect 24732 11734 24784 11786
rect 24784 11734 24786 11786
rect 24730 11732 24786 11734
rect 24522 10218 24578 10220
rect 24522 10166 24524 10218
rect 24524 10166 24576 10218
rect 24576 10166 24578 10218
rect 24522 10164 24578 10166
rect 24626 10218 24682 10220
rect 24626 10166 24628 10218
rect 24628 10166 24680 10218
rect 24680 10166 24682 10218
rect 24626 10164 24682 10166
rect 24730 10218 24786 10220
rect 24730 10166 24732 10218
rect 24732 10166 24784 10218
rect 24784 10166 24786 10218
rect 24730 10164 24786 10166
rect 24522 8650 24578 8652
rect 24522 8598 24524 8650
rect 24524 8598 24576 8650
rect 24576 8598 24578 8650
rect 24522 8596 24578 8598
rect 24626 8650 24682 8652
rect 24626 8598 24628 8650
rect 24628 8598 24680 8650
rect 24680 8598 24682 8650
rect 24626 8596 24682 8598
rect 24730 8650 24786 8652
rect 24730 8598 24732 8650
rect 24732 8598 24784 8650
rect 24784 8598 24786 8650
rect 24730 8596 24786 8598
rect 24522 7082 24578 7084
rect 24522 7030 24524 7082
rect 24524 7030 24576 7082
rect 24576 7030 24578 7082
rect 24522 7028 24578 7030
rect 24626 7082 24682 7084
rect 24626 7030 24628 7082
rect 24628 7030 24680 7082
rect 24680 7030 24682 7082
rect 24626 7028 24682 7030
rect 24730 7082 24786 7084
rect 24730 7030 24732 7082
rect 24732 7030 24784 7082
rect 24784 7030 24786 7082
rect 24730 7028 24786 7030
rect 24522 5514 24578 5516
rect 24522 5462 24524 5514
rect 24524 5462 24576 5514
rect 24576 5462 24578 5514
rect 24522 5460 24578 5462
rect 24626 5514 24682 5516
rect 24626 5462 24628 5514
rect 24628 5462 24680 5514
rect 24680 5462 24682 5514
rect 24626 5460 24682 5462
rect 24730 5514 24786 5516
rect 24730 5462 24732 5514
rect 24732 5462 24784 5514
rect 24784 5462 24786 5514
rect 24730 5460 24786 5462
rect 25452 13746 25508 13748
rect 25452 13694 25454 13746
rect 25454 13694 25506 13746
rect 25506 13694 25508 13746
rect 25452 13692 25508 13694
rect 25900 13132 25956 13188
rect 24892 4508 24948 4564
rect 25788 10332 25844 10388
rect 25004 4396 25060 4452
rect 23884 3388 23940 3444
rect 25228 4956 25284 5012
rect 24522 3946 24578 3948
rect 24522 3894 24524 3946
rect 24524 3894 24576 3946
rect 24576 3894 24578 3946
rect 24522 3892 24578 3894
rect 24626 3946 24682 3948
rect 24626 3894 24628 3946
rect 24628 3894 24680 3946
rect 24680 3894 24682 3946
rect 24626 3892 24682 3894
rect 24730 3946 24786 3948
rect 24730 3894 24732 3946
rect 24732 3894 24784 3946
rect 24784 3894 24786 3946
rect 24730 3892 24786 3894
rect 24892 3500 24948 3556
rect 25004 3388 25060 3444
rect 25452 3554 25508 3556
rect 25452 3502 25454 3554
rect 25454 3502 25506 3554
rect 25506 3502 25508 3554
rect 25452 3500 25508 3502
rect 26796 15820 26852 15876
rect 26348 15372 26404 15428
rect 26012 12236 26068 12292
rect 26572 12908 26628 12964
rect 25900 4956 25956 5012
rect 26124 3500 26180 3556
rect 26348 3388 26404 3444
rect 27468 17388 27524 17444
rect 28140 12908 28196 12964
rect 28252 13132 28308 13188
rect 27356 12796 27412 12852
rect 27132 4562 27188 4564
rect 27132 4510 27134 4562
rect 27134 4510 27186 4562
rect 27186 4510 27188 4562
rect 27132 4508 27188 4510
rect 27244 3724 27300 3780
rect 27468 3554 27524 3556
rect 27468 3502 27470 3554
rect 27470 3502 27522 3554
rect 27522 3502 27524 3554
rect 27468 3500 27524 3502
rect 27916 3500 27972 3556
rect 28140 3500 28196 3556
rect 27692 3388 27748 3444
rect 29260 17554 29316 17556
rect 29260 17502 29262 17554
rect 29262 17502 29314 17554
rect 29314 17502 29316 17554
rect 29260 17500 29316 17502
rect 29596 17500 29652 17556
rect 29184 17274 29240 17276
rect 29184 17222 29186 17274
rect 29186 17222 29238 17274
rect 29238 17222 29240 17274
rect 29184 17220 29240 17222
rect 29288 17274 29344 17276
rect 29288 17222 29290 17274
rect 29290 17222 29342 17274
rect 29342 17222 29344 17274
rect 29288 17220 29344 17222
rect 29392 17274 29448 17276
rect 29392 17222 29394 17274
rect 29394 17222 29446 17274
rect 29446 17222 29448 17274
rect 29392 17220 29448 17222
rect 36540 17554 36596 17556
rect 36540 17502 36542 17554
rect 36542 17502 36594 17554
rect 36594 17502 36596 17554
rect 36540 17500 36596 17502
rect 37212 17052 37268 17108
rect 29596 16940 29652 16996
rect 38220 18172 38276 18228
rect 38220 17554 38276 17556
rect 38220 17502 38222 17554
rect 38222 17502 38274 17554
rect 38274 17502 38276 17554
rect 38220 17500 38276 17502
rect 38508 17274 38564 17276
rect 38508 17222 38510 17274
rect 38510 17222 38562 17274
rect 38562 17222 38564 17274
rect 38508 17220 38564 17222
rect 38612 17274 38668 17276
rect 38612 17222 38614 17274
rect 38614 17222 38666 17274
rect 38666 17222 38668 17274
rect 38612 17220 38668 17222
rect 38716 17274 38772 17276
rect 38716 17222 38718 17274
rect 38718 17222 38770 17274
rect 38770 17222 38772 17274
rect 38716 17220 38772 17222
rect 37324 16940 37380 16996
rect 37212 16882 37268 16884
rect 37212 16830 37214 16882
rect 37214 16830 37266 16882
rect 37266 16830 37268 16882
rect 37212 16828 37268 16830
rect 33846 16490 33902 16492
rect 33846 16438 33848 16490
rect 33848 16438 33900 16490
rect 33900 16438 33902 16490
rect 33846 16436 33902 16438
rect 33950 16490 34006 16492
rect 33950 16438 33952 16490
rect 33952 16438 34004 16490
rect 34004 16438 34006 16490
rect 33950 16436 34006 16438
rect 34054 16490 34110 16492
rect 34054 16438 34056 16490
rect 34056 16438 34108 16490
rect 34108 16438 34110 16490
rect 34054 16436 34110 16438
rect 29184 15706 29240 15708
rect 29184 15654 29186 15706
rect 29186 15654 29238 15706
rect 29238 15654 29240 15706
rect 29184 15652 29240 15654
rect 29288 15706 29344 15708
rect 29288 15654 29290 15706
rect 29290 15654 29342 15706
rect 29342 15654 29344 15706
rect 29288 15652 29344 15654
rect 29392 15706 29448 15708
rect 29392 15654 29394 15706
rect 29394 15654 29446 15706
rect 29446 15654 29448 15706
rect 29392 15652 29448 15654
rect 33846 14922 33902 14924
rect 33846 14870 33848 14922
rect 33848 14870 33900 14922
rect 33900 14870 33902 14922
rect 33846 14868 33902 14870
rect 33950 14922 34006 14924
rect 33950 14870 33952 14922
rect 33952 14870 34004 14922
rect 34004 14870 34006 14922
rect 33950 14868 34006 14870
rect 34054 14922 34110 14924
rect 34054 14870 34056 14922
rect 34056 14870 34108 14922
rect 34108 14870 34110 14922
rect 34054 14868 34110 14870
rect 29036 14252 29092 14308
rect 31052 14476 31108 14532
rect 29184 14138 29240 14140
rect 29184 14086 29186 14138
rect 29186 14086 29238 14138
rect 29238 14086 29240 14138
rect 29184 14084 29240 14086
rect 29288 14138 29344 14140
rect 29288 14086 29290 14138
rect 29290 14086 29342 14138
rect 29342 14086 29344 14138
rect 29288 14084 29344 14086
rect 29392 14138 29448 14140
rect 29392 14086 29394 14138
rect 29394 14086 29446 14138
rect 29446 14086 29448 14138
rect 29392 14084 29448 14086
rect 30380 13580 30436 13636
rect 29184 12570 29240 12572
rect 29184 12518 29186 12570
rect 29186 12518 29238 12570
rect 29238 12518 29240 12570
rect 29184 12516 29240 12518
rect 29288 12570 29344 12572
rect 29288 12518 29290 12570
rect 29290 12518 29342 12570
rect 29342 12518 29344 12570
rect 29288 12516 29344 12518
rect 29392 12570 29448 12572
rect 29392 12518 29394 12570
rect 29394 12518 29446 12570
rect 29446 12518 29448 12570
rect 29392 12516 29448 12518
rect 29184 11002 29240 11004
rect 29184 10950 29186 11002
rect 29186 10950 29238 11002
rect 29238 10950 29240 11002
rect 29184 10948 29240 10950
rect 29288 11002 29344 11004
rect 29288 10950 29290 11002
rect 29290 10950 29342 11002
rect 29342 10950 29344 11002
rect 29288 10948 29344 10950
rect 29392 11002 29448 11004
rect 29392 10950 29394 11002
rect 29394 10950 29446 11002
rect 29446 10950 29448 11002
rect 29392 10948 29448 10950
rect 28476 10668 28532 10724
rect 29184 9434 29240 9436
rect 29184 9382 29186 9434
rect 29186 9382 29238 9434
rect 29238 9382 29240 9434
rect 29184 9380 29240 9382
rect 29288 9434 29344 9436
rect 29288 9382 29290 9434
rect 29290 9382 29342 9434
rect 29342 9382 29344 9434
rect 29288 9380 29344 9382
rect 29392 9434 29448 9436
rect 29392 9382 29394 9434
rect 29394 9382 29446 9434
rect 29446 9382 29448 9434
rect 29392 9380 29448 9382
rect 29184 7866 29240 7868
rect 29184 7814 29186 7866
rect 29186 7814 29238 7866
rect 29238 7814 29240 7866
rect 29184 7812 29240 7814
rect 29288 7866 29344 7868
rect 29288 7814 29290 7866
rect 29290 7814 29342 7866
rect 29342 7814 29344 7866
rect 29288 7812 29344 7814
rect 29392 7866 29448 7868
rect 29392 7814 29394 7866
rect 29394 7814 29446 7866
rect 29446 7814 29448 7866
rect 29392 7812 29448 7814
rect 29184 6298 29240 6300
rect 29184 6246 29186 6298
rect 29186 6246 29238 6298
rect 29238 6246 29240 6298
rect 29184 6244 29240 6246
rect 29288 6298 29344 6300
rect 29288 6246 29290 6298
rect 29290 6246 29342 6298
rect 29342 6246 29344 6298
rect 29288 6244 29344 6246
rect 29392 6298 29448 6300
rect 29392 6246 29394 6298
rect 29394 6246 29446 6298
rect 29446 6246 29448 6298
rect 29392 6244 29448 6246
rect 29036 4956 29092 5012
rect 28812 3500 28868 3556
rect 28588 3388 28644 3444
rect 29184 4730 29240 4732
rect 29184 4678 29186 4730
rect 29186 4678 29238 4730
rect 29238 4678 29240 4730
rect 29184 4676 29240 4678
rect 29288 4730 29344 4732
rect 29288 4678 29290 4730
rect 29290 4678 29342 4730
rect 29342 4678 29344 4730
rect 29288 4676 29344 4678
rect 29392 4730 29448 4732
rect 29392 4678 29394 4730
rect 29394 4678 29446 4730
rect 29446 4678 29448 4730
rect 29392 4676 29448 4678
rect 29708 4396 29764 4452
rect 29372 3442 29428 3444
rect 29372 3390 29374 3442
rect 29374 3390 29426 3442
rect 29426 3390 29428 3442
rect 29372 3388 29428 3390
rect 29596 3388 29652 3444
rect 29184 3162 29240 3164
rect 29184 3110 29186 3162
rect 29186 3110 29238 3162
rect 29238 3110 29240 3162
rect 29184 3108 29240 3110
rect 29288 3162 29344 3164
rect 29288 3110 29290 3162
rect 29290 3110 29342 3162
rect 29342 3110 29344 3162
rect 29288 3108 29344 3110
rect 29392 3162 29448 3164
rect 29392 3110 29394 3162
rect 29394 3110 29446 3162
rect 29446 3110 29448 3162
rect 29392 3108 29448 3110
rect 30156 3388 30212 3444
rect 30604 3388 30660 3444
rect 33846 13354 33902 13356
rect 33846 13302 33848 13354
rect 33848 13302 33900 13354
rect 33900 13302 33902 13354
rect 33846 13300 33902 13302
rect 33950 13354 34006 13356
rect 33950 13302 33952 13354
rect 33952 13302 34004 13354
rect 34004 13302 34006 13354
rect 33950 13300 34006 13302
rect 34054 13354 34110 13356
rect 34054 13302 34056 13354
rect 34056 13302 34108 13354
rect 34108 13302 34110 13354
rect 34054 13300 34110 13302
rect 37212 12850 37268 12852
rect 37212 12798 37214 12850
rect 37214 12798 37266 12850
rect 37266 12798 37268 12850
rect 37212 12796 37268 12798
rect 36540 12738 36596 12740
rect 36540 12686 36542 12738
rect 36542 12686 36594 12738
rect 36594 12686 36596 12738
rect 36540 12684 36596 12686
rect 37212 12066 37268 12068
rect 37212 12014 37214 12066
rect 37214 12014 37266 12066
rect 37266 12014 37268 12066
rect 37212 12012 37268 12014
rect 37548 16994 37604 16996
rect 37548 16942 37550 16994
rect 37550 16942 37602 16994
rect 37602 16942 37604 16994
rect 37548 16940 37604 16942
rect 37884 16716 37940 16772
rect 38220 16882 38276 16884
rect 38220 16830 38222 16882
rect 38222 16830 38274 16882
rect 38274 16830 38276 16882
rect 38220 16828 38276 16830
rect 38220 16156 38276 16212
rect 37884 15874 37940 15876
rect 37884 15822 37886 15874
rect 37886 15822 37938 15874
rect 37938 15822 37940 15874
rect 37884 15820 37940 15822
rect 37660 15484 37716 15540
rect 38508 15706 38564 15708
rect 38508 15654 38510 15706
rect 38510 15654 38562 15706
rect 38562 15654 38564 15706
rect 38508 15652 38564 15654
rect 38612 15706 38668 15708
rect 38612 15654 38614 15706
rect 38614 15654 38666 15706
rect 38666 15654 38668 15706
rect 38612 15652 38668 15654
rect 38716 15706 38772 15708
rect 38716 15654 38718 15706
rect 38718 15654 38770 15706
rect 38770 15654 38772 15706
rect 38716 15652 38772 15654
rect 38220 15484 38276 15540
rect 37884 15426 37940 15428
rect 37884 15374 37886 15426
rect 37886 15374 37938 15426
rect 37938 15374 37940 15426
rect 37884 15372 37940 15374
rect 38220 14812 38276 14868
rect 37660 14418 37716 14420
rect 37660 14366 37662 14418
rect 37662 14366 37714 14418
rect 37714 14366 37716 14418
rect 37660 14364 37716 14366
rect 37884 14306 37940 14308
rect 37884 14254 37886 14306
rect 37886 14254 37938 14306
rect 37938 14254 37940 14306
rect 37884 14252 37940 14254
rect 38220 14252 38276 14308
rect 38508 14138 38564 14140
rect 38508 14086 38510 14138
rect 38510 14086 38562 14138
rect 38562 14086 38564 14138
rect 38508 14084 38564 14086
rect 38612 14138 38668 14140
rect 38612 14086 38614 14138
rect 38614 14086 38666 14138
rect 38666 14086 38668 14138
rect 38612 14084 38668 14086
rect 38716 14138 38772 14140
rect 38716 14086 38718 14138
rect 38718 14086 38770 14138
rect 38770 14086 38772 14138
rect 38716 14084 38772 14086
rect 37884 13970 37940 13972
rect 37884 13918 37886 13970
rect 37886 13918 37938 13970
rect 37938 13918 37940 13970
rect 37884 13916 37940 13918
rect 37660 13468 37716 13524
rect 38220 13468 38276 13524
rect 37884 12908 37940 12964
rect 38220 12850 38276 12852
rect 38220 12798 38222 12850
rect 38222 12798 38274 12850
rect 38274 12798 38276 12850
rect 38220 12796 38276 12798
rect 38508 12570 38564 12572
rect 38508 12518 38510 12570
rect 38510 12518 38562 12570
rect 38562 12518 38564 12570
rect 38508 12516 38564 12518
rect 38612 12570 38668 12572
rect 38612 12518 38614 12570
rect 38614 12518 38666 12570
rect 38666 12518 38668 12570
rect 38612 12516 38668 12518
rect 38716 12570 38772 12572
rect 38716 12518 38718 12570
rect 38718 12518 38770 12570
rect 38770 12518 38772 12570
rect 38716 12516 38772 12518
rect 37884 12290 37940 12292
rect 37884 12238 37886 12290
rect 37886 12238 37938 12290
rect 37938 12238 37940 12290
rect 37884 12236 37940 12238
rect 37548 12178 37604 12180
rect 37548 12126 37550 12178
rect 37550 12126 37602 12178
rect 37602 12126 37604 12178
rect 37548 12124 37604 12126
rect 38220 12012 38276 12068
rect 33846 11786 33902 11788
rect 33846 11734 33848 11786
rect 33848 11734 33900 11786
rect 33900 11734 33902 11786
rect 33846 11732 33902 11734
rect 33950 11786 34006 11788
rect 33950 11734 33952 11786
rect 33952 11734 34004 11786
rect 34004 11734 34006 11786
rect 33950 11732 34006 11734
rect 34054 11786 34110 11788
rect 34054 11734 34056 11786
rect 34056 11734 34108 11786
rect 34108 11734 34110 11786
rect 34054 11732 34110 11734
rect 38220 11452 38276 11508
rect 37660 10780 37716 10836
rect 38508 11002 38564 11004
rect 38508 10950 38510 11002
rect 38510 10950 38562 11002
rect 38562 10950 38564 11002
rect 38508 10948 38564 10950
rect 38612 11002 38668 11004
rect 38612 10950 38614 11002
rect 38614 10950 38666 11002
rect 38666 10950 38668 11002
rect 38612 10948 38668 10950
rect 38716 11002 38772 11004
rect 38716 10950 38718 11002
rect 38718 10950 38770 11002
rect 38770 10950 38772 11002
rect 38716 10948 38772 10950
rect 38220 10780 38276 10836
rect 37884 10722 37940 10724
rect 37884 10670 37886 10722
rect 37886 10670 37938 10722
rect 37938 10670 37940 10722
rect 37884 10668 37940 10670
rect 37660 10610 37716 10612
rect 37660 10558 37662 10610
rect 37662 10558 37714 10610
rect 37714 10558 37716 10610
rect 37660 10556 37716 10558
rect 38220 10610 38276 10612
rect 38220 10558 38222 10610
rect 38222 10558 38274 10610
rect 38274 10558 38276 10610
rect 38220 10556 38276 10558
rect 33846 10218 33902 10220
rect 33846 10166 33848 10218
rect 33848 10166 33900 10218
rect 33900 10166 33902 10218
rect 33846 10164 33902 10166
rect 33950 10218 34006 10220
rect 33950 10166 33952 10218
rect 33952 10166 34004 10218
rect 34004 10166 34006 10218
rect 33950 10164 34006 10166
rect 34054 10218 34110 10220
rect 34054 10166 34056 10218
rect 34056 10166 34108 10218
rect 34108 10166 34110 10218
rect 34054 10164 34110 10166
rect 38220 10108 38276 10164
rect 38508 9434 38564 9436
rect 38508 9382 38510 9434
rect 38510 9382 38562 9434
rect 38562 9382 38564 9434
rect 38508 9380 38564 9382
rect 38612 9434 38668 9436
rect 38612 9382 38614 9434
rect 38614 9382 38666 9434
rect 38666 9382 38668 9434
rect 38612 9380 38668 9382
rect 38716 9434 38772 9436
rect 38716 9382 38718 9434
rect 38718 9382 38770 9434
rect 38770 9382 38772 9434
rect 38716 9380 38772 9382
rect 33846 8650 33902 8652
rect 33846 8598 33848 8650
rect 33848 8598 33900 8650
rect 33900 8598 33902 8650
rect 33846 8596 33902 8598
rect 33950 8650 34006 8652
rect 33950 8598 33952 8650
rect 33952 8598 34004 8650
rect 34004 8598 34006 8650
rect 33950 8596 34006 8598
rect 34054 8650 34110 8652
rect 34054 8598 34056 8650
rect 34056 8598 34108 8650
rect 34108 8598 34110 8650
rect 34054 8596 34110 8598
rect 38508 7866 38564 7868
rect 38508 7814 38510 7866
rect 38510 7814 38562 7866
rect 38562 7814 38564 7866
rect 38508 7812 38564 7814
rect 38612 7866 38668 7868
rect 38612 7814 38614 7866
rect 38614 7814 38666 7866
rect 38666 7814 38668 7866
rect 38612 7812 38668 7814
rect 38716 7866 38772 7868
rect 38716 7814 38718 7866
rect 38718 7814 38770 7866
rect 38770 7814 38772 7866
rect 38716 7812 38772 7814
rect 33846 7082 33902 7084
rect 33846 7030 33848 7082
rect 33848 7030 33900 7082
rect 33900 7030 33902 7082
rect 33846 7028 33902 7030
rect 33950 7082 34006 7084
rect 33950 7030 33952 7082
rect 33952 7030 34004 7082
rect 34004 7030 34006 7082
rect 33950 7028 34006 7030
rect 34054 7082 34110 7084
rect 34054 7030 34056 7082
rect 34056 7030 34108 7082
rect 34108 7030 34110 7082
rect 34054 7028 34110 7030
rect 38508 6298 38564 6300
rect 38508 6246 38510 6298
rect 38510 6246 38562 6298
rect 38562 6246 38564 6298
rect 38508 6244 38564 6246
rect 38612 6298 38668 6300
rect 38612 6246 38614 6298
rect 38614 6246 38666 6298
rect 38666 6246 38668 6298
rect 38612 6244 38668 6246
rect 38716 6298 38772 6300
rect 38716 6246 38718 6298
rect 38718 6246 38770 6298
rect 38770 6246 38772 6298
rect 38716 6244 38772 6246
rect 33846 5514 33902 5516
rect 33846 5462 33848 5514
rect 33848 5462 33900 5514
rect 33900 5462 33902 5514
rect 33846 5460 33902 5462
rect 33950 5514 34006 5516
rect 33950 5462 33952 5514
rect 33952 5462 34004 5514
rect 34004 5462 34006 5514
rect 33950 5460 34006 5462
rect 34054 5514 34110 5516
rect 34054 5462 34056 5514
rect 34056 5462 34108 5514
rect 34108 5462 34110 5514
rect 34054 5460 34110 5462
rect 38508 4730 38564 4732
rect 38508 4678 38510 4730
rect 38510 4678 38562 4730
rect 38562 4678 38564 4730
rect 38508 4676 38564 4678
rect 38612 4730 38668 4732
rect 38612 4678 38614 4730
rect 38614 4678 38666 4730
rect 38666 4678 38668 4730
rect 38612 4676 38668 4678
rect 38716 4730 38772 4732
rect 38716 4678 38718 4730
rect 38718 4678 38770 4730
rect 38770 4678 38772 4730
rect 38716 4676 38772 4678
rect 33846 3946 33902 3948
rect 33846 3894 33848 3946
rect 33848 3894 33900 3946
rect 33900 3894 33902 3946
rect 33846 3892 33902 3894
rect 33950 3946 34006 3948
rect 33950 3894 33952 3946
rect 33952 3894 34004 3946
rect 34004 3894 34006 3946
rect 33950 3892 34006 3894
rect 34054 3946 34110 3948
rect 34054 3894 34056 3946
rect 34056 3894 34108 3946
rect 34108 3894 34110 3946
rect 34054 3892 34110 3894
rect 38508 3162 38564 3164
rect 38508 3110 38510 3162
rect 38510 3110 38562 3162
rect 38562 3110 38564 3162
rect 38508 3108 38564 3110
rect 38612 3162 38668 3164
rect 38612 3110 38614 3162
rect 38614 3110 38666 3162
rect 38666 3110 38668 3162
rect 38612 3108 38668 3110
rect 38716 3162 38772 3164
rect 38716 3110 38718 3162
rect 38718 3110 38770 3162
rect 38770 3110 38772 3162
rect 38716 3108 38772 3110
<< metal3 >>
rect 10770 36876 10780 36932
rect 10836 36876 11452 36932
rect 11508 36876 11518 36932
rect 20178 36876 20188 36932
rect 20244 36876 21420 36932
rect 21476 36876 21486 36932
rect 26226 36876 26236 36932
rect 26292 36876 27468 36932
rect 27524 36876 28476 36932
rect 28532 36876 28542 36932
rect 5864 36820 5874 36876
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 6138 36820 6148 36876
rect 15188 36820 15198 36876
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15462 36820 15472 36876
rect 24512 36820 24522 36876
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24786 36820 24796 36876
rect 33836 36820 33846 36876
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 34110 36820 34120 36876
rect 24210 36764 24220 36820
rect 24276 36764 24286 36820
rect 24220 36708 24276 36764
rect 16146 36652 16156 36708
rect 16212 36652 17164 36708
rect 17220 36652 17230 36708
rect 20850 36652 20860 36708
rect 20916 36652 22092 36708
rect 22148 36652 22158 36708
rect 24220 36652 25452 36708
rect 25508 36652 25518 36708
rect 24882 36540 24892 36596
rect 24948 36540 26292 36596
rect 26236 36484 26292 36540
rect 16146 36428 16156 36484
rect 16212 36428 16492 36484
rect 16548 36428 16828 36484
rect 16884 36428 16894 36484
rect 22866 36428 22876 36484
rect 22932 36428 24780 36484
rect 24836 36428 24846 36484
rect 26226 36428 26236 36484
rect 26292 36428 26302 36484
rect 10658 36316 10668 36372
rect 10724 36316 11676 36372
rect 11732 36316 11742 36372
rect 11890 36204 11900 36260
rect 11956 36204 19628 36260
rect 19684 36204 19694 36260
rect 24994 36204 25004 36260
rect 25060 36204 26572 36260
rect 26628 36204 26638 36260
rect 10526 36036 10536 36092
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10800 36036 10810 36092
rect 19850 36036 19860 36092
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 20124 36036 20134 36092
rect 29174 36036 29184 36092
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29448 36036 29458 36092
rect 38498 36036 38508 36092
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38772 36036 38782 36092
rect 18050 35756 18060 35812
rect 18116 35756 19292 35812
rect 19348 35756 19358 35812
rect 22194 35756 22204 35812
rect 22260 35756 23100 35812
rect 23156 35756 23548 35812
rect 23604 35756 23614 35812
rect 23986 35756 23996 35812
rect 24052 35756 24062 35812
rect 23996 35700 24052 35756
rect 22754 35644 22764 35700
rect 22820 35644 24052 35700
rect 24210 35420 24220 35476
rect 24276 35420 25228 35476
rect 25284 35420 25294 35476
rect 19394 35308 19404 35364
rect 19460 35308 20860 35364
rect 20916 35308 20926 35364
rect 5864 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6148 35308
rect 15188 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15472 35308
rect 24512 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24796 35308
rect 33836 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34120 35308
rect 22642 34860 22652 34916
rect 22708 34860 24332 34916
rect 24388 34860 24398 34916
rect 10526 34468 10536 34524
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10800 34468 10810 34524
rect 19850 34468 19860 34524
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 20124 34468 20134 34524
rect 29174 34468 29184 34524
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29448 34468 29458 34524
rect 38498 34468 38508 34524
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38772 34468 38782 34524
rect 5864 33684 5874 33740
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 6138 33684 6148 33740
rect 15188 33684 15198 33740
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15462 33684 15472 33740
rect 24512 33684 24522 33740
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24786 33684 24796 33740
rect 33836 33684 33846 33740
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 34110 33684 34120 33740
rect 24882 33516 24892 33572
rect 24948 33516 27468 33572
rect 27524 33516 27534 33572
rect 23986 33404 23996 33460
rect 24052 33404 27132 33460
rect 27188 33404 27198 33460
rect 10526 32900 10536 32956
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10800 32900 10810 32956
rect 19850 32900 19860 32956
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 20124 32900 20134 32956
rect 29174 32900 29184 32956
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29448 32900 29458 32956
rect 38498 32900 38508 32956
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38772 32900 38782 32956
rect 21858 32284 21868 32340
rect 21924 32284 25788 32340
rect 25844 32284 25854 32340
rect 5864 32116 5874 32172
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 6138 32116 6148 32172
rect 15188 32116 15198 32172
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15462 32116 15472 32172
rect 24512 32116 24522 32172
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24786 32116 24796 32172
rect 33836 32116 33846 32172
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 34110 32116 34120 32172
rect 20626 31948 20636 32004
rect 20692 31948 22092 32004
rect 22148 31948 22158 32004
rect 22194 31500 22204 31556
rect 22260 31500 23324 31556
rect 23380 31500 23390 31556
rect 10526 31332 10536 31388
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10800 31332 10810 31388
rect 19850 31332 19860 31388
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 20124 31332 20134 31388
rect 29174 31332 29184 31388
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29448 31332 29458 31388
rect 38498 31332 38508 31388
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38772 31332 38782 31388
rect 5864 30548 5874 30604
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 6138 30548 6148 30604
rect 15188 30548 15198 30604
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15462 30548 15472 30604
rect 24512 30548 24522 30604
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24786 30548 24796 30604
rect 33836 30548 33846 30604
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 34110 30548 34120 30604
rect 39200 30324 40000 30352
rect 38210 30268 38220 30324
rect 38276 30268 40000 30324
rect 39200 30240 40000 30268
rect 37650 30044 37660 30100
rect 37716 30044 38220 30100
rect 38276 30044 38286 30100
rect 37874 29932 37884 29988
rect 37940 29932 38892 29988
rect 38948 29932 38958 29988
rect 10526 29764 10536 29820
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10800 29764 10810 29820
rect 19850 29764 19860 29820
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 20124 29764 20134 29820
rect 29174 29764 29184 29820
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29448 29764 29458 29820
rect 38498 29764 38508 29820
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38772 29764 38782 29820
rect 39200 29652 40000 29680
rect 38210 29596 38220 29652
rect 38276 29596 40000 29652
rect 39200 29568 40000 29596
rect 4274 29372 4284 29428
rect 4340 29372 16100 29428
rect 1922 29148 1932 29204
rect 1988 29148 1998 29204
rect 14354 29148 14364 29204
rect 14420 29148 15820 29204
rect 15876 29148 15886 29204
rect 0 28980 800 29008
rect 1932 28980 1988 29148
rect 16044 29092 16100 29372
rect 15922 29036 15932 29092
rect 15988 29036 16100 29092
rect 5864 28980 5874 29036
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 6138 28980 6148 29036
rect 15188 28980 15198 29036
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15462 28980 15472 29036
rect 24512 28980 24522 29036
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24786 28980 24796 29036
rect 33836 28980 33846 29036
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 34110 28980 34120 29036
rect 39200 28980 40000 29008
rect 0 28924 1988 28980
rect 38210 28924 38220 28980
rect 38276 28924 40000 28980
rect 0 28896 800 28924
rect 39200 28896 40000 28924
rect 15026 28812 15036 28868
rect 15092 28812 15708 28868
rect 15764 28812 15774 28868
rect 28690 28700 28700 28756
rect 28756 28700 37884 28756
rect 37940 28700 37950 28756
rect 37650 28588 37660 28644
rect 37716 28588 38108 28644
rect 38164 28588 38948 28644
rect 0 28308 800 28336
rect 38892 28308 38948 28588
rect 39200 28308 40000 28336
rect 0 28252 1708 28308
rect 1764 28252 2492 28308
rect 2548 28252 2558 28308
rect 38892 28252 40000 28308
rect 0 28224 800 28252
rect 10526 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10810 28252
rect 19850 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20134 28252
rect 29174 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29458 28252
rect 38498 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38782 28252
rect 39200 28224 40000 28252
rect 15026 27804 15036 27860
rect 15092 27804 19516 27860
rect 19572 27804 19582 27860
rect 0 27636 800 27664
rect 39200 27636 40000 27664
rect 0 27580 1708 27636
rect 1764 27580 2940 27636
rect 2996 27580 3006 27636
rect 37202 27580 37212 27636
rect 37268 27580 38220 27636
rect 38276 27580 40000 27636
rect 0 27552 800 27580
rect 39200 27552 40000 27580
rect 5864 27412 5874 27468
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 6138 27412 6148 27468
rect 15188 27412 15198 27468
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15462 27412 15472 27468
rect 24512 27412 24522 27468
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24786 27412 24796 27468
rect 33836 27412 33846 27468
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 34110 27412 34120 27468
rect 2034 27244 2044 27300
rect 2100 27244 13580 27300
rect 13636 27244 13646 27300
rect 20402 27244 20412 27300
rect 20468 27244 21084 27300
rect 21140 27244 21150 27300
rect 12562 27132 12572 27188
rect 12628 27132 17500 27188
rect 17556 27132 17566 27188
rect 15092 27020 16492 27076
rect 16548 27020 17612 27076
rect 17668 27020 17678 27076
rect 37090 27020 37100 27076
rect 37156 27020 37660 27076
rect 37716 27020 37726 27076
rect 0 26964 800 26992
rect 15092 26964 15148 27020
rect 39200 26964 40000 26992
rect 0 26908 2380 26964
rect 2436 26908 3164 26964
rect 3220 26908 3230 26964
rect 12562 26908 12572 26964
rect 12628 26908 15148 26964
rect 20290 26908 20300 26964
rect 20356 26908 21308 26964
rect 21364 26908 21374 26964
rect 37314 26908 37324 26964
rect 37380 26908 37772 26964
rect 37828 26908 40000 26964
rect 0 26880 800 26908
rect 39200 26880 40000 26908
rect 10526 26628 10536 26684
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10800 26628 10810 26684
rect 19850 26628 19860 26684
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 20124 26628 20134 26684
rect 29174 26628 29184 26684
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29448 26628 29458 26684
rect 38498 26628 38508 26684
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38772 26628 38782 26684
rect 11218 26460 11228 26516
rect 11284 26460 17724 26516
rect 17780 26460 20188 26516
rect 2034 26348 2044 26404
rect 2100 26348 14364 26404
rect 14420 26348 14430 26404
rect 0 26292 800 26320
rect 20132 26292 20188 26460
rect 39200 26292 40000 26320
rect 0 26236 1820 26292
rect 1876 26236 1886 26292
rect 14802 26236 14812 26292
rect 14868 26236 16604 26292
rect 16660 26236 16670 26292
rect 20132 26236 20972 26292
rect 21028 26236 21038 26292
rect 38098 26236 38108 26292
rect 38164 26236 40000 26292
rect 0 26208 800 26236
rect 39200 26208 40000 26236
rect 1698 26124 1708 26180
rect 1764 26124 2492 26180
rect 2548 26124 2558 26180
rect 20626 26124 20636 26180
rect 20692 26124 21420 26180
rect 21476 26124 21756 26180
rect 21812 26124 21822 26180
rect 37202 26124 37212 26180
rect 37268 26124 38220 26180
rect 38276 26124 38286 26180
rect 5864 25844 5874 25900
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 6138 25844 6148 25900
rect 15188 25844 15198 25900
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15462 25844 15472 25900
rect 24512 25844 24522 25900
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24786 25844 24796 25900
rect 33836 25844 33846 25900
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 34110 25844 34120 25900
rect 0 25620 800 25648
rect 39200 25620 40000 25648
rect 0 25564 1708 25620
rect 1764 25564 1774 25620
rect 38210 25564 38220 25620
rect 38276 25564 40000 25620
rect 0 25536 800 25564
rect 39200 25536 40000 25564
rect 16482 25452 16492 25508
rect 16548 25452 17388 25508
rect 17444 25452 17454 25508
rect 12898 25340 12908 25396
rect 12964 25340 13692 25396
rect 13748 25340 13758 25396
rect 21522 25340 21532 25396
rect 21588 25340 22876 25396
rect 22932 25340 22942 25396
rect 37650 25340 37660 25396
rect 37716 25340 38220 25396
rect 38276 25340 38286 25396
rect 2034 25228 2044 25284
rect 2100 25228 12348 25284
rect 12404 25228 12414 25284
rect 17042 25228 17052 25284
rect 17108 25228 18620 25284
rect 18676 25228 18686 25284
rect 20178 25228 20188 25284
rect 20244 25228 21196 25284
rect 21252 25228 21262 25284
rect 21634 25228 21644 25284
rect 21700 25228 22540 25284
rect 22596 25228 22606 25284
rect 26450 25228 26460 25284
rect 26516 25228 37884 25284
rect 37940 25228 37950 25284
rect 10526 25060 10536 25116
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10800 25060 10810 25116
rect 19850 25060 19860 25116
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 20124 25060 20134 25116
rect 29174 25060 29184 25116
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29448 25060 29458 25116
rect 38498 25060 38508 25116
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38772 25060 38782 25116
rect 0 24948 800 24976
rect 39200 24948 40000 24976
rect 0 24892 1708 24948
rect 1764 24892 2492 24948
rect 2548 24892 2558 24948
rect 13794 24892 13804 24948
rect 13860 24892 17948 24948
rect 18004 24892 18014 24948
rect 21298 24892 21308 24948
rect 21364 24892 22876 24948
rect 22932 24892 22942 24948
rect 38210 24892 38220 24948
rect 38276 24892 40000 24948
rect 0 24864 800 24892
rect 39200 24864 40000 24892
rect 16258 24780 16268 24836
rect 16324 24780 22652 24836
rect 22708 24780 22718 24836
rect 22978 24780 22988 24836
rect 23044 24780 26572 24836
rect 26628 24780 26638 24836
rect 37986 24780 37996 24836
rect 38052 24780 38062 24836
rect 13122 24668 13132 24724
rect 13188 24668 14700 24724
rect 14756 24668 14766 24724
rect 19730 24668 19740 24724
rect 19796 24668 20300 24724
rect 20356 24668 20366 24724
rect 20962 24668 20972 24724
rect 21028 24668 21038 24724
rect 27794 24668 27804 24724
rect 27860 24668 36988 24724
rect 37044 24668 37054 24724
rect 20972 24612 21028 24668
rect 16706 24556 16716 24612
rect 16772 24556 21028 24612
rect 25554 24556 25564 24612
rect 25620 24556 37436 24612
rect 37492 24556 37502 24612
rect 37996 24500 38052 24780
rect 12450 24444 12460 24500
rect 12516 24444 14700 24500
rect 14756 24444 15596 24500
rect 15652 24444 15662 24500
rect 26338 24444 26348 24500
rect 26404 24444 38052 24500
rect 0 24276 800 24304
rect 5864 24276 5874 24332
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 6138 24276 6148 24332
rect 15188 24276 15198 24332
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15462 24276 15472 24332
rect 24512 24276 24522 24332
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24786 24276 24796 24332
rect 33836 24276 33846 24332
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 34110 24276 34120 24332
rect 39200 24276 40000 24304
rect 0 24220 1708 24276
rect 1764 24220 2492 24276
rect 2548 24220 2558 24276
rect 38210 24220 38220 24276
rect 38276 24220 40000 24276
rect 0 24192 800 24220
rect 39200 24192 40000 24220
rect 13346 24108 13356 24164
rect 13412 24108 17836 24164
rect 17892 24108 17902 24164
rect 2706 23996 2716 24052
rect 2772 23996 14364 24052
rect 14420 23996 14430 24052
rect 16706 23996 16716 24052
rect 16772 23996 18732 24052
rect 18788 23996 18798 24052
rect 16370 23884 16380 23940
rect 16436 23884 17500 23940
rect 17556 23884 17566 23940
rect 2034 23660 2044 23716
rect 2100 23660 12404 23716
rect 37650 23660 37660 23716
rect 37716 23660 38220 23716
rect 38276 23660 38948 23716
rect 0 23604 800 23632
rect 12348 23604 12404 23660
rect 38892 23604 38948 23660
rect 39200 23604 40000 23632
rect 0 23548 1708 23604
rect 1764 23548 2492 23604
rect 2548 23548 2558 23604
rect 12338 23548 12348 23604
rect 12404 23548 12414 23604
rect 38892 23548 40000 23604
rect 0 23520 800 23548
rect 10526 23492 10536 23548
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10800 23492 10810 23548
rect 19850 23492 19860 23548
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 20124 23492 20134 23548
rect 29174 23492 29184 23548
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29448 23492 29458 23548
rect 38498 23492 38508 23548
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38772 23492 38782 23548
rect 39200 23520 40000 23548
rect 15586 23436 15596 23492
rect 15652 23436 16492 23492
rect 16548 23436 17388 23492
rect 17444 23436 17454 23492
rect 21522 23324 21532 23380
rect 21588 23324 26460 23380
rect 26516 23324 26526 23380
rect 2034 23212 2044 23268
rect 2100 23212 8428 23268
rect 16706 23212 16716 23268
rect 16772 23212 20188 23268
rect 20244 23212 21756 23268
rect 21812 23212 21822 23268
rect 23538 23212 23548 23268
rect 23604 23212 27020 23268
rect 27076 23212 27086 23268
rect 28476 23212 37324 23268
rect 37380 23212 37390 23268
rect 0 22932 800 22960
rect 8372 22932 8428 23212
rect 28476 23156 28532 23212
rect 13122 23100 13132 23156
rect 13188 23100 13804 23156
rect 13860 23100 15596 23156
rect 15652 23100 15662 23156
rect 28466 23100 28476 23156
rect 28532 23100 28542 23156
rect 28802 23100 28812 23156
rect 28868 23100 37548 23156
rect 37604 23100 37614 23156
rect 25442 22988 25452 23044
rect 25508 22988 38332 23044
rect 38388 22988 38398 23044
rect 39200 22932 40000 22960
rect 0 22876 1708 22932
rect 1764 22876 2492 22932
rect 2548 22876 2558 22932
rect 8372 22876 17612 22932
rect 17668 22876 17678 22932
rect 27682 22876 27692 22932
rect 27748 22876 28812 22932
rect 28868 22876 28878 22932
rect 37650 22876 37660 22932
rect 37716 22876 38220 22932
rect 38276 22876 40000 22932
rect 0 22848 800 22876
rect 39200 22848 40000 22876
rect 5864 22708 5874 22764
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 6138 22708 6148 22764
rect 15188 22708 15198 22764
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15462 22708 15472 22764
rect 24512 22708 24522 22764
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24786 22708 24796 22764
rect 33836 22708 33846 22764
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 34110 22708 34120 22764
rect 15026 22428 15036 22484
rect 15092 22428 16828 22484
rect 16884 22428 17388 22484
rect 17444 22428 19068 22484
rect 19124 22428 19628 22484
rect 19684 22428 19694 22484
rect 2034 22316 2044 22372
rect 2100 22316 15932 22372
rect 15988 22316 15998 22372
rect 0 22260 800 22288
rect 39200 22260 40000 22288
rect 0 22204 1708 22260
rect 1764 22204 2492 22260
rect 2548 22204 2558 22260
rect 21970 22204 21980 22260
rect 22036 22204 25788 22260
rect 25844 22204 25854 22260
rect 36530 22204 36540 22260
rect 36596 22204 38220 22260
rect 38276 22204 40000 22260
rect 0 22176 800 22204
rect 39200 22176 40000 22204
rect 13570 22092 13580 22148
rect 13636 22092 19516 22148
rect 19572 22092 20636 22148
rect 20692 22092 20860 22148
rect 20916 22092 20926 22148
rect 21522 22092 21532 22148
rect 21588 22092 22204 22148
rect 22260 22092 22270 22148
rect 10526 21924 10536 21980
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10800 21924 10810 21980
rect 19850 21924 19860 21980
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 20124 21924 20134 21980
rect 29174 21924 29184 21980
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29448 21924 29458 21980
rect 38498 21924 38508 21980
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38772 21924 38782 21980
rect 2034 21644 2044 21700
rect 2100 21644 12236 21700
rect 12292 21644 12302 21700
rect 14466 21644 14476 21700
rect 14532 21644 15820 21700
rect 15876 21644 15886 21700
rect 18498 21644 18508 21700
rect 18564 21644 20412 21700
rect 20468 21644 20478 21700
rect 0 21588 800 21616
rect 39200 21588 40000 21616
rect 0 21532 2380 21588
rect 2436 21532 3164 21588
rect 3220 21532 3230 21588
rect 37538 21532 37548 21588
rect 37604 21532 40000 21588
rect 0 21504 800 21532
rect 39200 21504 40000 21532
rect 1698 21420 1708 21476
rect 1764 21420 2940 21476
rect 2996 21420 3006 21476
rect 17938 21420 17948 21476
rect 18004 21420 18956 21476
rect 19012 21420 19022 21476
rect 20066 21420 20076 21476
rect 20132 21420 20300 21476
rect 20356 21420 20366 21476
rect 23202 21420 23212 21476
rect 23268 21420 23436 21476
rect 23492 21420 23772 21476
rect 23828 21420 23838 21476
rect 24434 21420 24444 21476
rect 24500 21420 25004 21476
rect 25060 21420 25070 21476
rect 37202 21420 37212 21476
rect 37268 21420 38220 21476
rect 38276 21420 38286 21476
rect 2594 21308 2604 21364
rect 2660 21308 12124 21364
rect 12180 21308 15372 21364
rect 15428 21308 15438 21364
rect 5864 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6148 21196
rect 15188 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15472 21196
rect 24512 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24796 21196
rect 33836 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34120 21196
rect 12898 20972 12908 21028
rect 12964 20972 16268 21028
rect 16324 20972 18508 21028
rect 18564 20972 18574 21028
rect 23762 20972 23772 21028
rect 23828 20972 24332 21028
rect 24388 20972 28252 21028
rect 28308 20972 37100 21028
rect 37156 20972 37166 21028
rect 0 20916 800 20944
rect 39200 20916 40000 20944
rect 0 20860 1708 20916
rect 1764 20860 1774 20916
rect 2818 20860 2828 20916
rect 2884 20860 8428 20916
rect 12450 20860 12460 20916
rect 12516 20860 13580 20916
rect 13636 20860 13646 20916
rect 15810 20860 15820 20916
rect 15876 20860 16940 20916
rect 16996 20860 17006 20916
rect 27132 20860 37996 20916
rect 38052 20860 38062 20916
rect 38210 20860 38220 20916
rect 38276 20860 40000 20916
rect 0 20832 800 20860
rect 8372 20804 8428 20860
rect 27132 20804 27188 20860
rect 39200 20832 40000 20860
rect 8372 20748 11340 20804
rect 11396 20748 13468 20804
rect 13524 20748 13534 20804
rect 20178 20748 20188 20804
rect 20244 20748 21196 20804
rect 21252 20748 21262 20804
rect 24434 20748 24444 20804
rect 24500 20748 25004 20804
rect 25060 20748 25564 20804
rect 25620 20748 25630 20804
rect 27122 20748 27132 20804
rect 27188 20748 27198 20804
rect 27356 20748 37884 20804
rect 37940 20748 37950 20804
rect 27356 20692 27412 20748
rect 8372 20636 11788 20692
rect 11844 20636 16828 20692
rect 16884 20636 16894 20692
rect 18274 20636 18284 20692
rect 18340 20636 21420 20692
rect 21476 20636 21486 20692
rect 23090 20636 23100 20692
rect 23156 20636 23166 20692
rect 23426 20636 23436 20692
rect 23492 20636 27412 20692
rect 27794 20636 27804 20692
rect 27860 20636 38892 20692
rect 38948 20636 38958 20692
rect 8372 20580 8428 20636
rect 23100 20580 23156 20636
rect 27804 20580 27860 20636
rect 2258 20524 2268 20580
rect 2324 20524 8428 20580
rect 18610 20524 18620 20580
rect 18676 20524 23156 20580
rect 23986 20524 23996 20580
rect 24052 20524 27860 20580
rect 27916 20524 29652 20580
rect 27916 20468 27972 20524
rect 24882 20412 24892 20468
rect 24948 20412 25396 20468
rect 25554 20412 25564 20468
rect 25620 20412 25788 20468
rect 25844 20412 27972 20468
rect 10526 20356 10536 20412
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10800 20356 10810 20412
rect 19850 20356 19860 20412
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 20124 20356 20134 20412
rect 22754 20300 22764 20356
rect 22820 20300 25004 20356
rect 25060 20300 25070 20356
rect 0 20244 800 20272
rect 25340 20244 25396 20412
rect 29174 20356 29184 20412
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29448 20356 29458 20412
rect 29596 20356 29652 20524
rect 31892 20524 37884 20580
rect 37940 20524 37950 20580
rect 31892 20468 31948 20524
rect 29922 20412 29932 20468
rect 29988 20412 31948 20468
rect 38498 20356 38508 20412
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38772 20356 38782 20412
rect 29596 20300 37436 20356
rect 37492 20300 37502 20356
rect 39200 20244 40000 20272
rect 0 20188 1708 20244
rect 1764 20188 2492 20244
rect 2548 20188 2558 20244
rect 19954 20188 19964 20244
rect 20020 20188 20972 20244
rect 21028 20188 21038 20244
rect 25330 20188 25340 20244
rect 25396 20188 29932 20244
rect 29988 20188 29998 20244
rect 37650 20188 37660 20244
rect 37716 20188 38220 20244
rect 38276 20188 40000 20244
rect 0 20160 800 20188
rect 21746 20132 21756 20188
rect 21812 20132 21832 20188
rect 39200 20160 40000 20188
rect 2034 20076 2044 20132
rect 2100 20076 12236 20132
rect 12292 20076 12302 20132
rect 19730 20076 19740 20132
rect 19796 20076 20300 20132
rect 20356 20076 22876 20132
rect 22932 20076 22942 20132
rect 23202 20076 23212 20132
rect 23268 20076 24220 20132
rect 24276 20076 24286 20132
rect 36978 20076 36988 20132
rect 37044 20076 37884 20132
rect 37940 20076 37950 20132
rect 8372 19964 15372 20020
rect 15428 19964 15438 20020
rect 21634 19964 21644 20020
rect 21700 19964 22764 20020
rect 22820 19964 22830 20020
rect 23996 19964 26908 20020
rect 26964 19964 26974 20020
rect 29922 19964 29932 20020
rect 29988 19964 37324 20020
rect 37380 19964 37390 20020
rect 8372 19796 8428 19964
rect 23996 19908 24052 19964
rect 21858 19852 21868 19908
rect 21924 19852 23324 19908
rect 23380 19852 23996 19908
rect 24052 19852 24062 19908
rect 26562 19852 26572 19908
rect 26628 19852 37548 19908
rect 37604 19852 37614 19908
rect 2146 19740 2156 19796
rect 2212 19740 8428 19796
rect 21522 19740 21532 19796
rect 21588 19740 23548 19796
rect 23604 19740 24668 19796
rect 24724 19740 24734 19796
rect 25218 19740 25228 19796
rect 25284 19740 26236 19796
rect 26292 19740 28476 19796
rect 28532 19740 28542 19796
rect 0 19572 800 19600
rect 5864 19572 5874 19628
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 6138 19572 6148 19628
rect 15188 19572 15198 19628
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15462 19572 15472 19628
rect 24512 19572 24522 19628
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24786 19572 24796 19628
rect 33836 19572 33846 19628
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 34110 19572 34120 19628
rect 39200 19572 40000 19600
rect 0 19516 1708 19572
rect 1764 19516 2492 19572
rect 2548 19516 2558 19572
rect 21634 19516 21644 19572
rect 21700 19516 21868 19572
rect 21924 19516 21934 19572
rect 22082 19516 22092 19572
rect 22148 19516 24388 19572
rect 38210 19516 38220 19572
rect 38276 19516 40000 19572
rect 0 19488 800 19516
rect 24332 19460 24388 19516
rect 39200 19488 40000 19516
rect 12898 19404 12908 19460
rect 12964 19404 19292 19460
rect 19348 19404 19358 19460
rect 24332 19404 27692 19460
rect 27748 19404 27758 19460
rect 2706 19292 2716 19348
rect 2772 19292 13524 19348
rect 20402 19292 20412 19348
rect 20468 19292 20860 19348
rect 20916 19292 25228 19348
rect 25284 19292 25294 19348
rect 26236 19292 37884 19348
rect 37940 19292 37950 19348
rect 13468 19236 13524 19292
rect 26236 19236 26292 19292
rect 4274 19180 4284 19236
rect 4340 19180 8428 19236
rect 13458 19180 13468 19236
rect 13524 19180 13534 19236
rect 17724 19180 18732 19236
rect 18788 19180 18798 19236
rect 19618 19180 19628 19236
rect 19684 19180 21084 19236
rect 21140 19180 21150 19236
rect 26226 19180 26236 19236
rect 26292 19180 26302 19236
rect 27570 19180 27580 19236
rect 27636 19180 36988 19236
rect 37044 19180 37054 19236
rect 8372 19124 8428 19180
rect 17724 19124 17780 19180
rect 8372 19068 17780 19124
rect 18498 19068 18508 19124
rect 18564 19068 26348 19124
rect 26404 19068 26414 19124
rect 27458 18956 27468 19012
rect 27524 18956 28476 19012
rect 28532 18956 31948 19012
rect 37650 18956 37660 19012
rect 37716 18956 38220 19012
rect 38276 18956 38948 19012
rect 0 18900 800 18928
rect 31892 18900 31948 18956
rect 38892 18900 38948 18956
rect 39200 18900 40000 18928
rect 0 18844 1932 18900
rect 1988 18844 1998 18900
rect 31892 18844 37772 18900
rect 37828 18844 37838 18900
rect 38892 18844 40000 18900
rect 0 18816 800 18844
rect 10526 18788 10536 18844
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10800 18788 10810 18844
rect 19850 18788 19860 18844
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 20124 18788 20134 18844
rect 29174 18788 29184 18844
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29448 18788 29458 18844
rect 38498 18788 38508 18844
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38772 18788 38782 18844
rect 39200 18816 40000 18844
rect 14914 18620 14924 18676
rect 14980 18620 19180 18676
rect 19236 18620 19246 18676
rect 20132 18620 23212 18676
rect 23268 18620 23278 18676
rect 20132 18564 20188 18620
rect 18610 18508 18620 18564
rect 18676 18508 19740 18564
rect 19796 18508 20188 18564
rect 2034 18396 2044 18452
rect 2100 18396 16828 18452
rect 16884 18396 16894 18452
rect 18946 18396 18956 18452
rect 19012 18396 20412 18452
rect 20468 18396 20478 18452
rect 21522 18396 21532 18452
rect 21588 18396 22876 18452
rect 22932 18396 22942 18452
rect 13010 18284 13020 18340
rect 13076 18284 14924 18340
rect 14980 18284 15820 18340
rect 15876 18284 17388 18340
rect 17444 18284 17454 18340
rect 22530 18284 22540 18340
rect 22596 18284 22988 18340
rect 23044 18284 37884 18340
rect 37940 18284 37950 18340
rect 0 18228 800 18256
rect 39200 18228 40000 18256
rect 0 18172 1708 18228
rect 1764 18172 2492 18228
rect 2548 18172 2558 18228
rect 12562 18172 12572 18228
rect 12628 18172 19292 18228
rect 19348 18172 19358 18228
rect 37650 18172 37660 18228
rect 37716 18172 38220 18228
rect 38276 18172 40000 18228
rect 0 18144 800 18172
rect 39200 18144 40000 18172
rect 5864 18004 5874 18060
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 6138 18004 6148 18060
rect 15188 18004 15198 18060
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15462 18004 15472 18060
rect 24512 18004 24522 18060
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24786 18004 24796 18060
rect 33836 18004 33846 18060
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 34110 18004 34120 18060
rect 12786 17836 12796 17892
rect 12852 17836 13468 17892
rect 13524 17836 13534 17892
rect 16258 17836 16268 17892
rect 16324 17836 19628 17892
rect 19684 17836 19694 17892
rect 1922 17724 1932 17780
rect 1988 17724 1998 17780
rect 2146 17724 2156 17780
rect 2212 17724 13804 17780
rect 13860 17724 13870 17780
rect 0 17556 800 17584
rect 1932 17556 1988 17724
rect 2706 17612 2716 17668
rect 2772 17612 11788 17668
rect 11844 17612 11854 17668
rect 12226 17612 12236 17668
rect 12292 17612 14028 17668
rect 14084 17612 14094 17668
rect 19954 17612 19964 17668
rect 20020 17612 26348 17668
rect 26404 17612 26414 17668
rect 39200 17556 40000 17584
rect 0 17500 1988 17556
rect 18498 17500 18508 17556
rect 18564 17500 19068 17556
rect 19124 17500 19852 17556
rect 19908 17500 20412 17556
rect 20468 17500 20478 17556
rect 25330 17500 25340 17556
rect 25396 17500 29260 17556
rect 29316 17500 29596 17556
rect 29652 17500 29662 17556
rect 36530 17500 36540 17556
rect 36596 17500 38220 17556
rect 38276 17500 40000 17556
rect 0 17472 800 17500
rect 39200 17472 40000 17500
rect 16258 17388 16268 17444
rect 16324 17388 20188 17444
rect 20244 17388 20254 17444
rect 22194 17388 22204 17444
rect 22260 17388 22652 17444
rect 22708 17388 23884 17444
rect 23940 17388 23950 17444
rect 24210 17388 24220 17444
rect 24276 17388 26908 17444
rect 26964 17388 27468 17444
rect 27524 17388 27534 17444
rect 10526 17220 10536 17276
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10800 17220 10810 17276
rect 19850 17220 19860 17276
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 20124 17220 20134 17276
rect 29174 17220 29184 17276
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29448 17220 29458 17276
rect 38498 17220 38508 17276
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38772 17220 38782 17276
rect 20514 17164 20524 17220
rect 20580 17164 26908 17220
rect 26964 17164 26974 17220
rect 18050 17052 18060 17108
rect 18116 17052 19740 17108
rect 19796 17052 19806 17108
rect 20402 17052 20412 17108
rect 20468 17052 21308 17108
rect 21364 17052 21374 17108
rect 22082 17052 22092 17108
rect 22148 17052 22988 17108
rect 23044 17052 23054 17108
rect 23650 17052 23660 17108
rect 23716 17052 37212 17108
rect 37268 17052 37278 17108
rect 18498 16940 18508 16996
rect 18564 16940 22428 16996
rect 22484 16940 22494 16996
rect 29586 16940 29596 16996
rect 29652 16940 37324 16996
rect 37380 16940 37390 16996
rect 37538 16940 37548 16996
rect 37604 16940 38500 16996
rect 0 16884 800 16912
rect 38444 16884 38500 16940
rect 39200 16884 40000 16912
rect 0 16828 1708 16884
rect 1764 16828 2492 16884
rect 2548 16828 2558 16884
rect 13122 16828 13132 16884
rect 13188 16828 14700 16884
rect 14756 16828 14766 16884
rect 19170 16828 19180 16884
rect 19236 16828 19964 16884
rect 20020 16828 20030 16884
rect 23090 16828 23100 16884
rect 23156 16828 24220 16884
rect 24276 16828 24286 16884
rect 37202 16828 37212 16884
rect 37268 16828 38220 16884
rect 38276 16828 38286 16884
rect 38444 16828 40000 16884
rect 0 16800 800 16828
rect 39200 16800 40000 16828
rect 2370 16716 2380 16772
rect 2436 16716 3164 16772
rect 3220 16716 3230 16772
rect 3388 16716 12460 16772
rect 12516 16716 12526 16772
rect 17938 16716 17948 16772
rect 18004 16716 18956 16772
rect 19012 16716 19022 16772
rect 19282 16716 19292 16772
rect 19348 16716 21980 16772
rect 22036 16716 22046 16772
rect 22306 16716 22316 16772
rect 22372 16716 37884 16772
rect 37940 16716 37950 16772
rect 3388 16660 3444 16716
rect 2258 16604 2268 16660
rect 2324 16604 3444 16660
rect 4274 16604 4284 16660
rect 4340 16604 13916 16660
rect 13972 16604 13982 16660
rect 5864 16436 5874 16492
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 6138 16436 6148 16492
rect 15188 16436 15198 16492
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15462 16436 15472 16492
rect 24512 16436 24522 16492
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24786 16436 24796 16492
rect 33836 16436 33846 16492
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 34110 16436 34120 16492
rect 12786 16380 12796 16436
rect 12852 16380 14140 16436
rect 14196 16380 14206 16436
rect 18722 16380 18732 16436
rect 18788 16380 19068 16436
rect 19124 16380 19516 16436
rect 19572 16380 20188 16436
rect 20132 16324 20188 16380
rect 2034 16268 2044 16324
rect 2100 16268 8428 16324
rect 20132 16268 21644 16324
rect 21700 16268 21710 16324
rect 0 16212 800 16240
rect 8372 16212 8428 16268
rect 39200 16212 40000 16240
rect 0 16156 2380 16212
rect 2436 16156 2446 16212
rect 8372 16156 13804 16212
rect 13860 16156 13870 16212
rect 38210 16156 38220 16212
rect 38276 16156 40000 16212
rect 0 16128 800 16156
rect 39200 16128 40000 16156
rect 14242 16044 14252 16100
rect 14308 16044 15148 16100
rect 15204 16044 17388 16100
rect 17444 16044 17454 16100
rect 17938 16044 17948 16100
rect 18004 16044 18284 16100
rect 18340 16044 19740 16100
rect 19796 16044 19806 16100
rect 2034 15820 2044 15876
rect 2100 15820 15372 15876
rect 15428 15820 15438 15876
rect 18946 15820 18956 15876
rect 19012 15820 19516 15876
rect 19572 15820 19582 15876
rect 26786 15820 26796 15876
rect 26852 15820 37884 15876
rect 37940 15820 37950 15876
rect 10526 15652 10536 15708
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10800 15652 10810 15708
rect 19850 15652 19860 15708
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 20124 15652 20134 15708
rect 29174 15652 29184 15708
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29448 15652 29458 15708
rect 38498 15652 38508 15708
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38772 15652 38782 15708
rect 0 15540 800 15568
rect 39200 15540 40000 15568
rect 0 15484 1708 15540
rect 1764 15484 2940 15540
rect 2996 15484 3006 15540
rect 37650 15484 37660 15540
rect 37716 15484 38220 15540
rect 38276 15484 40000 15540
rect 0 15456 800 15484
rect 39200 15456 40000 15484
rect 2034 15372 2044 15428
rect 2100 15372 8428 15428
rect 14130 15372 14140 15428
rect 14196 15372 16100 15428
rect 8372 15316 8428 15372
rect 16044 15316 16100 15372
rect 19180 15372 21196 15428
rect 21252 15372 21262 15428
rect 26338 15372 26348 15428
rect 26404 15372 37884 15428
rect 37940 15372 37950 15428
rect 19180 15316 19236 15372
rect 8372 15260 14028 15316
rect 14084 15260 14094 15316
rect 16034 15260 16044 15316
rect 16100 15260 18060 15316
rect 18116 15260 18126 15316
rect 18610 15260 18620 15316
rect 18676 15260 19180 15316
rect 19236 15260 19246 15316
rect 20066 15260 20076 15316
rect 20132 15260 21532 15316
rect 21588 15260 21598 15316
rect 20178 15148 20188 15204
rect 20244 15148 20300 15204
rect 20356 15148 20366 15204
rect 18610 14924 18620 14980
rect 18676 14924 19292 14980
rect 19348 14924 19358 14980
rect 0 14868 800 14896
rect 5864 14868 5874 14924
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 6138 14868 6148 14924
rect 15188 14868 15198 14924
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15462 14868 15472 14924
rect 24512 14868 24522 14924
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24786 14868 24796 14924
rect 33836 14868 33846 14924
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 34110 14868 34120 14924
rect 39200 14868 40000 14896
rect 0 14812 1708 14868
rect 1764 14812 2492 14868
rect 2548 14812 2558 14868
rect 19394 14812 19404 14868
rect 19460 14812 21308 14868
rect 21364 14812 21374 14868
rect 38210 14812 38220 14868
rect 38276 14812 40000 14868
rect 0 14784 800 14812
rect 39200 14784 40000 14812
rect 20598 14700 20636 14756
rect 20692 14700 20702 14756
rect 20178 14588 20188 14644
rect 20244 14588 21420 14644
rect 21476 14588 21486 14644
rect 18050 14476 18060 14532
rect 18116 14476 20412 14532
rect 20468 14476 20478 14532
rect 20626 14476 20636 14532
rect 20692 14476 21532 14532
rect 21588 14476 21598 14532
rect 24994 14476 25004 14532
rect 25060 14476 31052 14532
rect 31108 14476 31118 14532
rect 19618 14364 19628 14420
rect 19684 14364 19964 14420
rect 20020 14364 21420 14420
rect 21476 14364 21486 14420
rect 37650 14364 37660 14420
rect 37716 14364 38276 14420
rect 38220 14308 38276 14364
rect 15810 14252 15820 14308
rect 15876 14252 20412 14308
rect 20468 14252 20478 14308
rect 21186 14252 21196 14308
rect 21252 14252 23772 14308
rect 23828 14252 23838 14308
rect 29026 14252 29036 14308
rect 29092 14252 37884 14308
rect 37940 14252 37950 14308
rect 38210 14252 38220 14308
rect 38276 14252 38948 14308
rect 0 14196 800 14224
rect 38892 14196 38948 14252
rect 39200 14196 40000 14224
rect 0 14140 1708 14196
rect 1764 14140 2492 14196
rect 2548 14140 2558 14196
rect 38892 14140 40000 14196
rect 0 14112 800 14140
rect 10526 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10810 14140
rect 19850 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20134 14140
rect 29174 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29458 14140
rect 38498 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38782 14140
rect 39200 14112 40000 14140
rect 17938 13916 17948 13972
rect 18004 13916 22204 13972
rect 22260 13916 22270 13972
rect 24882 13916 24892 13972
rect 24948 13916 37884 13972
rect 37940 13916 37950 13972
rect 2706 13804 2716 13860
rect 2772 13804 15708 13860
rect 15764 13804 15774 13860
rect 22082 13804 22092 13860
rect 22148 13804 22876 13860
rect 22932 13804 24220 13860
rect 24276 13804 24286 13860
rect 20514 13692 20524 13748
rect 20580 13692 20972 13748
rect 21028 13692 21038 13748
rect 22194 13692 22204 13748
rect 22260 13692 25452 13748
rect 25508 13692 26908 13748
rect 26852 13636 26908 13692
rect 18274 13580 18284 13636
rect 18340 13580 18956 13636
rect 19012 13580 19022 13636
rect 20626 13580 20636 13636
rect 20692 13580 21084 13636
rect 21140 13580 21150 13636
rect 26852 13580 30380 13636
rect 30436 13580 30446 13636
rect 0 13524 800 13552
rect 39200 13524 40000 13552
rect 0 13468 1708 13524
rect 1764 13468 3612 13524
rect 3668 13468 3678 13524
rect 18498 13468 18508 13524
rect 18564 13468 20300 13524
rect 20356 13468 21308 13524
rect 21364 13468 21374 13524
rect 37650 13468 37660 13524
rect 37716 13468 38220 13524
rect 38276 13468 40000 13524
rect 0 13440 800 13468
rect 39200 13440 40000 13468
rect 2370 13356 2380 13412
rect 2436 13356 3164 13412
rect 3220 13356 3230 13412
rect 5864 13300 5874 13356
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 6138 13300 6148 13356
rect 15188 13300 15198 13356
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15462 13300 15472 13356
rect 24512 13300 24522 13356
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24786 13300 24796 13356
rect 33836 13300 33846 13356
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 34110 13300 34120 13356
rect 14690 13132 14700 13188
rect 14756 13132 19292 13188
rect 19348 13132 19358 13188
rect 25890 13132 25900 13188
rect 25956 13132 28252 13188
rect 28308 13132 28318 13188
rect 4274 13020 4284 13076
rect 4340 13020 16828 13076
rect 16884 13020 16894 13076
rect 20066 13020 20076 13076
rect 20132 13020 21644 13076
rect 21700 13020 21710 13076
rect 22754 13020 22764 13076
rect 22820 13020 24332 13076
rect 24388 13020 24398 13076
rect 12674 12908 12684 12964
rect 12740 12908 19292 12964
rect 19348 12908 19358 12964
rect 23762 12908 23772 12964
rect 23828 12908 26572 12964
rect 26628 12908 26638 12964
rect 28130 12908 28140 12964
rect 28196 12908 37884 12964
rect 37940 12908 37950 12964
rect 0 12852 800 12880
rect 39200 12852 40000 12880
rect 0 12796 2380 12852
rect 2436 12796 2446 12852
rect 17826 12796 17836 12852
rect 17892 12796 23828 12852
rect 27346 12796 27356 12852
rect 27412 12796 37212 12852
rect 37268 12796 37278 12852
rect 38210 12796 38220 12852
rect 38276 12796 40000 12852
rect 0 12768 800 12796
rect 23772 12740 23828 12796
rect 38220 12740 38276 12796
rect 39200 12768 40000 12796
rect 18946 12684 18956 12740
rect 19012 12684 20748 12740
rect 20804 12684 20814 12740
rect 20962 12684 20972 12740
rect 21028 12684 21756 12740
rect 21812 12684 21822 12740
rect 23762 12684 23772 12740
rect 23828 12684 23838 12740
rect 36530 12684 36540 12740
rect 36596 12684 38276 12740
rect 10526 12516 10536 12572
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10800 12516 10810 12572
rect 19850 12516 19860 12572
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 20124 12516 20134 12572
rect 29174 12516 29184 12572
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29448 12516 29458 12572
rect 38498 12516 38508 12572
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38772 12516 38782 12572
rect 18946 12348 18956 12404
rect 19012 12348 21532 12404
rect 21588 12348 21598 12404
rect 26002 12236 26012 12292
rect 26068 12236 37884 12292
rect 37940 12236 37950 12292
rect 0 12180 800 12208
rect 39200 12180 40000 12208
rect 0 12124 1932 12180
rect 1988 12124 1998 12180
rect 4274 12124 4284 12180
rect 4340 12124 15932 12180
rect 15988 12124 15998 12180
rect 37538 12124 37548 12180
rect 37604 12124 40000 12180
rect 0 12096 800 12124
rect 39200 12096 40000 12124
rect 37202 12012 37212 12068
rect 37268 12012 38220 12068
rect 38276 12012 38286 12068
rect 18050 11788 18060 11844
rect 18116 11788 18732 11844
rect 18788 11788 18798 11844
rect 5864 11732 5874 11788
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 6138 11732 6148 11788
rect 15188 11732 15198 11788
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15462 11732 15472 11788
rect 24512 11732 24522 11788
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24786 11732 24796 11788
rect 33836 11732 33846 11788
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 34110 11732 34120 11788
rect 0 11508 800 11536
rect 39200 11508 40000 11536
rect 0 11452 1932 11508
rect 1988 11452 1998 11508
rect 38210 11452 38220 11508
rect 38276 11452 40000 11508
rect 0 11424 800 11452
rect 39200 11424 40000 11452
rect 20066 11116 20076 11172
rect 20132 11116 21084 11172
rect 21140 11116 21150 11172
rect 10526 10948 10536 11004
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10800 10948 10810 11004
rect 19850 10948 19860 11004
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 20124 10948 20134 11004
rect 29174 10948 29184 11004
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29448 10948 29458 11004
rect 38498 10948 38508 11004
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38772 10948 38782 11004
rect 39200 10836 40000 10864
rect 37650 10780 37660 10836
rect 37716 10780 38220 10836
rect 38276 10780 40000 10836
rect 39200 10752 40000 10780
rect 28466 10668 28476 10724
rect 28532 10668 37884 10724
rect 37940 10668 37950 10724
rect 37650 10556 37660 10612
rect 37716 10556 38220 10612
rect 38276 10556 38286 10612
rect 23650 10332 23660 10388
rect 23716 10332 25788 10388
rect 25844 10332 25854 10388
rect 5864 10164 5874 10220
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 6138 10164 6148 10220
rect 15188 10164 15198 10220
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15462 10164 15472 10220
rect 24512 10164 24522 10220
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24786 10164 24796 10220
rect 33836 10164 33846 10220
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 34110 10164 34120 10220
rect 39200 10164 40000 10192
rect 15586 10108 15596 10164
rect 15652 10108 19292 10164
rect 19348 10108 19358 10164
rect 38210 10108 38220 10164
rect 38276 10108 40000 10164
rect 39200 10080 40000 10108
rect 10526 9380 10536 9436
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10800 9380 10810 9436
rect 19850 9380 19860 9436
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 20124 9380 20134 9436
rect 29174 9380 29184 9436
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29448 9380 29458 9436
rect 38498 9380 38508 9436
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38772 9380 38782 9436
rect 5864 8596 5874 8652
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 6138 8596 6148 8652
rect 15188 8596 15198 8652
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15462 8596 15472 8652
rect 24512 8596 24522 8652
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24786 8596 24796 8652
rect 33836 8596 33846 8652
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 34110 8596 34120 8652
rect 10526 7812 10536 7868
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10800 7812 10810 7868
rect 19850 7812 19860 7868
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 20124 7812 20134 7868
rect 29174 7812 29184 7868
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29448 7812 29458 7868
rect 38498 7812 38508 7868
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38772 7812 38782 7868
rect 5864 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6148 7084
rect 15188 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15472 7084
rect 24512 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24796 7084
rect 33836 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34120 7084
rect 10526 6244 10536 6300
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10800 6244 10810 6300
rect 19850 6244 19860 6300
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 20124 6244 20134 6300
rect 29174 6244 29184 6300
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29448 6244 29458 6300
rect 38498 6244 38508 6300
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38772 6244 38782 6300
rect 5864 5460 5874 5516
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 6138 5460 6148 5516
rect 15188 5460 15198 5516
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15462 5460 15472 5516
rect 24512 5460 24522 5516
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24786 5460 24796 5516
rect 33836 5460 33846 5516
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 34110 5460 34120 5516
rect 14140 5068 14812 5124
rect 14868 5068 14878 5124
rect 14140 4900 14196 5068
rect 22978 4956 22988 5012
rect 23044 4956 25228 5012
rect 25284 4956 25294 5012
rect 25890 4956 25900 5012
rect 25956 4956 29036 5012
rect 29092 4956 29102 5012
rect 14130 4844 14140 4900
rect 14196 4844 14206 4900
rect 21410 4844 21420 4900
rect 21476 4844 23660 4900
rect 23716 4844 23726 4900
rect 10526 4676 10536 4732
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10800 4676 10810 4732
rect 19850 4676 19860 4732
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 20124 4676 20134 4732
rect 29174 4676 29184 4732
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29448 4676 29458 4732
rect 38498 4676 38508 4732
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38772 4676 38782 4732
rect 16370 4620 16380 4676
rect 16436 4620 18620 4676
rect 18676 4620 18686 4676
rect 16034 4508 16044 4564
rect 16100 4508 20636 4564
rect 20692 4508 20702 4564
rect 20850 4508 20860 4564
rect 20916 4508 22428 4564
rect 22484 4508 22494 4564
rect 24882 4508 24892 4564
rect 24948 4508 27132 4564
rect 27188 4508 27198 4564
rect 24994 4396 25004 4452
rect 25060 4396 29708 4452
rect 29764 4396 29774 4452
rect 14914 4284 14924 4340
rect 14980 4284 20300 4340
rect 20356 4284 20366 4340
rect 20850 4284 20860 4340
rect 20916 4284 21532 4340
rect 21588 4284 21980 4340
rect 22036 4284 22046 4340
rect 5864 3892 5874 3948
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 6138 3892 6148 3948
rect 15188 3892 15198 3948
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15462 3892 15472 3948
rect 24512 3892 24522 3948
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24786 3892 24796 3948
rect 33836 3892 33846 3948
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 34110 3892 34120 3948
rect 23538 3724 23548 3780
rect 23604 3724 27244 3780
rect 27300 3724 27310 3780
rect 19506 3612 19516 3668
rect 19572 3612 20972 3668
rect 21028 3612 21038 3668
rect 18162 3500 18172 3556
rect 18228 3500 18620 3556
rect 18676 3500 18686 3556
rect 24882 3500 24892 3556
rect 24948 3500 25452 3556
rect 25508 3500 25518 3556
rect 26114 3500 26124 3556
rect 26180 3500 27468 3556
rect 27524 3500 27916 3556
rect 27972 3500 27982 3556
rect 28130 3500 28140 3556
rect 28196 3500 28812 3556
rect 28868 3500 29428 3556
rect 29372 3444 29428 3500
rect 12338 3388 12348 3444
rect 12404 3388 13468 3444
rect 13524 3388 13534 3444
rect 17378 3388 17388 3444
rect 17444 3388 20300 3444
rect 20356 3388 20366 3444
rect 22978 3388 22988 3444
rect 23044 3388 23436 3444
rect 23492 3388 23884 3444
rect 23940 3388 23950 3444
rect 24994 3388 25004 3444
rect 25060 3388 26348 3444
rect 26404 3388 26414 3444
rect 27682 3388 27692 3444
rect 27748 3388 28588 3444
rect 28644 3388 28654 3444
rect 29362 3388 29372 3444
rect 29428 3388 29438 3444
rect 29586 3388 29596 3444
rect 29652 3388 30156 3444
rect 30212 3388 30604 3444
rect 30660 3388 30670 3444
rect 10526 3108 10536 3164
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10800 3108 10810 3164
rect 19850 3108 19860 3164
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 20124 3108 20134 3164
rect 29174 3108 29184 3164
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29448 3108 29458 3164
rect 38498 3108 38508 3164
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38772 3108 38782 3164
<< via3 >>
rect 5874 36820 5930 36876
rect 5978 36820 6034 36876
rect 6082 36820 6138 36876
rect 15198 36820 15254 36876
rect 15302 36820 15358 36876
rect 15406 36820 15462 36876
rect 24522 36820 24578 36876
rect 24626 36820 24682 36876
rect 24730 36820 24786 36876
rect 33846 36820 33902 36876
rect 33950 36820 34006 36876
rect 34054 36820 34110 36876
rect 10536 36036 10592 36092
rect 10640 36036 10696 36092
rect 10744 36036 10800 36092
rect 19860 36036 19916 36092
rect 19964 36036 20020 36092
rect 20068 36036 20124 36092
rect 29184 36036 29240 36092
rect 29288 36036 29344 36092
rect 29392 36036 29448 36092
rect 38508 36036 38564 36092
rect 38612 36036 38668 36092
rect 38716 36036 38772 36092
rect 5874 35252 5930 35308
rect 5978 35252 6034 35308
rect 6082 35252 6138 35308
rect 15198 35252 15254 35308
rect 15302 35252 15358 35308
rect 15406 35252 15462 35308
rect 24522 35252 24578 35308
rect 24626 35252 24682 35308
rect 24730 35252 24786 35308
rect 33846 35252 33902 35308
rect 33950 35252 34006 35308
rect 34054 35252 34110 35308
rect 10536 34468 10592 34524
rect 10640 34468 10696 34524
rect 10744 34468 10800 34524
rect 19860 34468 19916 34524
rect 19964 34468 20020 34524
rect 20068 34468 20124 34524
rect 29184 34468 29240 34524
rect 29288 34468 29344 34524
rect 29392 34468 29448 34524
rect 38508 34468 38564 34524
rect 38612 34468 38668 34524
rect 38716 34468 38772 34524
rect 5874 33684 5930 33740
rect 5978 33684 6034 33740
rect 6082 33684 6138 33740
rect 15198 33684 15254 33740
rect 15302 33684 15358 33740
rect 15406 33684 15462 33740
rect 24522 33684 24578 33740
rect 24626 33684 24682 33740
rect 24730 33684 24786 33740
rect 33846 33684 33902 33740
rect 33950 33684 34006 33740
rect 34054 33684 34110 33740
rect 10536 32900 10592 32956
rect 10640 32900 10696 32956
rect 10744 32900 10800 32956
rect 19860 32900 19916 32956
rect 19964 32900 20020 32956
rect 20068 32900 20124 32956
rect 29184 32900 29240 32956
rect 29288 32900 29344 32956
rect 29392 32900 29448 32956
rect 38508 32900 38564 32956
rect 38612 32900 38668 32956
rect 38716 32900 38772 32956
rect 5874 32116 5930 32172
rect 5978 32116 6034 32172
rect 6082 32116 6138 32172
rect 15198 32116 15254 32172
rect 15302 32116 15358 32172
rect 15406 32116 15462 32172
rect 24522 32116 24578 32172
rect 24626 32116 24682 32172
rect 24730 32116 24786 32172
rect 33846 32116 33902 32172
rect 33950 32116 34006 32172
rect 34054 32116 34110 32172
rect 10536 31332 10592 31388
rect 10640 31332 10696 31388
rect 10744 31332 10800 31388
rect 19860 31332 19916 31388
rect 19964 31332 20020 31388
rect 20068 31332 20124 31388
rect 29184 31332 29240 31388
rect 29288 31332 29344 31388
rect 29392 31332 29448 31388
rect 38508 31332 38564 31388
rect 38612 31332 38668 31388
rect 38716 31332 38772 31388
rect 5874 30548 5930 30604
rect 5978 30548 6034 30604
rect 6082 30548 6138 30604
rect 15198 30548 15254 30604
rect 15302 30548 15358 30604
rect 15406 30548 15462 30604
rect 24522 30548 24578 30604
rect 24626 30548 24682 30604
rect 24730 30548 24786 30604
rect 33846 30548 33902 30604
rect 33950 30548 34006 30604
rect 34054 30548 34110 30604
rect 10536 29764 10592 29820
rect 10640 29764 10696 29820
rect 10744 29764 10800 29820
rect 19860 29764 19916 29820
rect 19964 29764 20020 29820
rect 20068 29764 20124 29820
rect 29184 29764 29240 29820
rect 29288 29764 29344 29820
rect 29392 29764 29448 29820
rect 38508 29764 38564 29820
rect 38612 29764 38668 29820
rect 38716 29764 38772 29820
rect 5874 28980 5930 29036
rect 5978 28980 6034 29036
rect 6082 28980 6138 29036
rect 15198 28980 15254 29036
rect 15302 28980 15358 29036
rect 15406 28980 15462 29036
rect 24522 28980 24578 29036
rect 24626 28980 24682 29036
rect 24730 28980 24786 29036
rect 33846 28980 33902 29036
rect 33950 28980 34006 29036
rect 34054 28980 34110 29036
rect 10536 28196 10592 28252
rect 10640 28196 10696 28252
rect 10744 28196 10800 28252
rect 19860 28196 19916 28252
rect 19964 28196 20020 28252
rect 20068 28196 20124 28252
rect 29184 28196 29240 28252
rect 29288 28196 29344 28252
rect 29392 28196 29448 28252
rect 38508 28196 38564 28252
rect 38612 28196 38668 28252
rect 38716 28196 38772 28252
rect 5874 27412 5930 27468
rect 5978 27412 6034 27468
rect 6082 27412 6138 27468
rect 15198 27412 15254 27468
rect 15302 27412 15358 27468
rect 15406 27412 15462 27468
rect 24522 27412 24578 27468
rect 24626 27412 24682 27468
rect 24730 27412 24786 27468
rect 33846 27412 33902 27468
rect 33950 27412 34006 27468
rect 34054 27412 34110 27468
rect 10536 26628 10592 26684
rect 10640 26628 10696 26684
rect 10744 26628 10800 26684
rect 19860 26628 19916 26684
rect 19964 26628 20020 26684
rect 20068 26628 20124 26684
rect 29184 26628 29240 26684
rect 29288 26628 29344 26684
rect 29392 26628 29448 26684
rect 38508 26628 38564 26684
rect 38612 26628 38668 26684
rect 38716 26628 38772 26684
rect 5874 25844 5930 25900
rect 5978 25844 6034 25900
rect 6082 25844 6138 25900
rect 15198 25844 15254 25900
rect 15302 25844 15358 25900
rect 15406 25844 15462 25900
rect 24522 25844 24578 25900
rect 24626 25844 24682 25900
rect 24730 25844 24786 25900
rect 33846 25844 33902 25900
rect 33950 25844 34006 25900
rect 34054 25844 34110 25900
rect 10536 25060 10592 25116
rect 10640 25060 10696 25116
rect 10744 25060 10800 25116
rect 19860 25060 19916 25116
rect 19964 25060 20020 25116
rect 20068 25060 20124 25116
rect 29184 25060 29240 25116
rect 29288 25060 29344 25116
rect 29392 25060 29448 25116
rect 38508 25060 38564 25116
rect 38612 25060 38668 25116
rect 38716 25060 38772 25116
rect 5874 24276 5930 24332
rect 5978 24276 6034 24332
rect 6082 24276 6138 24332
rect 15198 24276 15254 24332
rect 15302 24276 15358 24332
rect 15406 24276 15462 24332
rect 24522 24276 24578 24332
rect 24626 24276 24682 24332
rect 24730 24276 24786 24332
rect 33846 24276 33902 24332
rect 33950 24276 34006 24332
rect 34054 24276 34110 24332
rect 10536 23492 10592 23548
rect 10640 23492 10696 23548
rect 10744 23492 10800 23548
rect 19860 23492 19916 23548
rect 19964 23492 20020 23548
rect 20068 23492 20124 23548
rect 29184 23492 29240 23548
rect 29288 23492 29344 23548
rect 29392 23492 29448 23548
rect 38508 23492 38564 23548
rect 38612 23492 38668 23548
rect 38716 23492 38772 23548
rect 5874 22708 5930 22764
rect 5978 22708 6034 22764
rect 6082 22708 6138 22764
rect 15198 22708 15254 22764
rect 15302 22708 15358 22764
rect 15406 22708 15462 22764
rect 24522 22708 24578 22764
rect 24626 22708 24682 22764
rect 24730 22708 24786 22764
rect 33846 22708 33902 22764
rect 33950 22708 34006 22764
rect 34054 22708 34110 22764
rect 10536 21924 10592 21980
rect 10640 21924 10696 21980
rect 10744 21924 10800 21980
rect 19860 21924 19916 21980
rect 19964 21924 20020 21980
rect 20068 21924 20124 21980
rect 29184 21924 29240 21980
rect 29288 21924 29344 21980
rect 29392 21924 29448 21980
rect 38508 21924 38564 21980
rect 38612 21924 38668 21980
rect 38716 21924 38772 21980
rect 5874 21140 5930 21196
rect 5978 21140 6034 21196
rect 6082 21140 6138 21196
rect 15198 21140 15254 21196
rect 15302 21140 15358 21196
rect 15406 21140 15462 21196
rect 24522 21140 24578 21196
rect 24626 21140 24682 21196
rect 24730 21140 24786 21196
rect 33846 21140 33902 21196
rect 33950 21140 34006 21196
rect 34054 21140 34110 21196
rect 10536 20356 10592 20412
rect 10640 20356 10696 20412
rect 10744 20356 10800 20412
rect 19860 20356 19916 20412
rect 19964 20356 20020 20412
rect 20068 20356 20124 20412
rect 29184 20356 29240 20412
rect 29288 20356 29344 20412
rect 29392 20356 29448 20412
rect 38508 20356 38564 20412
rect 38612 20356 38668 20412
rect 38716 20356 38772 20412
rect 5874 19572 5930 19628
rect 5978 19572 6034 19628
rect 6082 19572 6138 19628
rect 15198 19572 15254 19628
rect 15302 19572 15358 19628
rect 15406 19572 15462 19628
rect 24522 19572 24578 19628
rect 24626 19572 24682 19628
rect 24730 19572 24786 19628
rect 33846 19572 33902 19628
rect 33950 19572 34006 19628
rect 34054 19572 34110 19628
rect 10536 18788 10592 18844
rect 10640 18788 10696 18844
rect 10744 18788 10800 18844
rect 19860 18788 19916 18844
rect 19964 18788 20020 18844
rect 20068 18788 20124 18844
rect 29184 18788 29240 18844
rect 29288 18788 29344 18844
rect 29392 18788 29448 18844
rect 38508 18788 38564 18844
rect 38612 18788 38668 18844
rect 38716 18788 38772 18844
rect 5874 18004 5930 18060
rect 5978 18004 6034 18060
rect 6082 18004 6138 18060
rect 15198 18004 15254 18060
rect 15302 18004 15358 18060
rect 15406 18004 15462 18060
rect 24522 18004 24578 18060
rect 24626 18004 24682 18060
rect 24730 18004 24786 18060
rect 33846 18004 33902 18060
rect 33950 18004 34006 18060
rect 34054 18004 34110 18060
rect 10536 17220 10592 17276
rect 10640 17220 10696 17276
rect 10744 17220 10800 17276
rect 19860 17220 19916 17276
rect 19964 17220 20020 17276
rect 20068 17220 20124 17276
rect 29184 17220 29240 17276
rect 29288 17220 29344 17276
rect 29392 17220 29448 17276
rect 38508 17220 38564 17276
rect 38612 17220 38668 17276
rect 38716 17220 38772 17276
rect 5874 16436 5930 16492
rect 5978 16436 6034 16492
rect 6082 16436 6138 16492
rect 15198 16436 15254 16492
rect 15302 16436 15358 16492
rect 15406 16436 15462 16492
rect 24522 16436 24578 16492
rect 24626 16436 24682 16492
rect 24730 16436 24786 16492
rect 33846 16436 33902 16492
rect 33950 16436 34006 16492
rect 34054 16436 34110 16492
rect 10536 15652 10592 15708
rect 10640 15652 10696 15708
rect 10744 15652 10800 15708
rect 19860 15652 19916 15708
rect 19964 15652 20020 15708
rect 20068 15652 20124 15708
rect 29184 15652 29240 15708
rect 29288 15652 29344 15708
rect 29392 15652 29448 15708
rect 38508 15652 38564 15708
rect 38612 15652 38668 15708
rect 38716 15652 38772 15708
rect 20300 15148 20356 15204
rect 5874 14868 5930 14924
rect 5978 14868 6034 14924
rect 6082 14868 6138 14924
rect 15198 14868 15254 14924
rect 15302 14868 15358 14924
rect 15406 14868 15462 14924
rect 24522 14868 24578 14924
rect 24626 14868 24682 14924
rect 24730 14868 24786 14924
rect 33846 14868 33902 14924
rect 33950 14868 34006 14924
rect 34054 14868 34110 14924
rect 20636 14700 20692 14756
rect 10536 14084 10592 14140
rect 10640 14084 10696 14140
rect 10744 14084 10800 14140
rect 19860 14084 19916 14140
rect 19964 14084 20020 14140
rect 20068 14084 20124 14140
rect 29184 14084 29240 14140
rect 29288 14084 29344 14140
rect 29392 14084 29448 14140
rect 38508 14084 38564 14140
rect 38612 14084 38668 14140
rect 38716 14084 38772 14140
rect 20636 13580 20692 13636
rect 5874 13300 5930 13356
rect 5978 13300 6034 13356
rect 6082 13300 6138 13356
rect 15198 13300 15254 13356
rect 15302 13300 15358 13356
rect 15406 13300 15462 13356
rect 24522 13300 24578 13356
rect 24626 13300 24682 13356
rect 24730 13300 24786 13356
rect 33846 13300 33902 13356
rect 33950 13300 34006 13356
rect 34054 13300 34110 13356
rect 10536 12516 10592 12572
rect 10640 12516 10696 12572
rect 10744 12516 10800 12572
rect 19860 12516 19916 12572
rect 19964 12516 20020 12572
rect 20068 12516 20124 12572
rect 29184 12516 29240 12572
rect 29288 12516 29344 12572
rect 29392 12516 29448 12572
rect 38508 12516 38564 12572
rect 38612 12516 38668 12572
rect 38716 12516 38772 12572
rect 5874 11732 5930 11788
rect 5978 11732 6034 11788
rect 6082 11732 6138 11788
rect 15198 11732 15254 11788
rect 15302 11732 15358 11788
rect 15406 11732 15462 11788
rect 24522 11732 24578 11788
rect 24626 11732 24682 11788
rect 24730 11732 24786 11788
rect 33846 11732 33902 11788
rect 33950 11732 34006 11788
rect 34054 11732 34110 11788
rect 10536 10948 10592 11004
rect 10640 10948 10696 11004
rect 10744 10948 10800 11004
rect 19860 10948 19916 11004
rect 19964 10948 20020 11004
rect 20068 10948 20124 11004
rect 29184 10948 29240 11004
rect 29288 10948 29344 11004
rect 29392 10948 29448 11004
rect 38508 10948 38564 11004
rect 38612 10948 38668 11004
rect 38716 10948 38772 11004
rect 5874 10164 5930 10220
rect 5978 10164 6034 10220
rect 6082 10164 6138 10220
rect 15198 10164 15254 10220
rect 15302 10164 15358 10220
rect 15406 10164 15462 10220
rect 24522 10164 24578 10220
rect 24626 10164 24682 10220
rect 24730 10164 24786 10220
rect 33846 10164 33902 10220
rect 33950 10164 34006 10220
rect 34054 10164 34110 10220
rect 10536 9380 10592 9436
rect 10640 9380 10696 9436
rect 10744 9380 10800 9436
rect 19860 9380 19916 9436
rect 19964 9380 20020 9436
rect 20068 9380 20124 9436
rect 29184 9380 29240 9436
rect 29288 9380 29344 9436
rect 29392 9380 29448 9436
rect 38508 9380 38564 9436
rect 38612 9380 38668 9436
rect 38716 9380 38772 9436
rect 5874 8596 5930 8652
rect 5978 8596 6034 8652
rect 6082 8596 6138 8652
rect 15198 8596 15254 8652
rect 15302 8596 15358 8652
rect 15406 8596 15462 8652
rect 24522 8596 24578 8652
rect 24626 8596 24682 8652
rect 24730 8596 24786 8652
rect 33846 8596 33902 8652
rect 33950 8596 34006 8652
rect 34054 8596 34110 8652
rect 10536 7812 10592 7868
rect 10640 7812 10696 7868
rect 10744 7812 10800 7868
rect 19860 7812 19916 7868
rect 19964 7812 20020 7868
rect 20068 7812 20124 7868
rect 29184 7812 29240 7868
rect 29288 7812 29344 7868
rect 29392 7812 29448 7868
rect 38508 7812 38564 7868
rect 38612 7812 38668 7868
rect 38716 7812 38772 7868
rect 5874 7028 5930 7084
rect 5978 7028 6034 7084
rect 6082 7028 6138 7084
rect 15198 7028 15254 7084
rect 15302 7028 15358 7084
rect 15406 7028 15462 7084
rect 24522 7028 24578 7084
rect 24626 7028 24682 7084
rect 24730 7028 24786 7084
rect 33846 7028 33902 7084
rect 33950 7028 34006 7084
rect 34054 7028 34110 7084
rect 10536 6244 10592 6300
rect 10640 6244 10696 6300
rect 10744 6244 10800 6300
rect 19860 6244 19916 6300
rect 19964 6244 20020 6300
rect 20068 6244 20124 6300
rect 29184 6244 29240 6300
rect 29288 6244 29344 6300
rect 29392 6244 29448 6300
rect 38508 6244 38564 6300
rect 38612 6244 38668 6300
rect 38716 6244 38772 6300
rect 5874 5460 5930 5516
rect 5978 5460 6034 5516
rect 6082 5460 6138 5516
rect 15198 5460 15254 5516
rect 15302 5460 15358 5516
rect 15406 5460 15462 5516
rect 24522 5460 24578 5516
rect 24626 5460 24682 5516
rect 24730 5460 24786 5516
rect 33846 5460 33902 5516
rect 33950 5460 34006 5516
rect 34054 5460 34110 5516
rect 10536 4676 10592 4732
rect 10640 4676 10696 4732
rect 10744 4676 10800 4732
rect 19860 4676 19916 4732
rect 19964 4676 20020 4732
rect 20068 4676 20124 4732
rect 29184 4676 29240 4732
rect 29288 4676 29344 4732
rect 29392 4676 29448 4732
rect 38508 4676 38564 4732
rect 38612 4676 38668 4732
rect 38716 4676 38772 4732
rect 20300 4284 20356 4340
rect 5874 3892 5930 3948
rect 5978 3892 6034 3948
rect 6082 3892 6138 3948
rect 15198 3892 15254 3948
rect 15302 3892 15358 3948
rect 15406 3892 15462 3948
rect 24522 3892 24578 3948
rect 24626 3892 24682 3948
rect 24730 3892 24786 3948
rect 33846 3892 33902 3948
rect 33950 3892 34006 3948
rect 34054 3892 34110 3948
rect 10536 3108 10592 3164
rect 10640 3108 10696 3164
rect 10744 3108 10800 3164
rect 19860 3108 19916 3164
rect 19964 3108 20020 3164
rect 20068 3108 20124 3164
rect 29184 3108 29240 3164
rect 29288 3108 29344 3164
rect 29392 3108 29448 3164
rect 38508 3108 38564 3164
rect 38612 3108 38668 3164
rect 38716 3108 38772 3164
<< metal4 >>
rect 5846 36876 6166 36908
rect 5846 36820 5874 36876
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 6138 36820 6166 36876
rect 5846 35308 6166 36820
rect 5846 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6166 35308
rect 5846 33740 6166 35252
rect 5846 33684 5874 33740
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 6138 33684 6166 33740
rect 5846 32172 6166 33684
rect 5846 32116 5874 32172
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 6138 32116 6166 32172
rect 5846 30604 6166 32116
rect 5846 30548 5874 30604
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 6138 30548 6166 30604
rect 5846 29036 6166 30548
rect 5846 28980 5874 29036
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 6138 28980 6166 29036
rect 5846 27468 6166 28980
rect 5846 27412 5874 27468
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 6138 27412 6166 27468
rect 5846 25900 6166 27412
rect 5846 25844 5874 25900
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 6138 25844 6166 25900
rect 5846 24332 6166 25844
rect 5846 24276 5874 24332
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 6138 24276 6166 24332
rect 5846 22764 6166 24276
rect 5846 22708 5874 22764
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 6138 22708 6166 22764
rect 5846 21196 6166 22708
rect 5846 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6166 21196
rect 5846 19628 6166 21140
rect 5846 19572 5874 19628
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 6138 19572 6166 19628
rect 5846 18060 6166 19572
rect 5846 18004 5874 18060
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 6138 18004 6166 18060
rect 5846 16492 6166 18004
rect 5846 16436 5874 16492
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 6138 16436 6166 16492
rect 5846 14924 6166 16436
rect 5846 14868 5874 14924
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 6138 14868 6166 14924
rect 5846 13356 6166 14868
rect 5846 13300 5874 13356
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 6138 13300 6166 13356
rect 5846 11788 6166 13300
rect 5846 11732 5874 11788
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 6138 11732 6166 11788
rect 5846 10220 6166 11732
rect 5846 10164 5874 10220
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 6138 10164 6166 10220
rect 5846 8652 6166 10164
rect 5846 8596 5874 8652
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 6138 8596 6166 8652
rect 5846 7084 6166 8596
rect 5846 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6166 7084
rect 5846 5516 6166 7028
rect 5846 5460 5874 5516
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 6138 5460 6166 5516
rect 5846 3948 6166 5460
rect 5846 3892 5874 3948
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 6138 3892 6166 3948
rect 5846 3076 6166 3892
rect 10508 36092 10828 36908
rect 10508 36036 10536 36092
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10800 36036 10828 36092
rect 10508 34524 10828 36036
rect 10508 34468 10536 34524
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10800 34468 10828 34524
rect 10508 32956 10828 34468
rect 10508 32900 10536 32956
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10800 32900 10828 32956
rect 10508 31388 10828 32900
rect 10508 31332 10536 31388
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10800 31332 10828 31388
rect 10508 29820 10828 31332
rect 10508 29764 10536 29820
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10800 29764 10828 29820
rect 10508 28252 10828 29764
rect 10508 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10828 28252
rect 10508 26684 10828 28196
rect 10508 26628 10536 26684
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10800 26628 10828 26684
rect 10508 25116 10828 26628
rect 10508 25060 10536 25116
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10800 25060 10828 25116
rect 10508 23548 10828 25060
rect 10508 23492 10536 23548
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10800 23492 10828 23548
rect 10508 21980 10828 23492
rect 10508 21924 10536 21980
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10800 21924 10828 21980
rect 10508 20412 10828 21924
rect 10508 20356 10536 20412
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10800 20356 10828 20412
rect 10508 18844 10828 20356
rect 10508 18788 10536 18844
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10800 18788 10828 18844
rect 10508 17276 10828 18788
rect 10508 17220 10536 17276
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10800 17220 10828 17276
rect 10508 15708 10828 17220
rect 10508 15652 10536 15708
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10800 15652 10828 15708
rect 10508 14140 10828 15652
rect 10508 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10828 14140
rect 10508 12572 10828 14084
rect 10508 12516 10536 12572
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10800 12516 10828 12572
rect 10508 11004 10828 12516
rect 10508 10948 10536 11004
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10800 10948 10828 11004
rect 10508 9436 10828 10948
rect 10508 9380 10536 9436
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10800 9380 10828 9436
rect 10508 7868 10828 9380
rect 10508 7812 10536 7868
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10800 7812 10828 7868
rect 10508 6300 10828 7812
rect 10508 6244 10536 6300
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10800 6244 10828 6300
rect 10508 4732 10828 6244
rect 10508 4676 10536 4732
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10800 4676 10828 4732
rect 10508 3164 10828 4676
rect 10508 3108 10536 3164
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10800 3108 10828 3164
rect 10508 3076 10828 3108
rect 15170 36876 15490 36908
rect 15170 36820 15198 36876
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15462 36820 15490 36876
rect 15170 35308 15490 36820
rect 15170 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15490 35308
rect 15170 33740 15490 35252
rect 15170 33684 15198 33740
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15462 33684 15490 33740
rect 15170 32172 15490 33684
rect 15170 32116 15198 32172
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15462 32116 15490 32172
rect 15170 30604 15490 32116
rect 15170 30548 15198 30604
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15462 30548 15490 30604
rect 15170 29036 15490 30548
rect 15170 28980 15198 29036
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15462 28980 15490 29036
rect 15170 27468 15490 28980
rect 15170 27412 15198 27468
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15462 27412 15490 27468
rect 15170 25900 15490 27412
rect 15170 25844 15198 25900
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15462 25844 15490 25900
rect 15170 24332 15490 25844
rect 15170 24276 15198 24332
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15462 24276 15490 24332
rect 15170 22764 15490 24276
rect 15170 22708 15198 22764
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15462 22708 15490 22764
rect 15170 21196 15490 22708
rect 15170 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15490 21196
rect 15170 19628 15490 21140
rect 15170 19572 15198 19628
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15462 19572 15490 19628
rect 15170 18060 15490 19572
rect 15170 18004 15198 18060
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15462 18004 15490 18060
rect 15170 16492 15490 18004
rect 15170 16436 15198 16492
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15462 16436 15490 16492
rect 15170 14924 15490 16436
rect 15170 14868 15198 14924
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15462 14868 15490 14924
rect 15170 13356 15490 14868
rect 15170 13300 15198 13356
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15462 13300 15490 13356
rect 15170 11788 15490 13300
rect 15170 11732 15198 11788
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15462 11732 15490 11788
rect 15170 10220 15490 11732
rect 15170 10164 15198 10220
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15462 10164 15490 10220
rect 15170 8652 15490 10164
rect 15170 8596 15198 8652
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15462 8596 15490 8652
rect 15170 7084 15490 8596
rect 15170 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15490 7084
rect 15170 5516 15490 7028
rect 15170 5460 15198 5516
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15462 5460 15490 5516
rect 15170 3948 15490 5460
rect 15170 3892 15198 3948
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15462 3892 15490 3948
rect 15170 3076 15490 3892
rect 19832 36092 20152 36908
rect 19832 36036 19860 36092
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 20124 36036 20152 36092
rect 19832 34524 20152 36036
rect 19832 34468 19860 34524
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 20124 34468 20152 34524
rect 19832 32956 20152 34468
rect 19832 32900 19860 32956
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 20124 32900 20152 32956
rect 19832 31388 20152 32900
rect 19832 31332 19860 31388
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 20124 31332 20152 31388
rect 19832 29820 20152 31332
rect 19832 29764 19860 29820
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 20124 29764 20152 29820
rect 19832 28252 20152 29764
rect 19832 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20152 28252
rect 19832 26684 20152 28196
rect 19832 26628 19860 26684
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 20124 26628 20152 26684
rect 19832 25116 20152 26628
rect 19832 25060 19860 25116
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 20124 25060 20152 25116
rect 19832 23548 20152 25060
rect 19832 23492 19860 23548
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 20124 23492 20152 23548
rect 19832 21980 20152 23492
rect 19832 21924 19860 21980
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 20124 21924 20152 21980
rect 19832 20412 20152 21924
rect 19832 20356 19860 20412
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 20124 20356 20152 20412
rect 19832 18844 20152 20356
rect 19832 18788 19860 18844
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 20124 18788 20152 18844
rect 19832 17276 20152 18788
rect 19832 17220 19860 17276
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 20124 17220 20152 17276
rect 19832 15708 20152 17220
rect 19832 15652 19860 15708
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 20124 15652 20152 15708
rect 19832 14140 20152 15652
rect 24494 36876 24814 36908
rect 24494 36820 24522 36876
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24786 36820 24814 36876
rect 24494 35308 24814 36820
rect 24494 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24814 35308
rect 24494 33740 24814 35252
rect 24494 33684 24522 33740
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24786 33684 24814 33740
rect 24494 32172 24814 33684
rect 24494 32116 24522 32172
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24786 32116 24814 32172
rect 24494 30604 24814 32116
rect 24494 30548 24522 30604
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24786 30548 24814 30604
rect 24494 29036 24814 30548
rect 24494 28980 24522 29036
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24786 28980 24814 29036
rect 24494 27468 24814 28980
rect 24494 27412 24522 27468
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24786 27412 24814 27468
rect 24494 25900 24814 27412
rect 24494 25844 24522 25900
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24786 25844 24814 25900
rect 24494 24332 24814 25844
rect 24494 24276 24522 24332
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24786 24276 24814 24332
rect 24494 22764 24814 24276
rect 24494 22708 24522 22764
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24786 22708 24814 22764
rect 24494 21196 24814 22708
rect 24494 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24814 21196
rect 24494 19628 24814 21140
rect 24494 19572 24522 19628
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24786 19572 24814 19628
rect 24494 18060 24814 19572
rect 24494 18004 24522 18060
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24786 18004 24814 18060
rect 24494 16492 24814 18004
rect 24494 16436 24522 16492
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24786 16436 24814 16492
rect 19832 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20152 14140
rect 19832 12572 20152 14084
rect 19832 12516 19860 12572
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 20124 12516 20152 12572
rect 19832 11004 20152 12516
rect 19832 10948 19860 11004
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 20124 10948 20152 11004
rect 19832 9436 20152 10948
rect 19832 9380 19860 9436
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 20124 9380 20152 9436
rect 19832 7868 20152 9380
rect 19832 7812 19860 7868
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 20124 7812 20152 7868
rect 19832 6300 20152 7812
rect 19832 6244 19860 6300
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 20124 6244 20152 6300
rect 19832 4732 20152 6244
rect 19832 4676 19860 4732
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 20124 4676 20152 4732
rect 19832 3164 20152 4676
rect 20300 15204 20356 15214
rect 20300 4340 20356 15148
rect 24494 14924 24814 16436
rect 24494 14868 24522 14924
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24786 14868 24814 14924
rect 20636 14756 20692 14766
rect 20636 13636 20692 14700
rect 20636 13570 20692 13580
rect 20300 4274 20356 4284
rect 24494 13356 24814 14868
rect 24494 13300 24522 13356
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24786 13300 24814 13356
rect 24494 11788 24814 13300
rect 24494 11732 24522 11788
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24786 11732 24814 11788
rect 24494 10220 24814 11732
rect 24494 10164 24522 10220
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24786 10164 24814 10220
rect 24494 8652 24814 10164
rect 24494 8596 24522 8652
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24786 8596 24814 8652
rect 24494 7084 24814 8596
rect 24494 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24814 7084
rect 24494 5516 24814 7028
rect 24494 5460 24522 5516
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24786 5460 24814 5516
rect 19832 3108 19860 3164
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 20124 3108 20152 3164
rect 19832 3076 20152 3108
rect 24494 3948 24814 5460
rect 24494 3892 24522 3948
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24786 3892 24814 3948
rect 24494 3076 24814 3892
rect 29156 36092 29476 36908
rect 29156 36036 29184 36092
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29448 36036 29476 36092
rect 29156 34524 29476 36036
rect 29156 34468 29184 34524
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29448 34468 29476 34524
rect 29156 32956 29476 34468
rect 29156 32900 29184 32956
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29448 32900 29476 32956
rect 29156 31388 29476 32900
rect 29156 31332 29184 31388
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29448 31332 29476 31388
rect 29156 29820 29476 31332
rect 29156 29764 29184 29820
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29448 29764 29476 29820
rect 29156 28252 29476 29764
rect 29156 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29476 28252
rect 29156 26684 29476 28196
rect 29156 26628 29184 26684
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29448 26628 29476 26684
rect 29156 25116 29476 26628
rect 29156 25060 29184 25116
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29448 25060 29476 25116
rect 29156 23548 29476 25060
rect 29156 23492 29184 23548
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29448 23492 29476 23548
rect 29156 21980 29476 23492
rect 29156 21924 29184 21980
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29448 21924 29476 21980
rect 29156 20412 29476 21924
rect 29156 20356 29184 20412
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29448 20356 29476 20412
rect 29156 18844 29476 20356
rect 29156 18788 29184 18844
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29448 18788 29476 18844
rect 29156 17276 29476 18788
rect 29156 17220 29184 17276
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29448 17220 29476 17276
rect 29156 15708 29476 17220
rect 29156 15652 29184 15708
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29448 15652 29476 15708
rect 29156 14140 29476 15652
rect 29156 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29476 14140
rect 29156 12572 29476 14084
rect 29156 12516 29184 12572
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29448 12516 29476 12572
rect 29156 11004 29476 12516
rect 29156 10948 29184 11004
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29448 10948 29476 11004
rect 29156 9436 29476 10948
rect 29156 9380 29184 9436
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29448 9380 29476 9436
rect 29156 7868 29476 9380
rect 29156 7812 29184 7868
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29448 7812 29476 7868
rect 29156 6300 29476 7812
rect 29156 6244 29184 6300
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29448 6244 29476 6300
rect 29156 4732 29476 6244
rect 29156 4676 29184 4732
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29448 4676 29476 4732
rect 29156 3164 29476 4676
rect 29156 3108 29184 3164
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29448 3108 29476 3164
rect 29156 3076 29476 3108
rect 33818 36876 34138 36908
rect 33818 36820 33846 36876
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 34110 36820 34138 36876
rect 33818 35308 34138 36820
rect 33818 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34138 35308
rect 33818 33740 34138 35252
rect 33818 33684 33846 33740
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 34110 33684 34138 33740
rect 33818 32172 34138 33684
rect 33818 32116 33846 32172
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 34110 32116 34138 32172
rect 33818 30604 34138 32116
rect 33818 30548 33846 30604
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 34110 30548 34138 30604
rect 33818 29036 34138 30548
rect 33818 28980 33846 29036
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 34110 28980 34138 29036
rect 33818 27468 34138 28980
rect 33818 27412 33846 27468
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 34110 27412 34138 27468
rect 33818 25900 34138 27412
rect 33818 25844 33846 25900
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 34110 25844 34138 25900
rect 33818 24332 34138 25844
rect 33818 24276 33846 24332
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 34110 24276 34138 24332
rect 33818 22764 34138 24276
rect 33818 22708 33846 22764
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 34110 22708 34138 22764
rect 33818 21196 34138 22708
rect 33818 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34138 21196
rect 33818 19628 34138 21140
rect 33818 19572 33846 19628
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 34110 19572 34138 19628
rect 33818 18060 34138 19572
rect 33818 18004 33846 18060
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 34110 18004 34138 18060
rect 33818 16492 34138 18004
rect 33818 16436 33846 16492
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 34110 16436 34138 16492
rect 33818 14924 34138 16436
rect 33818 14868 33846 14924
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 34110 14868 34138 14924
rect 33818 13356 34138 14868
rect 33818 13300 33846 13356
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 34110 13300 34138 13356
rect 33818 11788 34138 13300
rect 33818 11732 33846 11788
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 34110 11732 34138 11788
rect 33818 10220 34138 11732
rect 33818 10164 33846 10220
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 34110 10164 34138 10220
rect 33818 8652 34138 10164
rect 33818 8596 33846 8652
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 34110 8596 34138 8652
rect 33818 7084 34138 8596
rect 33818 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34138 7084
rect 33818 5516 34138 7028
rect 33818 5460 33846 5516
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 34110 5460 34138 5516
rect 33818 3948 34138 5460
rect 33818 3892 33846 3948
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 34110 3892 34138 3948
rect 33818 3076 34138 3892
rect 38480 36092 38800 36908
rect 38480 36036 38508 36092
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38772 36036 38800 36092
rect 38480 34524 38800 36036
rect 38480 34468 38508 34524
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38772 34468 38800 34524
rect 38480 32956 38800 34468
rect 38480 32900 38508 32956
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38772 32900 38800 32956
rect 38480 31388 38800 32900
rect 38480 31332 38508 31388
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38772 31332 38800 31388
rect 38480 29820 38800 31332
rect 38480 29764 38508 29820
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38772 29764 38800 29820
rect 38480 28252 38800 29764
rect 38480 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38800 28252
rect 38480 26684 38800 28196
rect 38480 26628 38508 26684
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38772 26628 38800 26684
rect 38480 25116 38800 26628
rect 38480 25060 38508 25116
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38772 25060 38800 25116
rect 38480 23548 38800 25060
rect 38480 23492 38508 23548
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38772 23492 38800 23548
rect 38480 21980 38800 23492
rect 38480 21924 38508 21980
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38772 21924 38800 21980
rect 38480 20412 38800 21924
rect 38480 20356 38508 20412
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38772 20356 38800 20412
rect 38480 18844 38800 20356
rect 38480 18788 38508 18844
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38772 18788 38800 18844
rect 38480 17276 38800 18788
rect 38480 17220 38508 17276
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38772 17220 38800 17276
rect 38480 15708 38800 17220
rect 38480 15652 38508 15708
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38772 15652 38800 15708
rect 38480 14140 38800 15652
rect 38480 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38800 14140
rect 38480 12572 38800 14084
rect 38480 12516 38508 12572
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38772 12516 38800 12572
rect 38480 11004 38800 12516
rect 38480 10948 38508 11004
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38772 10948 38800 11004
rect 38480 9436 38800 10948
rect 38480 9380 38508 9436
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38772 9380 38800 9436
rect 38480 7868 38800 9380
rect 38480 7812 38508 7868
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38772 7812 38800 7868
rect 38480 6300 38800 7812
rect 38480 6244 38508 6300
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38772 6244 38800 6300
rect 38480 4732 38800 6244
rect 38480 4676 38508 4732
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38772 4676 38800 4732
rect 38480 3164 38800 4676
rect 38480 3108 38508 3164
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38772 3108 38800 3164
rect 38480 3076 38800 3108
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _102_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23408 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _103_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20496 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20944 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698431365
transform 1 0 24192 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _106_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _107_
timestamp 1698431365
transform -1 0 22736 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698431365
transform 1 0 23072 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _109_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25312 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _110_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21728 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _111_
timestamp 1698431365
transform -1 0 25984 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _112_
timestamp 1698431365
transform -1 0 13776 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _113_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15456 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _114_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _115_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _116_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23184 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _117_
timestamp 1698431365
transform -1 0 21840 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _118_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19824 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _119_
timestamp 1698431365
transform 1 0 19488 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _120_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18368 0 1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698431365
transform -1 0 22848 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _122_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19488 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _123_
timestamp 1698431365
transform -1 0 18144 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _124_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15008 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _125_
timestamp 1698431365
transform 1 0 14560 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _126_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20832 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _127_
timestamp 1698431365
transform -1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _128_
timestamp 1698431365
transform -1 0 20048 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _129_
timestamp 1698431365
transform 1 0 16128 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _130_
timestamp 1698431365
transform -1 0 13104 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _131_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16800 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _132_
timestamp 1698431365
transform 1 0 21728 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_
timestamp 1698431365
transform -1 0 21728 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _134_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17808 0 -1 25088
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _135_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 1 23520
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _136_
timestamp 1698431365
transform 1 0 17248 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _137_
timestamp 1698431365
transform -1 0 16800 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _138_
timestamp 1698431365
transform 1 0 21728 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _139_
timestamp 1698431365
transform -1 0 21840 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _140_
timestamp 1698431365
transform 1 0 17808 0 -1 26656
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _141_
timestamp 1698431365
transform 1 0 17248 0 1 25088
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _142_
timestamp 1698431365
transform 1 0 12208 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _143_
timestamp 1698431365
transform -1 0 15792 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _144_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _145_
timestamp 1698431365
transform 1 0 25424 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698431365
transform -1 0 23184 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _147_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13552 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _148_
timestamp 1698431365
transform -1 0 13104 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _149_
timestamp 1698431365
transform -1 0 15344 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _150_
timestamp 1698431365
transform 1 0 12208 0 -1 21952
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _151_
timestamp 1698431365
transform 1 0 13328 0 -1 25088
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _152_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _153_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21952 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _154_
timestamp 1698431365
transform 1 0 23520 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _155_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23856 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698431365
transform -1 0 22176 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_2  _157_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26432 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698431365
transform 1 0 21728 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698431365
transform -1 0 21728 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _160_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22736 0 -1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _161_
timestamp 1698431365
transform 1 0 18144 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _162_
timestamp 1698431365
transform 1 0 23856 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _163_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23072 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _164_
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _165_
timestamp 1698431365
transform 1 0 18368 0 -1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _166_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _167_
timestamp 1698431365
transform -1 0 18816 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _168_
timestamp 1698431365
transform -1 0 20160 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _169_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _170_
timestamp 1698431365
transform -1 0 21840 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _171_
timestamp 1698431365
transform -1 0 23744 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _172_
timestamp 1698431365
transform 1 0 22624 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _173_
timestamp 1698431365
transform -1 0 19152 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _174_
timestamp 1698431365
transform 1 0 18704 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _175_
timestamp 1698431365
transform -1 0 20720 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _176_
timestamp 1698431365
transform 1 0 20384 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _177_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20832 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _178_
timestamp 1698431365
transform 1 0 18256 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _179_
timestamp 1698431365
transform 1 0 21280 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _180_
timestamp 1698431365
transform 1 0 18704 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _181_
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _182_
timestamp 1698431365
transform -1 0 20832 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _183_
timestamp 1698431365
transform 1 0 18704 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _184_
timestamp 1698431365
transform 1 0 22624 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _185_
timestamp 1698431365
transform 1 0 18704 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _186_
timestamp 1698431365
transform -1 0 18704 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _187_
timestamp 1698431365
transform -1 0 22624 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _188_
timestamp 1698431365
transform 1 0 11984 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _189_
timestamp 1698431365
transform -1 0 18144 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _190_
timestamp 1698431365
transform -1 0 18144 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _191_
timestamp 1698431365
transform -1 0 15232 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _192_
timestamp 1698431365
transform -1 0 19600 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _193_
timestamp 1698431365
transform 1 0 23744 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _194_
timestamp 1698431365
transform 1 0 25200 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _195_
timestamp 1698431365
transform -1 0 18704 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _196_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _197_
timestamp 1698431365
transform -1 0 20944 0 -1 20384
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _198_
timestamp 1698431365
transform 1 0 12208 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _199_
timestamp 1698431365
transform -1 0 15456 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _200_
timestamp 1698431365
transform 1 0 25760 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _201_
timestamp 1698431365
transform -1 0 20720 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _202_
timestamp 1698431365
transform 1 0 12208 0 -1 20384
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _203_
timestamp 1698431365
transform 1 0 13328 0 -1 17248
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _204_
timestamp 1698431365
transform 1 0 13552 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _205_
timestamp 1698431365
transform -1 0 13104 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _206_
timestamp 1698431365
transform 1 0 25200 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _207_
timestamp 1698431365
transform -1 0 20160 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _208_
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _209_
timestamp 1698431365
transform 1 0 13328 0 -1 18816
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _210_
timestamp 1698431365
transform 1 0 15456 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _211_
timestamp 1698431365
transform -1 0 16352 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _212_
timestamp 1698431365
transform 1 0 21280 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _213_
timestamp 1698431365
transform -1 0 18704 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _214_
timestamp 1698431365
transform -1 0 19488 0 1 21952
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _215_
timestamp 1698431365
transform 1 0 15232 0 1 17248
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__I test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23408 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__I
timestamp 1698431365
transform -1 0 14000 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__114__A1
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__A2
timestamp 1698431365
transform -1 0 17808 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__A2
timestamp 1698431365
transform -1 0 12208 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__I
timestamp 1698431365
transform 1 0 24192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__S1
timestamp 1698431365
transform 1 0 26208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__I2
timestamp 1698431365
transform -1 0 27888 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__S0
timestamp 1698431365
transform -1 0 28336 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__I
timestamp 1698431365
transform -1 0 20496 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__I3
timestamp 1698431365
transform -1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__A2
timestamp 1698431365
transform 1 0 11760 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__B1
timestamp 1698431365
transform 1 0 11312 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I2
timestamp 1698431365
transform 1 0 29232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 37744 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 37744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 37744 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 37744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 26992 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 25536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 37744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 30912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 27888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 29568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 28448 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 37744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 37520 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 37520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 2464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 14560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 15232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 3136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 21616 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 20496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform -1 0 26432 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform -1 0 20048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 20944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 2464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform 1 0 3136 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 2912 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform 1 0 2464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 15904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 12768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 2464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 37744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 37296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 12096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform -1 0 14224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform 1 0 2464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform 1 0 3584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform 1 0 3136 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform -1 0 37296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform -1 0 25984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform 1 0 37520 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform -1 0 23184 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform -1 0 37744 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform -1 0 37744 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698431365
transform -1 0 24416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698431365
transform -1 0 23520 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698431365
transform -1 0 25536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1698431365
transform -1 0 37744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1698431365
transform -1 0 37296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1698431365
transform -1 0 37744 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1698431365
transform -1 0 22288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1698431365
transform -1 0 28560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1698431365
transform -1 0 37296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1698431365
transform -1 0 24416 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1698431365
transform -1 0 23856 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1698431365
transform -1 0 37744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1698431365
transform -1 0 37744 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1698431365
transform -1 0 26432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1698431365
transform -1 0 30240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1698431365
transform -1 0 25984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1698431365
transform -1 0 37744 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1698431365
transform -1 0 37744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1698431365
transform -1 0 26992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1698431365
transform -1 0 37744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1698431365
transform -1 0 37296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1698431365
transform 1 0 19824 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1698431365
transform -1 0 16576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1698431365
transform -1 0 10304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1698431365
transform 1 0 2912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1698431365
transform -1 0 18928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1698431365
transform -1 0 15568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1698431365
transform -1 0 18256 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1698431365
transform -1 0 17696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1698431365
transform -1 0 29008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1698431365
transform 1 0 2464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input83_I
timestamp 1698431365
transform -1 0 18256 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input84_I
timestamp 1698431365
transform 1 0 14000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input85_I
timestamp 1698431365
transform -1 0 10752 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input86_I
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input87_I
timestamp 1698431365
transform -1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input88_I
timestamp 1698431365
transform -1 0 16912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input89_I
timestamp 1698431365
transform -1 0 37744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input90_I
timestamp 1698431365
transform -1 0 18928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input91_I
timestamp 1698431365
transform 1 0 16576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input92_I
timestamp 1698431365
transform 1 0 2464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input93_I
timestamp 1698431365
transform 1 0 2912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input94_I
timestamp 1698431365
transform 1 0 3136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input95_I
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input96_I
timestamp 1698431365
transform -1 0 37744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input97_I
timestamp 1698431365
transform -1 0 37744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input98_I
timestamp 1698431365
transform -1 0 37744 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input99_I
timestamp 1698431365
transform -1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_70 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_86 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10976 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_163
timestamp 1698431365
transform 1 0 19600 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_270
timestamp 1698431365
transform 1 0 31584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_324 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_328
timestamp 1698431365
transform 1 0 38080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_330
timestamp 1698431365
transform 1 0 38304 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_88
timestamp 1698431365
transform 1 0 11200 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_96
timestamp 1698431365
transform 1 0 12096 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_123
timestamp 1698431365
transform 1 0 15120 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_133
timestamp 1698431365
transform 1 0 16240 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_146
timestamp 1698431365
transform 1 0 17696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_148
timestamp 1698431365
transform 1 0 17920 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_151
timestamp 1698431365
transform 1 0 18256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_157
timestamp 1698431365
transform 1 0 18928 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_167
timestamp 1698431365
transform 1 0 20048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_171
timestamp 1698431365
transform 1 0 20496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_193
timestamp 1698431365
transform 1 0 22960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_195
timestamp 1698431365
transform 1 0 23184 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_198
timestamp 1698431365
transform 1 0 23520 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_202
timestamp 1698431365
transform 1 0 23968 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_216
timestamp 1698431365
transform 1 0 25536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_224
timestamp 1698431365
transform 1 0 26432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_226
timestamp 1698431365
transform 1 0 26656 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_235
timestamp 1698431365
transform 1 0 27664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_239
timestamp 1698431365
transform 1 0 28112 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_243
timestamp 1698431365
transform 1 0 28560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_247
timestamp 1698431365
transform 1 0 29008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_249
timestamp 1698431365
transform 1 0 29232 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_252
timestamp 1698431365
transform 1 0 29568 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_258
timestamp 1698431365
transform 1 0 30240 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_264
timestamp 1698431365
transform 1 0 30912 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_314
timestamp 1698431365
transform 1 0 36512 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_330
timestamp 1698431365
transform 1 0 38304 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_111
timestamp 1698431365
transform 1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_127
timestamp 1698431365
transform 1 0 15568 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_135
timestamp 1698431365
transform 1 0 16464 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_138
timestamp 1698431365
transform 1 0 16800 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_170
timestamp 1698431365
transform 1 0 20384 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_187
timestamp 1698431365
transform 1 0 22288 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_219
timestamp 1698431365
transform 1 0 25872 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_235
timestamp 1698431365
transform 1 0 27664 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698431365
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_325
timestamp 1698431365
transform 1 0 37744 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_329
timestamp 1698431365
transform 1 0 38192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_314
timestamp 1698431365
transform 1 0 36512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_330
timestamp 1698431365
transform 1 0 38304 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_325
timestamp 1698431365
transform 1 0 37744 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_329
timestamp 1698431365
transform 1 0 38192 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_314
timestamp 1698431365
transform 1 0 36512 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_330
timestamp 1698431365
transform 1 0 38304 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_325
timestamp 1698431365
transform 1 0 37744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_329
timestamp 1698431365
transform 1 0 38192 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_314
timestamp 1698431365
transform 1 0 36512 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_330
timestamp 1698431365
transform 1 0 38304 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_329
timestamp 1698431365
transform 1 0 38192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_314
timestamp 1698431365
transform 1 0 36512 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_322
timestamp 1698431365
transform 1 0 37408 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_321
timestamp 1698431365
transform 1 0 37296 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_28
timestamp 1698431365
transform 1 0 4480 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_60
timestamp 1698431365
transform 1 0 8064 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_68
timestamp 1698431365
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_150
timestamp 1698431365
transform 1 0 18144 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_154
timestamp 1698431365
transform 1 0 18592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_180
timestamp 1698431365
transform 1 0 21504 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_196
timestamp 1698431365
transform 1 0 23296 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_204
timestamp 1698431365
transform 1 0 24192 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_314
timestamp 1698431365
transform 1 0 36512 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_318
timestamp 1698431365
transform 1 0 36960 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_321
timestamp 1698431365
transform 1 0 37296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_28
timestamp 1698431365
transform 1 0 4480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698431365
transform 1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_139
timestamp 1698431365
transform 1 0 16912 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_170
timestamp 1698431365
transform 1 0 20384 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_187
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_189
timestamp 1698431365
transform 1 0 22512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_222
timestamp 1698431365
transform 1 0 26208 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_238
timestamp 1698431365
transform 1 0 28000 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698431365
transform 1 0 28448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_14
timestamp 1698431365
transform 1 0 2912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_18
timestamp 1698431365
transform 1 0 3360 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_22
timestamp 1698431365
transform 1 0 3808 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_54
timestamp 1698431365
transform 1 0 7392 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_144
timestamp 1698431365
transform 1 0 17472 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_170
timestamp 1698431365
transform 1 0 20384 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_314
timestamp 1698431365
transform 1 0 36512 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_322
timestamp 1698431365
transform 1 0 37408 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_8
timestamp 1698431365
transform 1 0 2240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_12
timestamp 1698431365
transform 1 0 2688 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_28
timestamp 1698431365
transform 1 0 4480 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_32
timestamp 1698431365
transform 1 0 4928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_139
timestamp 1698431365
transform 1 0 16912 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_155
timestamp 1698431365
transform 1 0 18704 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_159
timestamp 1698431365
transform 1 0 19152 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_222
timestamp 1698431365
transform 1 0 26208 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_238
timestamp 1698431365
transform 1 0 28000 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698431365
transform 1 0 28448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_321
timestamp 1698431365
transform 1 0 37296 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_8
timestamp 1698431365
transform 1 0 2240 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_12
timestamp 1698431365
transform 1 0 2688 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_44
timestamp 1698431365
transform 1 0 6272 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_60
timestamp 1698431365
transform 1 0 8064 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1698431365
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_104
timestamp 1698431365
transform 1 0 12992 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_108
timestamp 1698431365
transform 1 0 13440 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_110
timestamp 1698431365
transform 1 0 13664 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_150
timestamp 1698431365
transform 1 0 18144 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_184
timestamp 1698431365
transform 1 0 21952 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_200
timestamp 1698431365
transform 1 0 23744 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698431365
transform 1 0 36512 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_322
timestamp 1698431365
transform 1 0 37408 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_8
timestamp 1698431365
transform 1 0 2240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_12
timestamp 1698431365
transform 1 0 2688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_16
timestamp 1698431365
transform 1 0 3136 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698431365
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_134
timestamp 1698431365
transform 1 0 16352 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_165
timestamp 1698431365
transform 1 0 19824 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698431365
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698431365
transform 1 0 37296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_14
timestamp 1698431365
transform 1 0 2912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_18
timestamp 1698431365
transform 1 0 3360 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_50
timestamp 1698431365
transform 1 0 6944 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_88
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_96
timestamp 1698431365
transform 1 0 12096 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_146
timestamp 1698431365
transform 1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_173
timestamp 1698431365
transform 1 0 20720 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_177
timestamp 1698431365
transform 1 0 21168 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_216
timestamp 1698431365
transform 1 0 25536 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_250
timestamp 1698431365
transform 1 0 29344 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_266
timestamp 1698431365
transform 1 0 31136 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_274
timestamp 1698431365
transform 1 0 32032 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698431365
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_314
timestamp 1698431365
transform 1 0 36512 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_318
timestamp 1698431365
transform 1 0 36960 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_321
timestamp 1698431365
transform 1 0 37296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698431365
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698431365
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_69
timestamp 1698431365
transform 1 0 9072 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_85
timestamp 1698431365
transform 1 0 10864 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_89
timestamp 1698431365
transform 1 0 11312 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698431365
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_183
timestamp 1698431365
transform 1 0 21840 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_185
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_206
timestamp 1698431365
transform 1 0 24416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_210
timestamp 1698431365
transform 1 0 24864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_212
timestamp 1698431365
transform 1 0 25088 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_251
timestamp 1698431365
transform 1 0 29456 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_283
timestamp 1698431365
transform 1 0 33040 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_299
timestamp 1698431365
transform 1 0 34832 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_307
timestamp 1698431365
transform 1 0 35728 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_8
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_12
timestamp 1698431365
transform 1 0 2688 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_44
timestamp 1698431365
transform 1 0 6272 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698431365
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_104
timestamp 1698431365
transform 1 0 12992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_106
timestamp 1698431365
transform 1 0 13216 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_150
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_167
timestamp 1698431365
transform 1 0 20048 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_171
timestamp 1698431365
transform 1 0 20496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_183
timestamp 1698431365
transform 1 0 21840 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_195
timestamp 1698431365
transform 1 0 23184 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_203
timestamp 1698431365
transform 1 0 24080 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_220
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_252
timestamp 1698431365
transform 1 0 29568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_268
timestamp 1698431365
transform 1 0 31360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698431365
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698431365
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698431365
transform 1 0 4480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698431365
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_69
timestamp 1698431365
transform 1 0 9072 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_85
timestamp 1698431365
transform 1 0 10864 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_93
timestamp 1698431365
transform 1 0 11760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_186
timestamp 1698431365
transform 1 0 22176 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_202
timestamp 1698431365
transform 1 0 23968 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_210
timestamp 1698431365
transform 1 0 24864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_212
timestamp 1698431365
transform 1 0 25088 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698431365
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698431365
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_8
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_12
timestamp 1698431365
transform 1 0 2688 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_44
timestamp 1698431365
transform 1 0 6272 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698431365
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698431365
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_88
timestamp 1698431365
transform 1 0 11200 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_96
timestamp 1698431365
transform 1 0 12096 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_175
timestamp 1698431365
transform 1 0 20944 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_201
timestamp 1698431365
transform 1 0 23856 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_203
timestamp 1698431365
transform 1 0 24080 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_220
timestamp 1698431365
transform 1 0 25984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_258
timestamp 1698431365
transform 1 0 30240 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_274
timestamp 1698431365
transform 1 0 32032 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698431365
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698431365
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698431365
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_8
timestamp 1698431365
transform 1 0 2240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_12
timestamp 1698431365
transform 1 0 2688 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698431365
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698431365
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_69
timestamp 1698431365
transform 1 0 9072 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_85
timestamp 1698431365
transform 1 0 10864 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_91
timestamp 1698431365
transform 1 0 11536 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_200
timestamp 1698431365
transform 1 0 23744 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_233
timestamp 1698431365
transform 1 0 27440 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_237
timestamp 1698431365
transform 1 0 27888 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698431365
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_8
timestamp 1698431365
transform 1 0 2240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_12
timestamp 1698431365
transform 1 0 2688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_16
timestamp 1698431365
transform 1 0 3136 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_48
timestamp 1698431365
transform 1 0 6720 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_64
timestamp 1698431365
transform 1 0 8512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_88
timestamp 1698431365
transform 1 0 11200 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_92
timestamp 1698431365
transform 1 0 11648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_94
timestamp 1698431365
transform 1 0 11872 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_197
timestamp 1698431365
transform 1 0 23408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698431365
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_220
timestamp 1698431365
transform 1 0 25984 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_252
timestamp 1698431365
transform 1 0 29568 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_268
timestamp 1698431365
transform 1 0 31360 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_314
timestamp 1698431365
transform 1 0 36512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_318
timestamp 1698431365
transform 1 0 36960 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_321
timestamp 1698431365
transform 1 0 37296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_14
timestamp 1698431365
transform 1 0 2912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_18
timestamp 1698431365
transform 1 0 3360 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_170
timestamp 1698431365
transform 1 0 20384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698431365
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_187
timestamp 1698431365
transform 1 0 22288 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_195
timestamp 1698431365
transform 1 0 23184 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_199
timestamp 1698431365
transform 1 0 23632 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_203
timestamp 1698431365
transform 1 0 24080 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_206
timestamp 1698431365
transform 1 0 24416 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_238
timestamp 1698431365
transform 1 0 28000 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698431365
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_311
timestamp 1698431365
transform 1 0 36176 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_8
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_12
timestamp 1698431365
transform 1 0 2688 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_44
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698431365
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698431365
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_88
timestamp 1698431365
transform 1 0 11200 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_96
timestamp 1698431365
transform 1 0 12096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_100
timestamp 1698431365
transform 1 0 12544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_102
timestamp 1698431365
transform 1 0 12768 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_125
timestamp 1698431365
transform 1 0 15344 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_150
timestamp 1698431365
transform 1 0 18144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_181
timestamp 1698431365
transform 1 0 21616 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_189
timestamp 1698431365
transform 1 0 22512 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_193
timestamp 1698431365
transform 1 0 22960 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_200
timestamp 1698431365
transform 1 0 23744 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_208
timestamp 1698431365
transform 1 0 24640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_246
timestamp 1698431365
transform 1 0 28896 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698431365
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698431365
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_8
timestamp 1698431365
transform 1 0 2240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_12
timestamp 1698431365
transform 1 0 2688 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_69
timestamp 1698431365
transform 1 0 9072 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_85
timestamp 1698431365
transform 1 0 10864 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_93
timestamp 1698431365
transform 1 0 11760 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_113
timestamp 1698431365
transform 1 0 14000 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_129
timestamp 1698431365
transform 1 0 15792 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_131
timestamp 1698431365
transform 1 0 16016 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_140
timestamp 1698431365
transform 1 0 17024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_214
timestamp 1698431365
transform 1 0 25312 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_230
timestamp 1698431365
transform 1 0 27104 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_238
timestamp 1698431365
transform 1 0 28000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698431365
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698431365
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_8
timestamp 1698431365
transform 1 0 2240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_12
timestamp 1698431365
transform 1 0 2688 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_44
timestamp 1698431365
transform 1 0 6272 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698431365
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698431365
transform 1 0 11200 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_96
timestamp 1698431365
transform 1 0 12096 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_146
timestamp 1698431365
transform 1 0 17696 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_195
timestamp 1698431365
transform 1 0 23184 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_203
timestamp 1698431365
transform 1 0 24080 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698431365
transform 1 0 24528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_214
timestamp 1698431365
transform 1 0 25312 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_247
timestamp 1698431365
transform 1 0 29008 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698431365
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698431365
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_8
timestamp 1698431365
transform 1 0 2240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_12
timestamp 1698431365
transform 1 0 2688 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_122
timestamp 1698431365
transform 1 0 15008 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_138
timestamp 1698431365
transform 1 0 16800 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_214
timestamp 1698431365
transform 1 0 25312 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_230
timestamp 1698431365
transform 1 0 27104 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698431365
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698431365
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698431365
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698431365
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_8
timestamp 1698431365
transform 1 0 2240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_12
timestamp 1698431365
transform 1 0 2688 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_44
timestamp 1698431365
transform 1 0 6272 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698431365
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_104
timestamp 1698431365
transform 1 0 12992 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_112
timestamp 1698431365
transform 1 0 13888 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_116
timestamp 1698431365
transform 1 0 14336 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_144
timestamp 1698431365
transform 1 0 17472 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_190
timestamp 1698431365
transform 1 0 22624 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_314
timestamp 1698431365
transform 1 0 36512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_318
timestamp 1698431365
transform 1 0 36960 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_321
timestamp 1698431365
transform 1 0 37296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_14
timestamp 1698431365
transform 1 0 2912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_18
timestamp 1698431365
transform 1 0 3360 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_123
timestamp 1698431365
transform 1 0 15120 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_131
timestamp 1698431365
transform 1 0 16016 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_183
timestamp 1698431365
transform 1 0 21840 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_215
timestamp 1698431365
transform 1 0 25424 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_231
timestamp 1698431365
transform 1 0 27216 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_239
timestamp 1698431365
transform 1 0 28112 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698431365
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_8
timestamp 1698431365
transform 1 0 2240 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_12
timestamp 1698431365
transform 1 0 2688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_16
timestamp 1698431365
transform 1 0 3136 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_48
timestamp 1698431365
transform 1 0 6720 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_64
timestamp 1698431365
transform 1 0 8512 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698431365
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_158
timestamp 1698431365
transform 1 0 19040 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_160
timestamp 1698431365
transform 1 0 19264 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_174
timestamp 1698431365
transform 1 0 20832 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_314
timestamp 1698431365
transform 1 0 36512 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_318
timestamp 1698431365
transform 1 0 36960 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_321
timestamp 1698431365
transform 1 0 37296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_8
timestamp 1698431365
transform 1 0 2240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_12
timestamp 1698431365
transform 1 0 2688 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_28
timestamp 1698431365
transform 1 0 4480 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_32
timestamp 1698431365
transform 1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_321
timestamp 1698431365
transform 1 0 37296 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_28
timestamp 1698431365
transform 1 0 4480 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_60
timestamp 1698431365
transform 1 0 8064 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698431365
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_314
timestamp 1698431365
transform 1 0 36512 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_322
timestamp 1698431365
transform 1 0 37408 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_321
timestamp 1698431365
transform 1 0 37296 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_314
timestamp 1698431365
transform 1 0 36512 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_322
timestamp 1698431365
transform 1 0 37408 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_325
timestamp 1698431365
transform 1 0 37744 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_329
timestamp 1698431365
transform 1 0 38192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_314
timestamp 1698431365
transform 1 0 36512 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_330
timestamp 1698431365
transform 1 0 38304 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_325
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_329
timestamp 1698431365
transform 1 0 38192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_314
timestamp 1698431365
transform 1 0 36512 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_330
timestamp 1698431365
transform 1 0 38304 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698431365
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_139
timestamp 1698431365
transform 1 0 16912 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_147
timestamp 1698431365
transform 1 0 17808 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_151
timestamp 1698431365
transform 1 0 18256 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_157
timestamp 1698431365
transform 1 0 18928 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_187
timestamp 1698431365
transform 1 0 22288 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_191
timestamp 1698431365
transform 1 0 22736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_195
timestamp 1698431365
transform 1 0 23184 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_201
timestamp 1698431365
transform 1 0 23856 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_203
timestamp 1698431365
transform 1 0 24080 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_206
timestamp 1698431365
transform 1 0 24416 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_238
timestamp 1698431365
transform 1 0 28000 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_242
timestamp 1698431365
transform 1 0 28448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698431365
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_325
timestamp 1698431365
transform 1 0 37744 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_329
timestamp 1698431365
transform 1 0 38192 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_80
timestamp 1698431365
transform 1 0 10304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_84
timestamp 1698431365
transform 1 0 10752 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_111
timestamp 1698431365
transform 1 0 13776 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_115
timestamp 1698431365
transform 1 0 14224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_117
timestamp 1698431365
transform 1 0 14448 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_120
timestamp 1698431365
transform 1 0 14784 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_126
timestamp 1698431365
transform 1 0 15456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_132
timestamp 1698431365
transform 1 0 16128 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_144
timestamp 1698431365
transform 1 0 17472 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_163
timestamp 1698431365
transform 1 0 19600 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_167
timestamp 1698431365
transform 1 0 20048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_207
timestamp 1698431365
transform 1 0 24528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_209
timestamp 1698431365
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_216
timestamp 1698431365
transform 1 0 25536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_220
timestamp 1698431365
transform 1 0 25984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_224
timestamp 1698431365
transform 1 0 26432 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_226
timestamp 1698431365
transform 1 0 26656 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_235
timestamp 1698431365
transform 1 0 27664 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_267
timestamp 1698431365
transform 1 0 31248 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_275
timestamp 1698431365
transform 1 0 32144 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_314
timestamp 1698431365
transform 1 0 36512 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_330
timestamp 1698431365
transform 1 0 38304 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_36
timestamp 1698431365
transform 1 0 5376 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_70
timestamp 1698431365
transform 1 0 9184 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_80
timestamp 1698431365
transform 1 0 10304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_172
timestamp 1698431365
transform 1 0 20608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_201
timestamp 1698431365
transform 1 0 23856 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_203
timestamp 1698431365
transform 1 0 24080 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_236
timestamp 1698431365
transform 1 0 27776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_240
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_244
timestamp 1698431365
transform 1 0 28672 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_260
timestamp 1698431365
transform 1 0 30464 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_268
timestamp 1698431365
transform 1 0 31360 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_274
timestamp 1698431365
transform 1 0 32032 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_308
timestamp 1698431365
transform 1 0 35840 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_324
timestamp 1698431365
transform 1 0 37632 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_328
timestamp 1698431365
transform 1 0 38080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_330
timestamp 1698431365
transform 1 0 38304 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 38416 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 38416 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 38416 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 38416 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 27664 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 25760 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 37520 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform -1 0 38416 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 31584 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 27776 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform -1 0 30240 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 27776 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform -1 0 38416 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 38416 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform -1 0 37744 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 37744 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 13888 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 14560 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 2240 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform 1 0 21616 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 21616 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform -1 0 27104 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 22288 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 2240 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 15232 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 12096 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform -1 0 38416 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform -1 0 38416 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 12096 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 14896 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform 1 0 14224 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform 1 0 2240 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698431365
transform -1 0 38416 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698431365
transform -1 0 26432 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1698431365
transform -1 0 37744 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698431365
transform -1 0 23856 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698431365
transform -1 0 38416 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698431365
transform -1 0 38416 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1698431365
transform -1 0 25088 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1698431365
transform -1 0 24192 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1698431365
transform -1 0 25760 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1698431365
transform -1 0 38416 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input53
timestamp 1698431365
transform -1 0 38416 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1698431365
transform -1 0 38416 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1698431365
transform -1 0 22960 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input56
timestamp 1698431365
transform -1 0 28896 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input57
timestamp 1698431365
transform -1 0 38416 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input58
timestamp 1698431365
transform -1 0 25088 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input59
timestamp 1698431365
transform -1 0 24528 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1698431365
transform -1 0 38416 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1698431365
transform -1 0 38416 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input62
timestamp 1698431365
transform -1 0 27104 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input63
timestamp 1698431365
transform -1 0 30912 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input64
timestamp 1698431365
transform -1 0 26432 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input65
timestamp 1698431365
transform -1 0 38416 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input66
timestamp 1698431365
transform -1 0 38416 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input67
timestamp 1698431365
transform -1 0 27664 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input68
timestamp 1698431365
transform -1 0 38416 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input69
timestamp 1698431365
transform -1 0 38416 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input70
timestamp 1698431365
transform 1 0 19712 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input71
timestamp 1698431365
transform 1 0 15904 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input72
timestamp 1698431365
transform 1 0 10752 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input73
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input74
timestamp 1698431365
transform 1 0 18928 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input75
timestamp 1698431365
transform 1 0 15568 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input76
timestamp 1698431365
transform -1 0 18928 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input77
timestamp 1698431365
transform 1 0 17584 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input78
timestamp 1698431365
transform -1 0 29568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input79
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input80
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input81
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input82
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input83
timestamp 1698431365
transform 1 0 18256 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input84
timestamp 1698431365
transform 1 0 13216 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input85
timestamp 1698431365
transform 1 0 11424 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input86
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input87
timestamp 1698431365
transform 1 0 17584 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input88
timestamp 1698431365
transform 1 0 16912 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input89
timestamp 1698431365
transform -1 0 38416 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input90
timestamp 1698431365
transform -1 0 19600 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input91
timestamp 1698431365
transform 1 0 15904 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input92
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input93
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input94
timestamp 1698431365
transform 1 0 2240 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input95
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input96
timestamp 1698431365
transform -1 0 38416 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input97
timestamp 1698431365
transform -1 0 38416 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input98
timestamp 1698431365
transform -1 0 38416 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input99
timestamp 1698431365
transform -1 0 38416 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output100 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20272 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output101
timestamp 1698431365
transform -1 0 4480 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output102
timestamp 1698431365
transform -1 0 4480 0 1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output103
timestamp 1698431365
transform -1 0 13776 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output104
timestamp 1698431365
transform -1 0 19712 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output105
timestamp 1698431365
transform -1 0 4480 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output106
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output107
timestamp 1698431365
transform -1 0 15120 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output108
timestamp 1698431365
transform -1 0 15904 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output109
timestamp 1698431365
transform -1 0 23520 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output110
timestamp 1698431365
transform -1 0 4480 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output111
timestamp 1698431365
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_43 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_44
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 38640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_45
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 38640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_46
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_47
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_48
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 38640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_49
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 38640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_50
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 38640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_51
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_52
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 38640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_53
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 38640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 38640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 38640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 38640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 38640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 38640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 38640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 38640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 38640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 38640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 38640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 38640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 38640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 38640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 38640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 38640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 38640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 38640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 38640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 38640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_86 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_87
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_88
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_89
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_95
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_96
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_97
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_98
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_99
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_100
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_101
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_102
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_103
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_104
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_105
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_106
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_107
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_108
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_109
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_110
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_111
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_112
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_113
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_114
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_115
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_116
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_117
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_118
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_119
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_120
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_121
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_122
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_123
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_124
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_125
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_126
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_127
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_128
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_129
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_130
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_131
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_132
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_133
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_134
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_135
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_136
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_137
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_138
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_139
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_140
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_141
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_142
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_143
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_144
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_145
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_146
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_147
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_148
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_149
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_150
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_151
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_152
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_153
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_154
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_155
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_156
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_157
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_158
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_159
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_160
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_161
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_162
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_163
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_164
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_165
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_166
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_167
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_168
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_169
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_170
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_171
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_172
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_173
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_174
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_175
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_176
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_177
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_178
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_179
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_180
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_181
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_182
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_183
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_184
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_185
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_186
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_187
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_188
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_189
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_190
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_191
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_192
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_193
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_194
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_195
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_196
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_197
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_198
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_199
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_200
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_201
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_202
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_203
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_204
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_205
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_206
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_207
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_208
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_209
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_210
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_211
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_212
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_213
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_214
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_215
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_216
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_217
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_218
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_219
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_220
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_221
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_222
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_223
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_224
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_225
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_226
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_227
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_228
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_229
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_230
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_231
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_232
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_233
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_234
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_235
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_236
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_237
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_238
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_239
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_240
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_241
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_242
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_243
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_244
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_245
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_246
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_247
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_248
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_249
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_250
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_251
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_252
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_253
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_254
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_255
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_256
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_257
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_258
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_259
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_260
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_261
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_262
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_263
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_264
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_265
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_266
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_267
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_268
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_269
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_270
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_271
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_272
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_273
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_274
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_275
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_276
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_277
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_278
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_279
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_280
timestamp 1698431365
transform 1 0 8960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_281
timestamp 1698431365
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_282
timestamp 1698431365
transform 1 0 16576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_283
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698431365
transform 1 0 24192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698431365
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698431365
transform 1 0 31808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 310 870
<< labels >>
flabel metal2 s 20160 39200 20272 40000 0 FreeSans 448 90 0 0 out[0]
port 0 nsew signal tristate
flabel metal3 s 0 11424 800 11536 0 FreeSans 448 0 0 0 out[10]
port 1 nsew signal tristate
flabel metal3 s 0 12096 800 12208 0 FreeSans 448 0 0 0 out[11]
port 2 nsew signal tristate
flabel metal2 s 10752 39200 10864 40000 0 FreeSans 448 90 0 0 out[1]
port 3 nsew signal tristate
flabel metal2 s 16128 39200 16240 40000 0 FreeSans 448 90 0 0 out[2]
port 4 nsew signal tristate
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 out[3]
port 5 nsew signal tristate
flabel metal2 s 20832 39200 20944 40000 0 FreeSans 448 90 0 0 out[4]
port 6 nsew signal tristate
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 out[5]
port 7 nsew signal tristate
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 out[6]
port 8 nsew signal tristate
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 out[7]
port 9 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 out[8]
port 10 nsew signal tristate
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 out[9]
port 11 nsew signal tristate
flabel metal3 s 39200 30240 40000 30352 0 FreeSans 448 0 0 0 proj_out[0]
port 12 nsew signal input
flabel metal3 s 39200 10080 40000 10192 0 FreeSans 448 0 0 0 proj_out[10]
port 13 nsew signal input
flabel metal3 s 39200 13440 40000 13552 0 FreeSans 448 0 0 0 proj_out[11]
port 14 nsew signal input
flabel metal3 s 39200 24192 40000 24304 0 FreeSans 448 0 0 0 proj_out[12]
port 15 nsew signal input
flabel metal2 s 26880 39200 26992 40000 0 FreeSans 448 90 0 0 proj_out[13]
port 16 nsew signal input
flabel metal2 s 24192 39200 24304 40000 0 FreeSans 448 90 0 0 proj_out[14]
port 17 nsew signal input
flabel metal3 s 39200 26880 40000 26992 0 FreeSans 448 0 0 0 proj_out[15]
port 18 nsew signal input
flabel metal3 s 39200 22176 40000 22288 0 FreeSans 448 0 0 0 proj_out[16]
port 19 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 proj_out[17]
port 20 nsew signal input
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 proj_out[18]
port 21 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 proj_out[19]
port 22 nsew signal input
flabel metal2 s 26208 39200 26320 40000 0 FreeSans 448 90 0 0 proj_out[1]
port 23 nsew signal input
flabel metal3 s 39200 19488 40000 19600 0 FreeSans 448 0 0 0 proj_out[20]
port 24 nsew signal input
flabel metal3 s 39200 12768 40000 12880 0 FreeSans 448 0 0 0 proj_out[21]
port 25 nsew signal input
flabel metal3 s 39200 12096 40000 12208 0 FreeSans 448 0 0 0 proj_out[22]
port 26 nsew signal input
flabel metal3 s 39200 16800 40000 16912 0 FreeSans 448 0 0 0 proj_out[23]
port 27 nsew signal input
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 proj_out[24]
port 28 nsew signal input
flabel metal2 s 14112 39200 14224 40000 0 FreeSans 448 90 0 0 proj_out[25]
port 29 nsew signal input
flabel metal2 s 14784 39200 14896 40000 0 FreeSans 448 90 0 0 proj_out[26]
port 30 nsew signal input
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 proj_out[27]
port 31 nsew signal input
flabel metal2 s 21504 39200 21616 40000 0 FreeSans 448 90 0 0 proj_out[28]
port 32 nsew signal input
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 proj_out[29]
port 33 nsew signal input
flabel metal2 s 25536 39200 25648 40000 0 FreeSans 448 90 0 0 proj_out[2]
port 34 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 proj_out[30]
port 35 nsew signal input
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 proj_out[31]
port 36 nsew signal input
flabel metal3 s 0 14112 800 14224 0 FreeSans 448 0 0 0 proj_out[32]
port 37 nsew signal input
flabel metal3 s 0 14784 800 14896 0 FreeSans 448 0 0 0 proj_out[33]
port 38 nsew signal input
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 proj_out[34]
port 39 nsew signal input
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 proj_out[35]
port 40 nsew signal input
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 proj_out[36]
port 41 nsew signal input
flabel metal2 s 15456 39200 15568 40000 0 FreeSans 448 90 0 0 proj_out[37]
port 42 nsew signal input
flabel metal2 s 12768 39200 12880 40000 0 FreeSans 448 90 0 0 proj_out[38]
port 43 nsew signal input
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 proj_out[39]
port 44 nsew signal input
flabel metal3 s 39200 28224 40000 28336 0 FreeSans 448 0 0 0 proj_out[3]
port 45 nsew signal input
flabel metal3 s 39200 20832 40000 20944 0 FreeSans 448 0 0 0 proj_out[40]
port 46 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 proj_out[41]
port 47 nsew signal input
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 proj_out[42]
port 48 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 proj_out[43]
port 49 nsew signal input
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 proj_out[44]
port 50 nsew signal input
flabel metal3 s 0 13440 800 13552 0 FreeSans 448 0 0 0 proj_out[45]
port 51 nsew signal input
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 proj_out[46]
port 52 nsew signal input
flabel metal3 s 0 12768 800 12880 0 FreeSans 448 0 0 0 proj_out[47]
port 53 nsew signal input
flabel metal3 s 39200 27552 40000 27664 0 FreeSans 448 0 0 0 proj_out[48]
port 54 nsew signal input
flabel metal2 s 24864 39200 24976 40000 0 FreeSans 448 90 0 0 proj_out[49]
port 55 nsew signal input
flabel metal3 s 39200 21504 40000 21616 0 FreeSans 448 0 0 0 proj_out[4]
port 56 nsew signal input
flabel metal2 s 22176 39200 22288 40000 0 FreeSans 448 90 0 0 proj_out[50]
port 57 nsew signal input
flabel metal3 s 39200 28896 40000 29008 0 FreeSans 448 0 0 0 proj_out[51]
port 58 nsew signal input
flabel metal3 s 39200 23520 40000 23632 0 FreeSans 448 0 0 0 proj_out[52]
port 59 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 proj_out[53]
port 60 nsew signal input
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 proj_out[54]
port 61 nsew signal input
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 proj_out[55]
port 62 nsew signal input
flabel metal3 s 39200 20160 40000 20272 0 FreeSans 448 0 0 0 proj_out[56]
port 63 nsew signal input
flabel metal3 s 39200 11424 40000 11536 0 FreeSans 448 0 0 0 proj_out[57]
port 64 nsew signal input
flabel metal3 s 39200 10752 40000 10864 0 FreeSans 448 0 0 0 proj_out[58]
port 65 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 proj_out[59]
port 66 nsew signal input
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 proj_out[5]
port 67 nsew signal input
flabel metal3 s 39200 25536 40000 25648 0 FreeSans 448 0 0 0 proj_out[60]
port 68 nsew signal input
flabel metal2 s 22848 39200 22960 40000 0 FreeSans 448 90 0 0 proj_out[61]
port 69 nsew signal input
flabel metal2 s 23520 39200 23632 40000 0 FreeSans 448 90 0 0 proj_out[62]
port 70 nsew signal input
flabel metal3 s 39200 24864 40000 24976 0 FreeSans 448 0 0 0 proj_out[63]
port 71 nsew signal input
flabel metal3 s 39200 29568 40000 29680 0 FreeSans 448 0 0 0 proj_out[64]
port 72 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 proj_out[65]
port 73 nsew signal input
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 proj_out[66]
port 74 nsew signal input
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 proj_out[67]
port 75 nsew signal input
flabel metal3 s 39200 18816 40000 18928 0 FreeSans 448 0 0 0 proj_out[68]
port 76 nsew signal input
flabel metal3 s 39200 15456 40000 15568 0 FreeSans 448 0 0 0 proj_out[69]
port 77 nsew signal input
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 proj_out[6]
port 78 nsew signal input
flabel metal3 s 39200 14784 40000 14896 0 FreeSans 448 0 0 0 proj_out[70]
port 79 nsew signal input
flabel metal3 s 39200 16128 40000 16240 0 FreeSans 448 0 0 0 proj_out[71]
port 80 nsew signal input
flabel metal2 s 19488 39200 19600 40000 0 FreeSans 448 90 0 0 proj_out[72]
port 81 nsew signal input
flabel metal2 s 16800 39200 16912 40000 0 FreeSans 448 90 0 0 proj_out[73]
port 82 nsew signal input
flabel metal2 s 11424 39200 11536 40000 0 FreeSans 448 90 0 0 proj_out[74]
port 83 nsew signal input
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 proj_out[75]
port 84 nsew signal input
flabel metal2 s 18816 39200 18928 40000 0 FreeSans 448 90 0 0 proj_out[76]
port 85 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 proj_out[77]
port 86 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 proj_out[78]
port 87 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 proj_out[79]
port 88 nsew signal input
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 proj_out[7]
port 89 nsew signal input
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 proj_out[80]
port 90 nsew signal input
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 proj_out[81]
port 91 nsew signal input
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 proj_out[82]
port 92 nsew signal input
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 proj_out[83]
port 93 nsew signal input
flabel metal2 s 18144 39200 18256 40000 0 FreeSans 448 90 0 0 proj_out[84]
port 94 nsew signal input
flabel metal2 s 13440 39200 13552 40000 0 FreeSans 448 90 0 0 proj_out[85]
port 95 nsew signal input
flabel metal2 s 12096 39200 12208 40000 0 FreeSans 448 90 0 0 proj_out[86]
port 96 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 proj_out[87]
port 97 nsew signal input
flabel metal2 s 17472 39200 17584 40000 0 FreeSans 448 90 0 0 proj_out[88]
port 98 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 proj_out[89]
port 99 nsew signal input
flabel metal3 s 39200 18144 40000 18256 0 FreeSans 448 0 0 0 proj_out[8]
port 100 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 proj_out[90]
port 101 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 proj_out[91]
port 102 nsew signal input
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 proj_out[92]
port 103 nsew signal input
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 proj_out[93]
port 104 nsew signal input
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 proj_out[94]
port 105 nsew signal input
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 proj_out[95]
port 106 nsew signal input
flabel metal3 s 39200 14112 40000 14224 0 FreeSans 448 0 0 0 proj_out[9]
port 107 nsew signal input
flabel metal3 s 39200 22848 40000 22960 0 FreeSans 448 0 0 0 sel[0]
port 108 nsew signal input
flabel metal3 s 39200 26208 40000 26320 0 FreeSans 448 0 0 0 sel[1]
port 109 nsew signal input
flabel metal3 s 39200 17472 40000 17584 0 FreeSans 448 0 0 0 sel[2]
port 110 nsew signal input
flabel metal4 s 5846 3076 6166 36908 0 FreeSans 1280 90 0 0 vdd
port 111 nsew power bidirectional
flabel metal4 s 15170 3076 15490 36908 0 FreeSans 1280 90 0 0 vdd
port 111 nsew power bidirectional
flabel metal4 s 24494 3076 24814 36908 0 FreeSans 1280 90 0 0 vdd
port 111 nsew power bidirectional
flabel metal4 s 33818 3076 34138 36908 0 FreeSans 1280 90 0 0 vdd
port 111 nsew power bidirectional
flabel metal4 s 10508 3076 10828 36908 0 FreeSans 1280 90 0 0 vss
port 112 nsew ground bidirectional
flabel metal4 s 19832 3076 20152 36908 0 FreeSans 1280 90 0 0 vss
port 112 nsew ground bidirectional
flabel metal4 s 29156 3076 29476 36908 0 FreeSans 1280 90 0 0 vss
port 112 nsew ground bidirectional
flabel metal4 s 38480 3076 38800 36908 0 FreeSans 1280 90 0 0 vss
port 112 nsew ground bidirectional
rlabel metal1 19992 36848 19992 36848 0 vdd
rlabel via1 20072 36064 20072 36064 0 vss
rlabel metal2 20328 19656 20328 19656 0 _000_
rlabel metal2 21000 21672 21000 21672 0 _001_
rlabel metal2 21448 25480 21448 25480 0 _002_
rlabel metal2 25256 20860 25256 20860 0 _003_
rlabel metal2 25816 22344 25816 22344 0 _004_
rlabel metal2 23352 21644 23352 21644 0 _005_
rlabel metal2 27048 23912 27048 23912 0 _006_
rlabel metal3 24024 23352 24024 23352 0 _007_
rlabel metal2 21168 23912 21168 23912 0 _008_
rlabel metal3 20776 22120 20776 22120 0 _009_
rlabel metal2 13160 23072 13160 23072 0 _010_
rlabel metal3 21056 26152 21056 26152 0 _011_
rlabel metal2 18536 21224 18536 21224 0 _012_
rlabel metal2 18760 25480 18760 25480 0 _013_
rlabel metal2 21448 18424 21448 18424 0 _014_
rlabel metal2 21336 20552 21336 20552 0 _015_
rlabel metal2 16856 22400 16856 22400 0 _016_
rlabel metal2 20328 25480 20328 25480 0 _017_
rlabel metal2 19880 27608 19880 27608 0 _018_
rlabel metal2 22344 17248 22344 17248 0 _019_
rlabel metal2 17864 21644 17864 21644 0 _020_
rlabel metal2 15624 23688 15624 23688 0 _021_
rlabel metal2 14728 25984 14728 25984 0 _022_
rlabel metal2 15064 27160 15064 27160 0 _023_
rlabel metal2 24304 21336 24304 21336 0 _024_
rlabel metal2 12600 25816 12600 25816 0 _025_
rlabel metal3 17864 25256 17864 25256 0 _026_
rlabel metal2 15624 25872 15624 25872 0 _027_
rlabel metal3 16968 23912 16968 23912 0 _028_
rlabel metal3 22232 25368 22232 25368 0 _029_
rlabel metal2 20216 25088 20216 25088 0 _030_
rlabel metal2 19656 24192 19656 24192 0 _031_
rlabel metal2 18424 25480 18424 25480 0 _032_
rlabel metal2 16520 25536 16520 25536 0 _033_
rlabel metal2 22736 23688 22736 23688 0 _034_
rlabel metal2 20104 25928 20104 25928 0 _035_
rlabel metal2 19656 25760 19656 25760 0 _036_
rlabel metal3 13944 24696 13944 24696 0 _037_
rlabel metal2 14616 24360 14616 24360 0 _038_
rlabel metal2 25816 24696 25816 24696 0 _039_
rlabel metal3 24808 24808 24808 24808 0 _040_
rlabel metal3 19488 24808 19488 24808 0 _041_
rlabel metal2 15848 21560 15848 21560 0 _042_
rlabel metal2 13608 21168 13608 21168 0 _043_
rlabel metal2 14560 23016 14560 23016 0 _044_
rlabel metal2 15736 23016 15736 23016 0 _045_
rlabel metal2 18984 21112 18984 21112 0 _046_
rlabel metal3 22232 19992 22232 19992 0 _047_
rlabel metal2 23968 21672 23968 21672 0 _048_
rlabel metal2 22680 19880 22680 19880 0 _049_
rlabel metal2 21560 19208 21560 19208 0 _050_
rlabel metal2 22064 21560 22064 21560 0 _051_
rlabel metal2 22288 22120 22288 22120 0 _052_
rlabel metal2 21112 21896 21112 21896 0 _053_
rlabel metal2 20104 21112 20104 21112 0 _054_
rlabel metal3 23128 20608 23128 20608 0 _055_
rlabel metal3 23912 20328 23912 20328 0 _056_
rlabel metal2 22120 20272 22120 20272 0 _057_
rlabel metal3 20720 20776 20720 20776 0 _058_
rlabel metal2 20216 22064 20216 22064 0 _059_
rlabel metal2 18088 16968 18088 16968 0 _060_
rlabel metal2 21224 15344 21224 15344 0 _061_
rlabel metal3 20832 15288 20832 15288 0 _062_
rlabel metal3 20888 17080 20888 17080 0 _063_
rlabel metal2 21896 16968 21896 16968 0 _064_
rlabel metal2 21224 13328 21224 13328 0 _065_
rlabel metal3 18144 16072 18144 16072 0 _066_
rlabel metal2 20776 12432 20776 12432 0 _067_
rlabel metal2 20272 16856 20272 16856 0 _068_
rlabel metal2 21112 12992 21112 12992 0 _069_
rlabel metal2 19208 14392 19208 14392 0 _070_
rlabel metal2 22008 13104 22008 13104 0 _071_
rlabel metal3 20272 12376 20272 12376 0 _072_
rlabel metal2 21840 13048 21840 13048 0 _073_
rlabel metal3 20384 14840 20384 14840 0 _074_
rlabel metal3 23800 12768 23800 12768 0 _075_
rlabel metal3 18648 13608 18648 13608 0 _076_
rlabel metal3 20104 13944 20104 13944 0 _077_
rlabel metal2 12936 19376 12936 19376 0 _078_
rlabel metal3 13160 17640 13160 17640 0 _079_
rlabel metal2 14952 17976 14952 17976 0 _080_
rlabel metal2 14840 18200 14840 18200 0 _081_
rlabel metal3 18816 17528 18816 17528 0 _082_
rlabel metal2 24248 17136 24248 17136 0 _083_
rlabel metal3 22456 19096 22456 19096 0 _084_
rlabel metal2 18200 19656 18200 19656 0 _085_
rlabel metal2 17416 20580 17416 20580 0 _086_
rlabel metal3 13944 16856 13944 16856 0 _087_
rlabel metal2 14616 16072 14616 16072 0 _088_
rlabel metal2 26936 17136 26936 17136 0 _089_
rlabel metal2 16296 17192 16296 17192 0 _090_
rlabel metal2 15736 18312 15736 18312 0 _091_
rlabel metal2 14504 17304 14504 17304 0 _092_
rlabel metal3 13160 17864 13160 17864 0 _093_
rlabel metal2 26376 17584 26376 17584 0 _094_
rlabel metal2 19656 17752 19656 17752 0 _095_
rlabel metal2 15624 18872 15624 18872 0 _096_
rlabel metal2 16408 16520 16408 16520 0 _097_
rlabel metal2 15624 16968 15624 16968 0 _098_
rlabel metal2 18536 16520 18536 16520 0 _099_
rlabel metal2 18200 16800 18200 16800 0 _100_
rlabel metal2 17752 20048 17752 20048 0 _101_
rlabel metal3 28504 23184 28504 23184 0 net1
rlabel metal2 27272 3584 27272 3584 0 net10
rlabel metal2 20552 31864 20552 31864 0 net100
rlabel metal3 10136 12152 10136 12152 0 net101
rlabel metal2 4312 12992 4312 12992 0 net102
rlabel metal3 15624 24136 15624 24136 0 net103
rlabel metal2 19208 31024 19208 31024 0 net104
rlabel metal2 15904 24472 15904 24472 0 net105
rlabel metal2 20720 21000 20720 21000 0 net106
rlabel metal3 20272 15176 20272 15176 0 net107
rlabel metal2 15792 3528 15792 3528 0 net108
rlabel metal2 22904 6216 22904 6216 0 net109
rlabel metal2 29736 3920 29736 3920 0 net11
rlabel metal3 6356 19208 6356 19208 0 net110
rlabel metal2 4312 17136 4312 17136 0 net111
rlabel metal2 27496 34888 27496 34888 0 net12
rlabel metal2 37016 19656 37016 19656 0 net13
rlabel metal2 28168 14896 28168 14896 0 net14
rlabel metal2 27384 15232 27384 15232 0 net15
rlabel metal2 23688 16968 23688 16968 0 net16
rlabel metal2 2072 27104 2072 27104 0 net17
rlabel metal2 14392 32704 14392 32704 0 net18
rlabel metal2 15064 32536 15064 32536 0 net19
rlabel metal2 28504 14168 28504 14168 0 net2
rlabel metal2 2744 25424 2744 25424 0 net20
rlabel metal2 20608 27272 20608 27272 0 net21
rlabel metal2 20104 12768 20104 12768 0 net22
rlabel metal3 25816 36232 25816 36232 0 net23
rlabel metal2 19824 3416 19824 3416 0 net24
rlabel metal2 20104 13440 20104 13440 0 net25
rlabel metal2 2016 14392 2016 14392 0 net26
rlabel metal3 5236 15400 5236 15400 0 net27
rlabel metal2 2744 17360 2744 17360 0 net28
rlabel metal2 15400 16016 15400 16016 0 net29
rlabel metal2 24752 16856 24752 16856 0 net3
rlabel metal2 14392 26040 14392 26040 0 net30
rlabel metal2 16296 28224 16296 28224 0 net31
rlabel metal2 12600 31696 12600 31696 0 net32
rlabel metal2 12376 24976 12376 24976 0 net33
rlabel metal2 28728 26712 28728 26712 0 net34
rlabel metal2 23464 20720 23464 20720 0 net35
rlabel metal2 12656 3416 12656 3416 0 net36
rlabel metal2 15400 5152 15400 5152 0 net37
rlabel metal2 14728 9072 14728 9072 0 net38
rlabel metal2 12264 19712 12264 19712 0 net39
rlabel metal2 27720 23016 27720 23016 0 net4
rlabel metal2 2128 13944 2128 13944 0 net40
rlabel metal2 2072 16632 2072 16632 0 net41
rlabel metal3 9240 13832 9240 13832 0 net42
rlabel metal2 38360 25144 38360 25144 0 net43
rlabel metal3 23856 32312 23856 32312 0 net44
rlabel metal2 37296 22120 37296 22120 0 net45
rlabel metal2 21952 24024 21952 24024 0 net46
rlabel metal2 37464 27048 37464 27048 0 net47
rlabel metal3 27160 20832 27160 20832 0 net48
rlabel metal2 24416 3416 24416 3416 0 net49
rlabel metal2 27160 34608 27160 34608 0 net5
rlabel metal2 23688 4144 23688 4144 0 net50
rlabel metal2 25256 4200 25256 4200 0 net51
rlabel metal3 27664 20216 27664 20216 0 net52
rlabel metal2 25984 16744 25984 16744 0 net53
rlabel metal3 27328 17528 27328 17528 0 net54
rlabel metal3 21672 4536 21672 4536 0 net55
rlabel metal2 28336 3416 28336 3416 0 net56
rlabel metal2 26376 23800 26376 23800 0 net57
rlabel metal2 22680 26180 22680 26180 0 net58
rlabel metal3 23408 35672 23408 35672 0 net59
rlabel metal2 24136 25396 24136 25396 0 net6
rlabel metal2 26488 24976 26488 24976 0 net60
rlabel metal2 24024 20608 24024 20608 0 net61
rlabel metal2 23688 13832 23688 13832 0 net62
rlabel metal2 30408 8512 30408 8512 0 net63
rlabel metal2 23688 11648 23688 11648 0 net64
rlabel metal3 26264 19264 26264 19264 0 net65
rlabel metal2 26824 16352 26824 16352 0 net66
rlabel metal2 24920 9128 24920 9128 0 net67
rlabel metal2 26376 16240 26376 16240 0 net68
rlabel metal2 22344 16800 22344 16800 0 net69
rlabel metal2 37016 25760 37016 25760 0 net7
rlabel metal2 20216 31640 20216 31640 0 net70
rlabel metal3 21000 24640 21000 24640 0 net71
rlabel metal3 20580 26264 20580 26264 0 net72
rlabel metal2 2632 24640 2632 24640 0 net73
rlabel metal2 20440 22848 20440 22848 0 net74
rlabel metal2 20888 15064 20888 15064 0 net75
rlabel metal2 18424 9240 18424 9240 0 net76
rlabel metal2 18816 16072 18816 16072 0 net77
rlabel metal2 29064 4144 29064 4144 0 net78
rlabel metal2 2296 22680 2296 22680 0 net79
rlabel metal2 37632 21112 37632 21112 0 net8
rlabel metal2 2128 20552 2128 20552 0 net80
rlabel metal2 2072 18480 2072 18480 0 net81
rlabel metal2 2072 22288 2072 22288 0 net82
rlabel metal2 18760 31416 18760 31416 0 net83
rlabel metal3 15904 24920 15904 24920 0 net84
rlabel metal2 19544 26572 19544 26572 0 net85
rlabel metal3 12376 23632 12376 23632 0 net86
rlabel metal2 19264 23128 19264 23128 0 net87
rlabel metal3 20832 14616 20832 14616 0 net88
rlabel metal2 28504 19096 28504 19096 0 net89
rlabel metal2 31080 8960 31080 8960 0 net9
rlabel metal2 18984 12152 18984 12152 0 net90
rlabel metal3 17528 4648 17528 4648 0 net91
rlabel metal2 2856 24472 2856 24472 0 net92
rlabel metal2 12264 21392 12264 21392 0 net93
rlabel metal2 2744 20720 2744 20720 0 net94
rlabel metal3 5236 23240 5236 23240 0 net95
rlabel metal2 29064 15568 29064 15568 0 net96
rlabel metal2 25816 20328 25816 20328 0 net97
rlabel metal2 28280 20944 28280 20944 0 net98
rlabel metal2 22568 18368 22568 18368 0 net99
rlabel metal2 20216 38066 20216 38066 0 out[0]
rlabel metal3 1358 11480 1358 11480 0 out[10]
rlabel metal3 1358 12152 1358 12152 0 out[11]
rlabel metal2 10808 38066 10808 38066 0 out[1]
rlabel metal3 16688 36680 16688 36680 0 out[2]
rlabel metal3 1358 28952 1358 28952 0 out[3]
rlabel metal2 20888 37954 20888 37954 0 out[4]
rlabel metal2 12152 854 12152 854 0 out[5]
rlabel metal2 12824 854 12824 854 0 out[6]
rlabel metal3 20272 3640 20272 3640 0 out[7]
rlabel metal3 1358 18872 1358 18872 0 out[8]
rlabel metal3 1358 17528 1358 17528 0 out[9]
rlabel metal2 38248 30632 38248 30632 0 proj_out[0]
rlabel metal2 38248 10360 38248 10360 0 proj_out[10]
rlabel metal2 38248 13608 38248 13608 0 proj_out[11]
rlabel metal2 38248 24472 38248 24472 0 proj_out[12]
rlabel metal2 26992 35896 26992 35896 0 proj_out[13]
rlabel metal2 25480 36568 25480 36568 0 proj_out[14]
rlabel metal3 38290 26936 38290 26936 0 proj_out[15]
rlabel metal3 38738 22232 38738 22232 0 proj_out[16]
rlabel metal2 31304 2128 31304 2128 0 proj_out[17]
rlabel metal2 27944 3864 27944 3864 0 proj_out[18]
rlabel metal2 29960 3192 29960 3192 0 proj_out[19]
rlabel metal2 27496 36680 27496 36680 0 proj_out[1]
rlabel metal2 38248 19768 38248 19768 0 proj_out[20]
rlabel metal3 38738 12824 38738 12824 0 proj_out[21]
rlabel metal3 38402 12152 38402 12152 0 proj_out[22]
rlabel metal3 38024 16968 38024 16968 0 proj_out[23]
rlabel metal2 1848 26656 1848 26656 0 proj_out[24]
rlabel metal2 14168 37842 14168 37842 0 proj_out[25]
rlabel metal2 14840 37842 14840 37842 0 proj_out[26]
rlabel metal3 1582 26936 1582 26936 0 proj_out[27]
rlabel metal2 21560 37114 21560 37114 0 proj_out[28]
rlabel metal2 20664 2856 20664 2856 0 proj_out[29]
rlabel metal2 26824 36568 26824 36568 0 proj_out[2]
rlabel metal2 20216 2058 20216 2058 0 proj_out[30]
rlabel metal3 21448 4312 21448 4312 0 proj_out[31]
rlabel metal2 1736 14280 1736 14280 0 proj_out[32]
rlabel metal2 1736 15064 1736 15064 0 proj_out[33]
rlabel metal2 2408 16520 2408 16520 0 proj_out[34]
rlabel metal2 1736 15736 1736 15736 0 proj_out[35]
rlabel metal2 1736 25928 1736 25928 0 proj_out[36]
rlabel metal2 15568 36456 15568 36456 0 proj_out[37]
rlabel metal2 12600 36456 12600 36456 0 proj_out[38]
rlabel metal2 1736 25144 1736 25144 0 proj_out[39]
rlabel metal3 38528 28616 38528 28616 0 proj_out[3]
rlabel metal2 38248 21224 38248 21224 0 proj_out[40]
rlabel metal2 12376 3472 12376 3472 0 proj_out[41]
rlabel metal2 14952 5096 14952 5096 0 proj_out[42]
rlabel metal2 14392 4648 14392 4648 0 proj_out[43]
rlabel metal2 1736 19768 1736 19768 0 proj_out[44]
rlabel metal2 1736 13608 1736 13608 0 proj_out[45]
rlabel metal3 1246 16856 1246 16856 0 proj_out[46]
rlabel metal2 2408 13272 2408 13272 0 proj_out[47]
rlabel metal2 38248 27720 38248 27720 0 proj_out[48]
rlabel metal3 26264 36512 26264 36512 0 proj_out[49]
rlabel metal3 38402 21560 38402 21560 0 proj_out[4]
rlabel metal2 23576 35728 23576 35728 0 proj_out[50]
rlabel metal2 38248 29176 38248 29176 0 proj_out[51]
rlabel metal2 38248 23744 38248 23744 0 proj_out[52]
rlabel metal2 24192 2520 24192 2520 0 proj_out[53]
rlabel metal2 22904 2058 22904 2058 0 proj_out[54]
rlabel metal2 24584 2296 24584 2296 0 proj_out[55]
rlabel metal2 38248 20440 38248 20440 0 proj_out[56]
rlabel metal2 38248 11816 38248 11816 0 proj_out[57]
rlabel metal2 38248 11032 38248 11032 0 proj_out[58]
rlabel metal2 22680 4592 22680 4592 0 proj_out[59]
rlabel metal2 28616 3472 28616 3472 0 proj_out[5]
rlabel metal2 38248 25928 38248 25928 0 proj_out[60]
rlabel metal3 23856 36456 23856 36456 0 proj_out[61]
rlabel metal2 24248 36120 24248 36120 0 proj_out[62]
rlabel metal2 38248 25144 38248 25144 0 proj_out[63]
rlabel metal2 38248 29848 38248 29848 0 proj_out[64]
rlabel metal2 26824 3808 26824 3808 0 proj_out[65]
rlabel metal2 30632 3472 30632 3472 0 proj_out[66]
rlabel metal2 24976 2184 24976 2184 0 proj_out[67]
rlabel metal2 38248 19040 38248 19040 0 proj_out[68]
rlabel metal2 38248 15736 38248 15736 0 proj_out[69]
rlabel metal2 26992 4200 26992 4200 0 proj_out[6]
rlabel metal2 38248 15064 38248 15064 0 proj_out[70]
rlabel metal2 38248 16520 38248 16520 0 proj_out[71]
rlabel metal2 19880 36736 19880 36736 0 proj_out[72]
rlabel via2 16520 36456 16520 36456 0 proj_out[73]
rlabel metal2 11032 36792 11032 36792 0 proj_out[74]
rlabel metal2 1736 27720 1736 27720 0 proj_out[75]
rlabel metal2 18984 35784 18984 35784 0 proj_out[76]
rlabel metal2 15512 2058 15512 2058 0 proj_out[77]
rlabel metal3 18424 3528 18424 3528 0 proj_out[78]
rlabel metal2 17528 2058 17528 2058 0 proj_out[79]
rlabel metal3 29400 3472 29400 3472 0 proj_out[7]
rlabel metal2 1736 24472 1736 24472 0 proj_out[80]
rlabel metal2 1736 20384 1736 20384 0 proj_out[81]
rlabel metal2 1736 18312 1736 18312 0 proj_out[82]
rlabel metal3 1246 22232 1246 22232 0 proj_out[83]
rlabel metal2 18312 35784 18312 35784 0 proj_out[84]
rlabel metal2 13496 37842 13496 37842 0 proj_out[85]
rlabel metal2 11760 36456 11760 36456 0 proj_out[86]
rlabel metal2 1736 23632 1736 23632 0 proj_out[87]
rlabel metal2 17640 35784 17640 35784 0 proj_out[88]
rlabel metal2 16968 3528 16968 3528 0 proj_out[89]
rlabel metal2 38248 18312 38248 18312 0 proj_out[8]
rlabel metal2 19096 2520 19096 2520 0 proj_out[90]
rlabel metal2 16408 4872 16408 4872 0 proj_out[91]
rlabel metal2 1736 28448 1736 28448 0 proj_out[92]
rlabel metal2 1736 21224 1736 21224 0 proj_out[93]
rlabel metal2 2408 21840 2408 21840 0 proj_out[94]
rlabel metal2 1736 23016 1736 23016 0 proj_out[95]
rlabel metal2 38248 14336 38248 14336 0 proj_out[9]
rlabel metal2 38248 23016 38248 23016 0 sel[0]
rlabel metal2 38136 26656 38136 26656 0 sel[1]
rlabel metal3 38738 17528 38738 17528 0 sel[2]
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
