magic
tech gf180mcuD
magscale 1 10
timestamp 1702441332
<< metal1 >>
rect 32274 37774 32286 37826
rect 32338 37823 32350 37826
rect 33506 37823 33518 37826
rect 32338 37777 33518 37823
rect 32338 37774 32350 37777
rect 33506 37774 33518 37777
rect 33570 37774 33582 37826
rect 33618 37662 33630 37714
rect 33682 37711 33694 37714
rect 34850 37711 34862 37714
rect 33682 37665 34862 37711
rect 33682 37662 33694 37665
rect 34850 37662 34862 37665
rect 34914 37662 34926 37714
rect 1344 36874 38640 36908
rect 1344 36822 5876 36874
rect 5928 36822 5980 36874
rect 6032 36822 6084 36874
rect 6136 36822 15200 36874
rect 15252 36822 15304 36874
rect 15356 36822 15408 36874
rect 15460 36822 24524 36874
rect 24576 36822 24628 36874
rect 24680 36822 24732 36874
rect 24784 36822 33848 36874
rect 33900 36822 33952 36874
rect 34004 36822 34056 36874
rect 34108 36822 38640 36874
rect 1344 36788 38640 36822
rect 5742 36482 5794 36494
rect 2706 36430 2718 36482
rect 2770 36430 2782 36482
rect 4050 36430 4062 36482
rect 4114 36430 4126 36482
rect 4834 36430 4846 36482
rect 4898 36430 4910 36482
rect 6514 36430 6526 36482
rect 6578 36430 6590 36482
rect 7858 36430 7870 36482
rect 7922 36430 7934 36482
rect 9650 36430 9662 36482
rect 9714 36430 9726 36482
rect 10322 36430 10334 36482
rect 10386 36430 10398 36482
rect 10994 36430 11006 36482
rect 11058 36430 11070 36482
rect 11666 36430 11678 36482
rect 11730 36430 11742 36482
rect 14802 36430 14814 36482
rect 14866 36430 14878 36482
rect 15474 36430 15486 36482
rect 15538 36430 15550 36482
rect 17266 36430 17278 36482
rect 17330 36430 17342 36482
rect 17938 36430 17950 36482
rect 18002 36430 18014 36482
rect 19282 36430 19294 36482
rect 19346 36430 19358 36482
rect 22642 36430 22654 36482
rect 22706 36430 22718 36482
rect 23314 36430 23326 36482
rect 23378 36430 23390 36482
rect 25442 36430 25454 36482
rect 25506 36430 25518 36482
rect 26786 36430 26798 36482
rect 26850 36430 26862 36482
rect 27458 36430 27470 36482
rect 27522 36430 27534 36482
rect 29250 36430 29262 36482
rect 29314 36430 29326 36482
rect 32386 36430 32398 36482
rect 32450 36430 32462 36482
rect 33058 36430 33070 36482
rect 33122 36430 33134 36482
rect 34402 36430 34414 36482
rect 34466 36430 34478 36482
rect 36194 36430 36206 36482
rect 36258 36430 36270 36482
rect 36866 36430 36878 36482
rect 36930 36430 36942 36482
rect 37538 36430 37550 36482
rect 37602 36430 37614 36482
rect 5742 36418 5794 36430
rect 3278 36370 3330 36382
rect 3278 36306 3330 36318
rect 3614 36370 3666 36382
rect 3614 36306 3666 36318
rect 4622 36370 4674 36382
rect 4622 36306 4674 36318
rect 7086 36370 7138 36382
rect 7086 36306 7138 36318
rect 7422 36370 7474 36382
rect 7422 36306 7474 36318
rect 8094 36370 8146 36382
rect 8094 36306 8146 36318
rect 8430 36370 8482 36382
rect 8430 36306 8482 36318
rect 8766 36370 8818 36382
rect 8766 36306 8818 36318
rect 9886 36370 9938 36382
rect 9886 36306 9938 36318
rect 10558 36370 10610 36382
rect 10558 36306 10610 36318
rect 11230 36370 11282 36382
rect 11230 36306 11282 36318
rect 11902 36370 11954 36382
rect 11902 36306 11954 36318
rect 12238 36370 12290 36382
rect 12238 36306 12290 36318
rect 12574 36370 12626 36382
rect 12574 36306 12626 36318
rect 13358 36370 13410 36382
rect 13358 36306 13410 36318
rect 13694 36370 13746 36382
rect 13694 36306 13746 36318
rect 14030 36370 14082 36382
rect 14030 36306 14082 36318
rect 14366 36370 14418 36382
rect 14366 36306 14418 36318
rect 16046 36370 16098 36382
rect 16046 36306 16098 36318
rect 16382 36370 16434 36382
rect 16382 36306 16434 36318
rect 17502 36370 17554 36382
rect 17502 36306 17554 36318
rect 18174 36370 18226 36382
rect 18174 36306 18226 36318
rect 18510 36370 18562 36382
rect 18510 36306 18562 36318
rect 18846 36370 18898 36382
rect 18846 36306 18898 36318
rect 19518 36370 19570 36382
rect 19518 36306 19570 36318
rect 19854 36370 19906 36382
rect 19854 36306 19906 36318
rect 20190 36370 20242 36382
rect 20190 36306 20242 36318
rect 21086 36370 21138 36382
rect 21086 36306 21138 36318
rect 21422 36370 21474 36382
rect 21422 36306 21474 36318
rect 21758 36370 21810 36382
rect 21758 36306 21810 36318
rect 22094 36370 22146 36382
rect 22094 36306 22146 36318
rect 22430 36370 22482 36382
rect 22430 36306 22482 36318
rect 23102 36370 23154 36382
rect 23102 36306 23154 36318
rect 24558 36370 24610 36382
rect 24558 36306 24610 36318
rect 24894 36370 24946 36382
rect 24894 36306 24946 36318
rect 25230 36370 25282 36382
rect 25230 36306 25282 36318
rect 25902 36370 25954 36382
rect 25902 36306 25954 36318
rect 26238 36370 26290 36382
rect 26238 36306 26290 36318
rect 26574 36370 26626 36382
rect 26574 36306 26626 36318
rect 27246 36370 27298 36382
rect 27246 36306 27298 36318
rect 28366 36370 28418 36382
rect 28366 36306 28418 36318
rect 28702 36370 28754 36382
rect 28702 36306 28754 36318
rect 29710 36370 29762 36382
rect 29710 36306 29762 36318
rect 30046 36370 30098 36382
rect 30046 36306 30098 36318
rect 30718 36370 30770 36382
rect 30718 36306 30770 36318
rect 31054 36370 31106 36382
rect 31054 36306 31106 36318
rect 31390 36370 31442 36382
rect 31390 36306 31442 36318
rect 32174 36370 32226 36382
rect 32174 36306 32226 36318
rect 32846 36370 32898 36382
rect 32846 36306 32898 36318
rect 33518 36370 33570 36382
rect 33518 36306 33570 36318
rect 33854 36370 33906 36382
rect 33854 36306 33906 36318
rect 34190 36370 34242 36382
rect 34190 36306 34242 36318
rect 34862 36370 34914 36382
rect 34862 36306 34914 36318
rect 35198 36370 35250 36382
rect 35198 36306 35250 36318
rect 35982 36370 36034 36382
rect 35982 36306 36034 36318
rect 36654 36370 36706 36382
rect 36654 36306 36706 36318
rect 37326 36370 37378 36382
rect 37326 36306 37378 36318
rect 4286 36258 4338 36270
rect 2930 36206 2942 36258
rect 2994 36206 3006 36258
rect 4286 36194 4338 36206
rect 6078 36258 6130 36270
rect 6078 36194 6130 36206
rect 6750 36258 6802 36270
rect 6750 36194 6802 36206
rect 15038 36258 15090 36270
rect 15038 36194 15090 36206
rect 15710 36258 15762 36270
rect 15710 36194 15762 36206
rect 29038 36258 29090 36270
rect 29038 36194 29090 36206
rect 30382 36258 30434 36270
rect 30382 36194 30434 36206
rect 38110 36258 38162 36270
rect 38110 36194 38162 36206
rect 1344 36090 38800 36124
rect 1344 36038 10538 36090
rect 10590 36038 10642 36090
rect 10694 36038 10746 36090
rect 10798 36038 19862 36090
rect 19914 36038 19966 36090
rect 20018 36038 20070 36090
rect 20122 36038 29186 36090
rect 29238 36038 29290 36090
rect 29342 36038 29394 36090
rect 29446 36038 38510 36090
rect 38562 36038 38614 36090
rect 38666 36038 38718 36090
rect 38770 36038 38800 36090
rect 1344 36004 38800 36038
rect 3166 35922 3218 35934
rect 3166 35858 3218 35870
rect 4510 35922 4562 35934
rect 4510 35858 4562 35870
rect 5406 35922 5458 35934
rect 5406 35858 5458 35870
rect 5630 35922 5682 35934
rect 5630 35858 5682 35870
rect 6974 35922 7026 35934
rect 6974 35858 7026 35870
rect 9102 35922 9154 35934
rect 9102 35858 9154 35870
rect 9662 35922 9714 35934
rect 9662 35858 9714 35870
rect 15262 35922 15314 35934
rect 15262 35858 15314 35870
rect 15934 35922 15986 35934
rect 15934 35858 15986 35870
rect 16382 35922 16434 35934
rect 16382 35858 16434 35870
rect 27134 35922 27186 35934
rect 27134 35858 27186 35870
rect 33742 35922 33794 35934
rect 33742 35858 33794 35870
rect 34526 35922 34578 35934
rect 34526 35858 34578 35870
rect 37550 35810 37602 35822
rect 5954 35758 5966 35810
rect 6018 35758 6030 35810
rect 9986 35758 9998 35810
rect 10050 35758 10062 35810
rect 37550 35746 37602 35758
rect 38222 35810 38274 35822
rect 38222 35746 38274 35758
rect 37214 35698 37266 35710
rect 16594 35646 16606 35698
rect 16658 35646 16670 35698
rect 27346 35646 27358 35698
rect 27410 35646 27422 35698
rect 34738 35646 34750 35698
rect 34802 35646 34814 35698
rect 37214 35634 37266 35646
rect 37886 35698 37938 35710
rect 37886 35634 37938 35646
rect 3614 35586 3666 35598
rect 3614 35522 3666 35534
rect 4174 35586 4226 35598
rect 4174 35522 4226 35534
rect 6414 35586 6466 35598
rect 6414 35522 6466 35534
rect 10446 35586 10498 35598
rect 10446 35522 10498 35534
rect 32510 35586 32562 35598
rect 32510 35522 32562 35534
rect 33182 35586 33234 35598
rect 33182 35522 33234 35534
rect 34190 35586 34242 35598
rect 34190 35522 34242 35534
rect 35310 35586 35362 35598
rect 35310 35522 35362 35534
rect 35758 35586 35810 35598
rect 35758 35522 35810 35534
rect 36318 35586 36370 35598
rect 36318 35522 36370 35534
rect 36878 35586 36930 35598
rect 36878 35522 36930 35534
rect 4162 35422 4174 35474
rect 4226 35471 4238 35474
rect 4610 35471 4622 35474
rect 4226 35425 4622 35471
rect 4226 35422 4238 35425
rect 4610 35422 4622 35425
rect 4674 35422 4686 35474
rect 1344 35306 38640 35340
rect 1344 35254 5876 35306
rect 5928 35254 5980 35306
rect 6032 35254 6084 35306
rect 6136 35254 15200 35306
rect 15252 35254 15304 35306
rect 15356 35254 15408 35306
rect 15460 35254 24524 35306
rect 24576 35254 24628 35306
rect 24680 35254 24732 35306
rect 24784 35254 33848 35306
rect 33900 35254 33952 35306
rect 34004 35254 34056 35306
rect 34108 35254 38640 35306
rect 1344 35220 38640 35254
rect 37662 34802 37714 34814
rect 37662 34738 37714 34750
rect 37886 34802 37938 34814
rect 37886 34738 37938 34750
rect 37102 34690 37154 34702
rect 37102 34626 37154 34638
rect 38222 34690 38274 34702
rect 38222 34626 38274 34638
rect 1344 34522 38800 34556
rect 1344 34470 10538 34522
rect 10590 34470 10642 34522
rect 10694 34470 10746 34522
rect 10798 34470 19862 34522
rect 19914 34470 19966 34522
rect 20018 34470 20070 34522
rect 20122 34470 29186 34522
rect 29238 34470 29290 34522
rect 29342 34470 29394 34522
rect 29446 34470 38510 34522
rect 38562 34470 38614 34522
rect 38666 34470 38718 34522
rect 38770 34470 38800 34522
rect 1344 34436 38800 34470
rect 38222 34242 38274 34254
rect 38222 34178 38274 34190
rect 37986 34078 37998 34130
rect 38050 34078 38062 34130
rect 37550 34018 37602 34030
rect 37550 33954 37602 33966
rect 1344 33738 38640 33772
rect 1344 33686 5876 33738
rect 5928 33686 5980 33738
rect 6032 33686 6084 33738
rect 6136 33686 15200 33738
rect 15252 33686 15304 33738
rect 15356 33686 15408 33738
rect 15460 33686 24524 33738
rect 24576 33686 24628 33738
rect 24680 33686 24732 33738
rect 24784 33686 33848 33738
rect 33900 33686 33952 33738
rect 34004 33686 34056 33738
rect 34108 33686 38640 33738
rect 1344 33652 38640 33686
rect 37886 33234 37938 33246
rect 37886 33170 37938 33182
rect 1710 33122 1762 33134
rect 2494 33122 2546 33134
rect 2034 33070 2046 33122
rect 2098 33070 2110 33122
rect 1710 33058 1762 33070
rect 2494 33058 2546 33070
rect 37662 33122 37714 33134
rect 37662 33058 37714 33070
rect 38222 33122 38274 33134
rect 38222 33058 38274 33070
rect 1344 32954 38800 32988
rect 1344 32902 10538 32954
rect 10590 32902 10642 32954
rect 10694 32902 10746 32954
rect 10798 32902 19862 32954
rect 19914 32902 19966 32954
rect 20018 32902 20070 32954
rect 20122 32902 29186 32954
rect 29238 32902 29290 32954
rect 29342 32902 29394 32954
rect 29446 32902 38510 32954
rect 38562 32902 38614 32954
rect 38666 32902 38718 32954
rect 38770 32902 38800 32954
rect 1344 32868 38800 32902
rect 1710 32674 1762 32686
rect 1710 32610 1762 32622
rect 38222 32674 38274 32686
rect 38222 32610 38274 32622
rect 2046 32562 2098 32574
rect 2046 32498 2098 32510
rect 37550 32562 37602 32574
rect 37986 32510 37998 32562
rect 38050 32510 38062 32562
rect 37550 32498 37602 32510
rect 2606 32450 2658 32462
rect 2606 32386 2658 32398
rect 2942 32450 2994 32462
rect 2942 32386 2994 32398
rect 2258 32286 2270 32338
rect 2322 32335 2334 32338
rect 2930 32335 2942 32338
rect 2322 32289 2942 32335
rect 2322 32286 2334 32289
rect 2930 32286 2942 32289
rect 2994 32286 3006 32338
rect 1344 32170 38640 32204
rect 1344 32118 5876 32170
rect 5928 32118 5980 32170
rect 6032 32118 6084 32170
rect 6136 32118 15200 32170
rect 15252 32118 15304 32170
rect 15356 32118 15408 32170
rect 15460 32118 24524 32170
rect 24576 32118 24628 32170
rect 24680 32118 24732 32170
rect 24784 32118 33848 32170
rect 33900 32118 33952 32170
rect 34004 32118 34056 32170
rect 34108 32118 38640 32170
rect 1344 32084 38640 32118
rect 2046 31666 2098 31678
rect 2046 31602 2098 31614
rect 2382 31666 2434 31678
rect 2382 31602 2434 31614
rect 2718 31666 2770 31678
rect 2718 31602 2770 31614
rect 37214 31666 37266 31678
rect 37214 31602 37266 31614
rect 37550 31666 37602 31678
rect 37550 31602 37602 31614
rect 37886 31666 37938 31678
rect 37886 31602 37938 31614
rect 1710 31554 1762 31566
rect 1710 31490 1762 31502
rect 3278 31554 3330 31566
rect 3278 31490 3330 31502
rect 38222 31554 38274 31566
rect 38222 31490 38274 31502
rect 1344 31386 38800 31420
rect 1344 31334 10538 31386
rect 10590 31334 10642 31386
rect 10694 31334 10746 31386
rect 10798 31334 19862 31386
rect 19914 31334 19966 31386
rect 20018 31334 20070 31386
rect 20122 31334 29186 31386
rect 29238 31334 29290 31386
rect 29342 31334 29394 31386
rect 29446 31334 38510 31386
rect 38562 31334 38614 31386
rect 38666 31334 38718 31386
rect 38770 31334 38800 31386
rect 1344 31300 38800 31334
rect 1710 31106 1762 31118
rect 1710 31042 1762 31054
rect 38222 31106 38274 31118
rect 38222 31042 38274 31054
rect 37886 30994 37938 31006
rect 1922 30942 1934 30994
rect 1986 30942 1998 30994
rect 37886 30930 37938 30942
rect 2494 30882 2546 30894
rect 2494 30818 2546 30830
rect 1344 30602 38640 30636
rect 1344 30550 5876 30602
rect 5928 30550 5980 30602
rect 6032 30550 6084 30602
rect 6136 30550 15200 30602
rect 15252 30550 15304 30602
rect 15356 30550 15408 30602
rect 15460 30550 24524 30602
rect 24576 30550 24628 30602
rect 24680 30550 24732 30602
rect 24784 30550 33848 30602
rect 33900 30550 33952 30602
rect 34004 30550 34056 30602
rect 34108 30550 38640 30602
rect 1344 30516 38640 30550
rect 18946 30158 18958 30210
rect 19010 30158 19022 30210
rect 21522 30158 21534 30210
rect 21586 30158 21598 30210
rect 24098 30158 24110 30210
rect 24162 30158 24174 30210
rect 25554 30158 25566 30210
rect 25618 30158 25630 30210
rect 28018 30158 28030 30210
rect 28082 30158 28094 30210
rect 2046 30098 2098 30110
rect 2046 30034 2098 30046
rect 13694 30098 13746 30110
rect 13694 30034 13746 30046
rect 14030 30098 14082 30110
rect 14030 30034 14082 30046
rect 18734 30098 18786 30110
rect 18734 30034 18786 30046
rect 21758 30098 21810 30110
rect 21758 30034 21810 30046
rect 22094 30098 22146 30110
rect 22094 30034 22146 30046
rect 22430 30098 22482 30110
rect 22430 30034 22482 30046
rect 23326 30098 23378 30110
rect 23326 30034 23378 30046
rect 23662 30098 23714 30110
rect 23662 30034 23714 30046
rect 24334 30098 24386 30110
rect 24334 30034 24386 30046
rect 25790 30098 25842 30110
rect 25790 30034 25842 30046
rect 26126 30098 26178 30110
rect 26126 30034 26178 30046
rect 26462 30098 26514 30110
rect 26462 30034 26514 30046
rect 27246 30098 27298 30110
rect 27246 30034 27298 30046
rect 27582 30098 27634 30110
rect 27582 30034 27634 30046
rect 28254 30098 28306 30110
rect 28254 30034 28306 30046
rect 37886 30098 37938 30110
rect 37886 30034 37938 30046
rect 1710 29986 1762 29998
rect 1710 29922 1762 29934
rect 2606 29986 2658 29998
rect 2606 29922 2658 29934
rect 17390 29986 17442 29998
rect 17390 29922 17442 29934
rect 18398 29986 18450 29998
rect 18398 29922 18450 29934
rect 19630 29986 19682 29998
rect 19630 29922 19682 29934
rect 38222 29986 38274 29998
rect 38222 29922 38274 29934
rect 1344 29818 38800 29852
rect 1344 29766 10538 29818
rect 10590 29766 10642 29818
rect 10694 29766 10746 29818
rect 10798 29766 19862 29818
rect 19914 29766 19966 29818
rect 20018 29766 20070 29818
rect 20122 29766 29186 29818
rect 29238 29766 29290 29818
rect 29342 29766 29394 29818
rect 29446 29766 38510 29818
rect 38562 29766 38614 29818
rect 38666 29766 38718 29818
rect 38770 29766 38800 29818
rect 1344 29732 38800 29766
rect 14366 29650 14418 29662
rect 14366 29586 14418 29598
rect 18734 29650 18786 29662
rect 18734 29586 18786 29598
rect 19630 29650 19682 29662
rect 21522 29598 21534 29650
rect 21586 29598 21598 29650
rect 21858 29598 21870 29650
rect 21922 29598 21934 29650
rect 23314 29598 23326 29650
rect 23378 29598 23390 29650
rect 24210 29598 24222 29650
rect 24274 29598 24286 29650
rect 25778 29598 25790 29650
rect 25842 29598 25854 29650
rect 27122 29598 27134 29650
rect 27186 29598 27198 29650
rect 28018 29598 28030 29650
rect 28082 29598 28094 29650
rect 19630 29586 19682 29598
rect 1710 29538 1762 29550
rect 1710 29474 1762 29486
rect 14030 29538 14082 29550
rect 14030 29474 14082 29486
rect 19294 29538 19346 29550
rect 19294 29474 19346 29486
rect 19966 29538 20018 29550
rect 19966 29474 20018 29486
rect 20302 29538 20354 29550
rect 20302 29474 20354 29486
rect 38222 29538 38274 29550
rect 38222 29474 38274 29486
rect 2046 29426 2098 29438
rect 15822 29426 15874 29438
rect 13234 29374 13246 29426
rect 13298 29374 13310 29426
rect 14578 29374 14590 29426
rect 14642 29374 14654 29426
rect 2046 29362 2098 29374
rect 15822 29362 15874 29374
rect 16718 29426 16770 29438
rect 16718 29362 16770 29374
rect 17838 29426 17890 29438
rect 17838 29362 17890 29374
rect 17950 29426 18002 29438
rect 17950 29362 18002 29374
rect 18062 29426 18114 29438
rect 22430 29426 22482 29438
rect 18274 29374 18286 29426
rect 18338 29374 18350 29426
rect 18062 29362 18114 29374
rect 22430 29362 22482 29374
rect 37886 29426 37938 29438
rect 37886 29362 37938 29374
rect 2494 29314 2546 29326
rect 2494 29250 2546 29262
rect 15374 29314 15426 29326
rect 15374 29250 15426 29262
rect 16270 29314 16322 29326
rect 16270 29250 16322 29262
rect 20974 29314 21026 29326
rect 20974 29250 21026 29262
rect 22766 29314 22818 29326
rect 22766 29250 22818 29262
rect 23662 29314 23714 29326
rect 23662 29250 23714 29262
rect 25230 29314 25282 29326
rect 25230 29250 25282 29262
rect 26574 29314 26626 29326
rect 26574 29250 26626 29262
rect 27470 29314 27522 29326
rect 27470 29250 27522 29262
rect 13470 29202 13522 29214
rect 13470 29138 13522 29150
rect 13694 29202 13746 29214
rect 13694 29138 13746 29150
rect 13918 29202 13970 29214
rect 13918 29138 13970 29150
rect 16158 29202 16210 29214
rect 16158 29138 16210 29150
rect 16606 29202 16658 29214
rect 16606 29138 16658 29150
rect 21198 29202 21250 29214
rect 21198 29138 21250 29150
rect 22206 29202 22258 29214
rect 22206 29138 22258 29150
rect 22990 29202 23042 29214
rect 22990 29138 23042 29150
rect 23886 29202 23938 29214
rect 23886 29138 23938 29150
rect 25454 29202 25506 29214
rect 25454 29138 25506 29150
rect 26798 29202 26850 29214
rect 26798 29138 26850 29150
rect 27694 29202 27746 29214
rect 27694 29138 27746 29150
rect 1344 29034 38640 29068
rect 1344 28982 5876 29034
rect 5928 28982 5980 29034
rect 6032 28982 6084 29034
rect 6136 28982 15200 29034
rect 15252 28982 15304 29034
rect 15356 28982 15408 29034
rect 15460 28982 24524 29034
rect 24576 28982 24628 29034
rect 24680 28982 24732 29034
rect 24784 28982 33848 29034
rect 33900 28982 33952 29034
rect 34004 28982 34056 29034
rect 34108 28982 38640 29034
rect 1344 28948 38640 28982
rect 14254 28866 14306 28878
rect 14254 28802 14306 28814
rect 15486 28866 15538 28878
rect 15486 28802 15538 28814
rect 15822 28866 15874 28878
rect 15822 28802 15874 28814
rect 18734 28866 18786 28878
rect 18734 28802 18786 28814
rect 25230 28866 25282 28878
rect 25554 28814 25566 28866
rect 25618 28814 25630 28866
rect 25230 28802 25282 28814
rect 13918 28754 13970 28766
rect 13918 28690 13970 28702
rect 16494 28754 16546 28766
rect 16494 28690 16546 28702
rect 16942 28754 16994 28766
rect 16942 28690 16994 28702
rect 17390 28754 17442 28766
rect 17390 28690 17442 28702
rect 13582 28642 13634 28654
rect 13582 28578 13634 28590
rect 13694 28642 13746 28654
rect 13694 28578 13746 28590
rect 14142 28642 14194 28654
rect 14142 28578 14194 28590
rect 15598 28642 15650 28654
rect 17838 28642 17890 28654
rect 16034 28590 16046 28642
rect 16098 28590 16110 28642
rect 15598 28578 15650 28590
rect 17838 28578 17890 28590
rect 17950 28642 18002 28654
rect 17950 28578 18002 28590
rect 18062 28642 18114 28654
rect 19854 28642 19906 28654
rect 18386 28590 18398 28642
rect 18450 28590 18462 28642
rect 19170 28590 19182 28642
rect 19234 28590 19246 28642
rect 18062 28578 18114 28590
rect 19854 28578 19906 28590
rect 21758 28642 21810 28654
rect 21758 28578 21810 28590
rect 21870 28642 21922 28654
rect 21870 28578 21922 28590
rect 22430 28642 22482 28654
rect 22430 28578 22482 28590
rect 25006 28642 25058 28654
rect 26002 28590 26014 28642
rect 26066 28590 26078 28642
rect 25006 28578 25058 28590
rect 2046 28530 2098 28542
rect 2046 28466 2098 28478
rect 11454 28530 11506 28542
rect 11454 28466 11506 28478
rect 11790 28530 11842 28542
rect 23774 28530 23826 28542
rect 22082 28478 22094 28530
rect 22146 28478 22158 28530
rect 11790 28466 11842 28478
rect 23774 28466 23826 28478
rect 24110 28530 24162 28542
rect 24110 28466 24162 28478
rect 26238 28530 26290 28542
rect 26238 28466 26290 28478
rect 27358 28530 27410 28542
rect 27358 28466 27410 28478
rect 27694 28530 27746 28542
rect 27694 28466 27746 28478
rect 37886 28530 37938 28542
rect 37886 28466 37938 28478
rect 1710 28418 1762 28430
rect 1710 28354 1762 28366
rect 18958 28418 19010 28430
rect 18958 28354 19010 28366
rect 22654 28418 22706 28430
rect 22654 28354 22706 28366
rect 38222 28418 38274 28430
rect 38222 28354 38274 28366
rect 1344 28250 38800 28284
rect 1344 28198 10538 28250
rect 10590 28198 10642 28250
rect 10694 28198 10746 28250
rect 10798 28198 19862 28250
rect 19914 28198 19966 28250
rect 20018 28198 20070 28250
rect 20122 28198 29186 28250
rect 29238 28198 29290 28250
rect 29342 28198 29394 28250
rect 29446 28198 38510 28250
rect 38562 28198 38614 28250
rect 38666 28198 38718 28250
rect 38770 28198 38800 28250
rect 1344 28164 38800 28198
rect 12350 28082 12402 28094
rect 12350 28018 12402 28030
rect 19854 28082 19906 28094
rect 19854 28018 19906 28030
rect 23550 28082 23602 28094
rect 23550 28018 23602 28030
rect 24222 28082 24274 28094
rect 28926 28082 28978 28094
rect 26002 28030 26014 28082
rect 26066 28030 26078 28082
rect 24222 28018 24274 28030
rect 28926 28018 28978 28030
rect 1710 27970 1762 27982
rect 1710 27906 1762 27918
rect 14702 27970 14754 27982
rect 14702 27906 14754 27918
rect 15598 27970 15650 27982
rect 15598 27906 15650 27918
rect 18398 27970 18450 27982
rect 18398 27906 18450 27918
rect 20190 27970 20242 27982
rect 20190 27906 20242 27918
rect 20526 27970 20578 27982
rect 20526 27906 20578 27918
rect 22094 27970 22146 27982
rect 22094 27906 22146 27918
rect 22206 27970 22258 27982
rect 22206 27906 22258 27918
rect 25454 27970 25506 27982
rect 25454 27906 25506 27918
rect 26574 27970 26626 27982
rect 26574 27906 26626 27918
rect 27694 27970 27746 27982
rect 27694 27906 27746 27918
rect 38222 27970 38274 27982
rect 38222 27906 38274 27918
rect 2046 27858 2098 27870
rect 14814 27858 14866 27870
rect 15710 27858 15762 27870
rect 12562 27806 12574 27858
rect 12626 27806 12638 27858
rect 13122 27806 13134 27858
rect 13186 27806 13198 27858
rect 15250 27806 15262 27858
rect 15314 27806 15326 27858
rect 2046 27794 2098 27806
rect 14814 27794 14866 27806
rect 15710 27794 15762 27806
rect 16046 27858 16098 27870
rect 16046 27794 16098 27806
rect 18286 27858 18338 27870
rect 19070 27858 19122 27870
rect 18610 27806 18622 27858
rect 18674 27806 18686 27858
rect 18286 27794 18338 27806
rect 19070 27794 19122 27806
rect 19518 27858 19570 27870
rect 19518 27794 19570 27806
rect 21870 27858 21922 27870
rect 22878 27858 22930 27870
rect 22418 27806 22430 27858
rect 22482 27806 22494 27858
rect 21870 27794 21922 27806
rect 22878 27794 22930 27806
rect 23214 27858 23266 27870
rect 23214 27794 23266 27806
rect 23886 27858 23938 27870
rect 23886 27794 23938 27806
rect 25342 27858 25394 27870
rect 25342 27794 25394 27806
rect 25566 27858 25618 27870
rect 25566 27794 25618 27806
rect 26462 27858 26514 27870
rect 26462 27794 26514 27806
rect 26686 27858 26738 27870
rect 27806 27858 27858 27870
rect 28590 27858 28642 27870
rect 27458 27806 27470 27858
rect 27522 27806 27534 27858
rect 28242 27806 28254 27858
rect 28306 27806 28318 27858
rect 37986 27806 37998 27858
rect 38050 27806 38062 27858
rect 26686 27794 26738 27806
rect 27806 27794 27858 27806
rect 28590 27794 28642 27806
rect 12014 27746 12066 27758
rect 12014 27682 12066 27694
rect 16942 27746 16994 27758
rect 16942 27682 16994 27694
rect 17502 27746 17554 27758
rect 17502 27682 17554 27694
rect 18062 27746 18114 27758
rect 18062 27682 18114 27694
rect 37550 27746 37602 27758
rect 37550 27682 37602 27694
rect 11342 27634 11394 27646
rect 11342 27570 11394 27582
rect 11454 27634 11506 27646
rect 11454 27570 11506 27582
rect 11678 27634 11730 27646
rect 11678 27570 11730 27582
rect 11902 27634 11954 27646
rect 11902 27570 11954 27582
rect 13358 27634 13410 27646
rect 13358 27570 13410 27582
rect 13582 27634 13634 27646
rect 13582 27570 13634 27582
rect 13806 27634 13858 27646
rect 13806 27570 13858 27582
rect 13918 27634 13970 27646
rect 13918 27570 13970 27582
rect 15038 27634 15090 27646
rect 15038 27570 15090 27582
rect 15934 27634 15986 27646
rect 15934 27570 15986 27582
rect 17390 27634 17442 27646
rect 27122 27582 27134 27634
rect 27186 27582 27198 27634
rect 17390 27570 17442 27582
rect 1344 27466 38640 27500
rect 1344 27414 5876 27466
rect 5928 27414 5980 27466
rect 6032 27414 6084 27466
rect 6136 27414 15200 27466
rect 15252 27414 15304 27466
rect 15356 27414 15408 27466
rect 15460 27414 24524 27466
rect 24576 27414 24628 27466
rect 24680 27414 24732 27466
rect 24784 27414 33848 27466
rect 33900 27414 33952 27466
rect 34004 27414 34056 27466
rect 34108 27414 38640 27466
rect 1344 27380 38640 27414
rect 10446 27298 10498 27310
rect 10446 27234 10498 27246
rect 10670 27298 10722 27310
rect 10670 27234 10722 27246
rect 20190 27186 20242 27198
rect 15922 27134 15934 27186
rect 15986 27134 15998 27186
rect 20190 27122 20242 27134
rect 21758 27186 21810 27198
rect 21758 27122 21810 27134
rect 10222 27074 10274 27086
rect 12350 27074 12402 27086
rect 10882 27022 10894 27074
rect 10946 27022 10958 27074
rect 11218 27022 11230 27074
rect 11282 27022 11294 27074
rect 10222 27010 10274 27022
rect 12350 27010 12402 27022
rect 13918 27074 13970 27086
rect 15374 27074 15426 27086
rect 14914 27022 14926 27074
rect 14978 27022 14990 27074
rect 13918 27010 13970 27022
rect 15374 27010 15426 27022
rect 15710 27074 15762 27086
rect 17950 27074 18002 27086
rect 16146 27022 16158 27074
rect 16210 27022 16222 27074
rect 17378 27022 17390 27074
rect 17442 27022 17454 27074
rect 15710 27010 15762 27022
rect 17950 27010 18002 27022
rect 18174 27074 18226 27086
rect 21982 27074 22034 27086
rect 22990 27074 23042 27086
rect 24894 27074 24946 27086
rect 18498 27022 18510 27074
rect 18562 27022 18574 27074
rect 22306 27022 22318 27074
rect 22370 27022 22382 27074
rect 24658 27022 24670 27074
rect 24722 27022 24734 27074
rect 18174 27010 18226 27022
rect 21982 27010 22034 27022
rect 22990 27010 23042 27022
rect 24894 27010 24946 27022
rect 25006 27074 25058 27086
rect 37214 27074 37266 27086
rect 26898 27022 26910 27074
rect 26962 27022 26974 27074
rect 25006 27010 25058 27022
rect 37214 27010 37266 27022
rect 2046 26962 2098 26974
rect 2046 26898 2098 26910
rect 2382 26962 2434 26974
rect 2382 26898 2434 26910
rect 2718 26962 2770 26974
rect 2718 26898 2770 26910
rect 9438 26962 9490 26974
rect 9438 26898 9490 26910
rect 9774 26962 9826 26974
rect 9774 26898 9826 26910
rect 10110 26962 10162 26974
rect 13582 26962 13634 26974
rect 17614 26962 17666 26974
rect 18958 26962 19010 26974
rect 11330 26910 11342 26962
rect 11394 26910 11406 26962
rect 12786 26910 12798 26962
rect 12850 26910 12862 26962
rect 15138 26910 15150 26962
rect 15202 26910 15214 26962
rect 18386 26910 18398 26962
rect 18450 26910 18462 26962
rect 10110 26898 10162 26910
rect 13582 26898 13634 26910
rect 17614 26898 17666 26910
rect 18958 26898 19010 26910
rect 19406 26962 19458 26974
rect 19406 26898 19458 26910
rect 19742 26962 19794 26974
rect 22766 26962 22818 26974
rect 22194 26910 22206 26962
rect 22258 26910 22270 26962
rect 19742 26898 19794 26910
rect 22766 26898 22818 26910
rect 23326 26962 23378 26974
rect 25790 26962 25842 26974
rect 25442 26910 25454 26962
rect 25506 26910 25518 26962
rect 23326 26898 23378 26910
rect 25790 26898 25842 26910
rect 26126 26962 26178 26974
rect 26126 26898 26178 26910
rect 27134 26962 27186 26974
rect 27134 26898 27186 26910
rect 28254 26962 28306 26974
rect 28254 26898 28306 26910
rect 28590 26962 28642 26974
rect 28590 26898 28642 26910
rect 37550 26962 37602 26974
rect 37550 26898 37602 26910
rect 37886 26962 37938 26974
rect 37886 26898 37938 26910
rect 38222 26962 38274 26974
rect 38222 26898 38274 26910
rect 1710 26850 1762 26862
rect 11890 26798 11902 26850
rect 11954 26798 11966 26850
rect 1710 26786 1762 26798
rect 1344 26682 38800 26716
rect 1344 26630 10538 26682
rect 10590 26630 10642 26682
rect 10694 26630 10746 26682
rect 10798 26630 19862 26682
rect 19914 26630 19966 26682
rect 20018 26630 20070 26682
rect 20122 26630 29186 26682
rect 29238 26630 29290 26682
rect 29342 26630 29394 26682
rect 29446 26630 38510 26682
rect 38562 26630 38614 26682
rect 38666 26630 38718 26682
rect 38770 26630 38800 26682
rect 1344 26596 38800 26630
rect 10110 26514 10162 26526
rect 10110 26450 10162 26462
rect 11678 26514 11730 26526
rect 11678 26450 11730 26462
rect 13022 26514 13074 26526
rect 13022 26450 13074 26462
rect 14478 26514 14530 26526
rect 16606 26514 16658 26526
rect 15922 26462 15934 26514
rect 15986 26462 15998 26514
rect 14478 26450 14530 26462
rect 16606 26450 16658 26462
rect 17838 26514 17890 26526
rect 17838 26450 17890 26462
rect 18174 26514 18226 26526
rect 18174 26450 18226 26462
rect 21534 26514 21586 26526
rect 21534 26450 21586 26462
rect 23438 26514 23490 26526
rect 23438 26450 23490 26462
rect 26462 26514 26514 26526
rect 28130 26462 28142 26514
rect 28194 26462 28206 26514
rect 26462 26450 26514 26462
rect 1710 26402 1762 26414
rect 1710 26338 1762 26350
rect 10446 26402 10498 26414
rect 10446 26338 10498 26350
rect 15598 26402 15650 26414
rect 15598 26338 15650 26350
rect 17502 26402 17554 26414
rect 17502 26338 17554 26350
rect 19182 26402 19234 26414
rect 24110 26402 24162 26414
rect 21970 26350 21982 26402
rect 22034 26350 22046 26402
rect 19182 26338 19234 26350
rect 24110 26338 24162 26350
rect 38222 26402 38274 26414
rect 38222 26338 38274 26350
rect 2046 26290 2098 26302
rect 2046 26226 2098 26238
rect 9774 26290 9826 26302
rect 11342 26290 11394 26302
rect 10658 26238 10670 26290
rect 10722 26238 10734 26290
rect 11106 26238 11118 26290
rect 11170 26238 11182 26290
rect 9774 26226 9826 26238
rect 11342 26226 11394 26238
rect 12686 26290 12738 26302
rect 12686 26226 12738 26238
rect 13582 26290 13634 26302
rect 13582 26226 13634 26238
rect 14142 26290 14194 26302
rect 16270 26290 16322 26302
rect 18846 26290 18898 26302
rect 14690 26238 14702 26290
rect 14754 26238 14766 26290
rect 18386 26238 18398 26290
rect 18450 26238 18462 26290
rect 14142 26226 14194 26238
rect 16270 26226 16322 26238
rect 18846 26226 18898 26238
rect 19742 26290 19794 26302
rect 19742 26226 19794 26238
rect 19854 26290 19906 26302
rect 21870 26290 21922 26302
rect 20066 26238 20078 26290
rect 20130 26238 20142 26290
rect 21298 26238 21310 26290
rect 21362 26238 21374 26290
rect 19854 26226 19906 26238
rect 21870 26226 21922 26238
rect 22206 26290 22258 26302
rect 22878 26290 22930 26302
rect 22418 26238 22430 26290
rect 22482 26238 22494 26290
rect 22206 26226 22258 26238
rect 22878 26226 22930 26238
rect 23102 26290 23154 26302
rect 23102 26226 23154 26238
rect 23774 26290 23826 26302
rect 23774 26226 23826 26238
rect 26798 26290 26850 26302
rect 26798 26226 26850 26238
rect 27806 26290 27858 26302
rect 27806 26226 27858 26238
rect 37886 26290 37938 26302
rect 37886 26226 37938 26238
rect 11566 26178 11618 26190
rect 11566 26114 11618 26126
rect 13806 26178 13858 26190
rect 13806 26114 13858 26126
rect 16718 26178 16770 26190
rect 16718 26114 16770 26126
rect 19518 26178 19570 26190
rect 19518 26114 19570 26126
rect 27582 26178 27634 26190
rect 27582 26114 27634 26126
rect 11790 26066 11842 26078
rect 11790 26002 11842 26014
rect 13470 26066 13522 26078
rect 13470 26002 13522 26014
rect 14030 26066 14082 26078
rect 14030 26002 14082 26014
rect 20526 26066 20578 26078
rect 20526 26002 20578 26014
rect 1344 25898 38640 25932
rect 1344 25846 5876 25898
rect 5928 25846 5980 25898
rect 6032 25846 6084 25898
rect 6136 25846 15200 25898
rect 15252 25846 15304 25898
rect 15356 25846 15408 25898
rect 15460 25846 24524 25898
rect 24576 25846 24628 25898
rect 24680 25846 24732 25898
rect 24784 25846 33848 25898
rect 33900 25846 33952 25898
rect 34004 25846 34056 25898
rect 34108 25846 38640 25898
rect 1344 25812 38640 25846
rect 15262 25730 15314 25742
rect 15262 25666 15314 25678
rect 18398 25730 18450 25742
rect 18398 25666 18450 25678
rect 18958 25730 19010 25742
rect 18958 25666 19010 25678
rect 22766 25730 22818 25742
rect 22766 25666 22818 25678
rect 23326 25730 23378 25742
rect 23326 25666 23378 25678
rect 24670 25730 24722 25742
rect 24670 25666 24722 25678
rect 14926 25618 14978 25630
rect 14926 25554 14978 25566
rect 16158 25618 16210 25630
rect 16158 25554 16210 25566
rect 18846 25618 18898 25630
rect 18846 25554 18898 25566
rect 15150 25506 15202 25518
rect 17390 25506 17442 25518
rect 22878 25506 22930 25518
rect 11666 25454 11678 25506
rect 11730 25454 11742 25506
rect 16818 25454 16830 25506
rect 16882 25454 16894 25506
rect 17938 25454 17950 25506
rect 18002 25454 18014 25506
rect 20514 25454 20526 25506
rect 20578 25454 20590 25506
rect 15150 25442 15202 25454
rect 17390 25442 17442 25454
rect 22878 25442 22930 25454
rect 23102 25506 23154 25518
rect 23102 25442 23154 25454
rect 24446 25506 24498 25518
rect 26798 25506 26850 25518
rect 26562 25454 26574 25506
rect 26626 25454 26638 25506
rect 24446 25442 24498 25454
rect 26798 25442 26850 25454
rect 26910 25506 26962 25518
rect 26910 25442 26962 25454
rect 2046 25394 2098 25406
rect 2046 25330 2098 25342
rect 12462 25394 12514 25406
rect 12462 25330 12514 25342
rect 12798 25394 12850 25406
rect 12798 25330 12850 25342
rect 16382 25394 16434 25406
rect 16382 25330 16434 25342
rect 16494 25394 16546 25406
rect 16494 25330 16546 25342
rect 17614 25394 17666 25406
rect 17614 25330 17666 25342
rect 17726 25394 17778 25406
rect 17726 25330 17778 25342
rect 20750 25394 20802 25406
rect 20750 25330 20802 25342
rect 21310 25394 21362 25406
rect 21310 25330 21362 25342
rect 21646 25394 21698 25406
rect 21646 25330 21698 25342
rect 23438 25394 23490 25406
rect 23438 25330 23490 25342
rect 23774 25394 23826 25406
rect 23774 25330 23826 25342
rect 24110 25394 24162 25406
rect 25342 25394 25394 25406
rect 24994 25342 25006 25394
rect 25058 25342 25070 25394
rect 24110 25330 24162 25342
rect 25342 25330 25394 25342
rect 25678 25394 25730 25406
rect 27694 25394 27746 25406
rect 27346 25342 27358 25394
rect 27410 25342 27422 25394
rect 25678 25330 25730 25342
rect 27694 25330 27746 25342
rect 28030 25394 28082 25406
rect 28030 25330 28082 25342
rect 37886 25394 37938 25406
rect 37886 25330 37938 25342
rect 1710 25282 1762 25294
rect 1710 25218 1762 25230
rect 11454 25282 11506 25294
rect 11454 25218 11506 25230
rect 15262 25282 15314 25294
rect 15262 25218 15314 25230
rect 15822 25282 15874 25294
rect 15822 25218 15874 25230
rect 17166 25282 17218 25294
rect 17166 25218 17218 25230
rect 19406 25282 19458 25294
rect 19406 25218 19458 25230
rect 20078 25282 20130 25294
rect 20078 25218 20130 25230
rect 38222 25282 38274 25294
rect 38222 25218 38274 25230
rect 1344 25114 38800 25148
rect 1344 25062 10538 25114
rect 10590 25062 10642 25114
rect 10694 25062 10746 25114
rect 10798 25062 19862 25114
rect 19914 25062 19966 25114
rect 20018 25062 20070 25114
rect 20122 25062 29186 25114
rect 29238 25062 29290 25114
rect 29342 25062 29394 25114
rect 29446 25062 38510 25114
rect 38562 25062 38614 25114
rect 38666 25062 38718 25114
rect 38770 25062 38800 25114
rect 1344 25028 38800 25062
rect 13022 24946 13074 24958
rect 13022 24882 13074 24894
rect 14814 24946 14866 24958
rect 14814 24882 14866 24894
rect 17390 24946 17442 24958
rect 17390 24882 17442 24894
rect 22430 24946 22482 24958
rect 22430 24882 22482 24894
rect 29374 24946 29426 24958
rect 29374 24882 29426 24894
rect 1710 24834 1762 24846
rect 1710 24770 1762 24782
rect 2046 24834 2098 24846
rect 2046 24770 2098 24782
rect 9886 24834 9938 24846
rect 9886 24770 9938 24782
rect 10222 24834 10274 24846
rect 12014 24834 12066 24846
rect 11666 24782 11678 24834
rect 11730 24782 11742 24834
rect 10222 24770 10274 24782
rect 12014 24770 12066 24782
rect 12350 24834 12402 24846
rect 12350 24770 12402 24782
rect 20526 24834 20578 24846
rect 21198 24834 21250 24846
rect 20962 24782 20974 24834
rect 21026 24782 21038 24834
rect 20526 24770 20578 24782
rect 21198 24770 21250 24782
rect 24670 24834 24722 24846
rect 24670 24770 24722 24782
rect 26686 24834 26738 24846
rect 26686 24770 26738 24782
rect 27806 24834 27858 24846
rect 27806 24770 27858 24782
rect 38222 24834 38274 24846
rect 38222 24770 38274 24782
rect 10558 24722 10610 24734
rect 13358 24722 13410 24734
rect 9650 24670 9662 24722
rect 9714 24670 9726 24722
rect 11442 24670 11454 24722
rect 11506 24670 11518 24722
rect 10558 24658 10610 24670
rect 13358 24658 13410 24670
rect 13694 24722 13746 24734
rect 13694 24658 13746 24670
rect 13806 24722 13858 24734
rect 13806 24658 13858 24670
rect 14254 24722 14306 24734
rect 14254 24658 14306 24670
rect 15150 24722 15202 24734
rect 15150 24658 15202 24670
rect 15486 24722 15538 24734
rect 15486 24658 15538 24670
rect 16046 24722 16098 24734
rect 18958 24722 19010 24734
rect 17602 24670 17614 24722
rect 17666 24670 17678 24722
rect 16046 24658 16098 24670
rect 18958 24658 19010 24670
rect 20190 24722 20242 24734
rect 21870 24722 21922 24734
rect 21410 24670 21422 24722
rect 21474 24670 21486 24722
rect 20190 24658 20242 24670
rect 21870 24658 21922 24670
rect 22094 24722 22146 24734
rect 26574 24722 26626 24734
rect 27470 24722 27522 24734
rect 24434 24670 24446 24722
rect 24498 24670 24510 24722
rect 25218 24670 25230 24722
rect 25282 24670 25294 24722
rect 26338 24670 26350 24722
rect 26402 24670 26414 24722
rect 27122 24670 27134 24722
rect 27186 24670 27198 24722
rect 22094 24658 22146 24670
rect 26574 24658 26626 24670
rect 27470 24658 27522 24670
rect 28366 24722 28418 24734
rect 29038 24722 29090 24734
rect 28690 24670 28702 24722
rect 28754 24670 28766 24722
rect 28366 24658 28418 24670
rect 29038 24658 29090 24670
rect 37886 24722 37938 24734
rect 37886 24658 37938 24670
rect 16830 24610 16882 24622
rect 16830 24546 16882 24558
rect 18398 24610 18450 24622
rect 18398 24546 18450 24558
rect 19406 24610 19458 24622
rect 19406 24546 19458 24558
rect 20862 24610 20914 24622
rect 20862 24546 20914 24558
rect 25790 24610 25842 24622
rect 25790 24546 25842 24558
rect 28142 24610 28194 24622
rect 28142 24546 28194 24558
rect 14030 24498 14082 24510
rect 14030 24434 14082 24446
rect 14366 24498 14418 24510
rect 14366 24434 14418 24446
rect 15598 24498 15650 24510
rect 15598 24434 15650 24446
rect 15822 24498 15874 24510
rect 15822 24434 15874 24446
rect 16158 24498 16210 24510
rect 16158 24434 16210 24446
rect 18286 24498 18338 24510
rect 18286 24434 18338 24446
rect 18846 24498 18898 24510
rect 18846 24434 18898 24446
rect 19182 24498 19234 24510
rect 19182 24434 19234 24446
rect 19518 24498 19570 24510
rect 19518 24434 19570 24446
rect 25566 24498 25618 24510
rect 25566 24434 25618 24446
rect 1344 24330 38640 24364
rect 1344 24278 5876 24330
rect 5928 24278 5980 24330
rect 6032 24278 6084 24330
rect 6136 24278 15200 24330
rect 15252 24278 15304 24330
rect 15356 24278 15408 24330
rect 15460 24278 24524 24330
rect 24576 24278 24628 24330
rect 24680 24278 24732 24330
rect 24784 24278 33848 24330
rect 33900 24278 33952 24330
rect 34004 24278 34056 24330
rect 34108 24278 38640 24330
rect 1344 24244 38640 24278
rect 10222 24162 10274 24174
rect 10222 24098 10274 24110
rect 10670 24162 10722 24174
rect 10670 24098 10722 24110
rect 14478 24162 14530 24174
rect 14478 24098 14530 24110
rect 14702 24162 14754 24174
rect 14702 24098 14754 24110
rect 14814 24162 14866 24174
rect 14814 24098 14866 24110
rect 24446 24162 24498 24174
rect 24446 24098 24498 24110
rect 28142 24162 28194 24174
rect 28142 24098 28194 24110
rect 12350 24050 12402 24062
rect 12350 23986 12402 23998
rect 10446 23938 10498 23950
rect 12574 23938 12626 23950
rect 9426 23886 9438 23938
rect 9490 23886 9502 23938
rect 9986 23886 9998 23938
rect 10050 23886 10062 23938
rect 11554 23886 11566 23938
rect 11618 23886 11630 23938
rect 12114 23886 12126 23938
rect 12178 23886 12190 23938
rect 10446 23874 10498 23886
rect 12574 23874 12626 23886
rect 12798 23938 12850 23950
rect 12798 23874 12850 23886
rect 16606 23938 16658 23950
rect 16606 23874 16658 23886
rect 17278 23938 17330 23950
rect 18286 23938 18338 23950
rect 19518 23938 19570 23950
rect 24222 23938 24274 23950
rect 26574 23938 26626 23950
rect 17826 23886 17838 23938
rect 17890 23886 17902 23938
rect 18722 23886 18734 23938
rect 18786 23886 18798 23938
rect 23538 23886 23550 23938
rect 23602 23886 23614 23938
rect 26338 23886 26350 23938
rect 26402 23886 26414 23938
rect 17278 23874 17330 23886
rect 18286 23874 18338 23886
rect 19518 23874 19570 23886
rect 24222 23874 24274 23886
rect 26574 23874 26626 23886
rect 26686 23938 26738 23950
rect 26686 23874 26738 23886
rect 27918 23938 27970 23950
rect 27918 23874 27970 23886
rect 2046 23826 2098 23838
rect 2046 23762 2098 23774
rect 9662 23826 9714 23838
rect 9662 23762 9714 23774
rect 11790 23826 11842 23838
rect 11790 23762 11842 23774
rect 14366 23826 14418 23838
rect 14366 23762 14418 23774
rect 15374 23826 15426 23838
rect 15374 23762 15426 23774
rect 16270 23826 16322 23838
rect 19182 23826 19234 23838
rect 17378 23774 17390 23826
rect 17442 23774 17454 23826
rect 17714 23774 17726 23826
rect 17778 23774 17790 23826
rect 16270 23762 16322 23774
rect 19182 23762 19234 23774
rect 21310 23826 21362 23838
rect 21310 23762 21362 23774
rect 21646 23826 21698 23838
rect 21646 23762 21698 23774
rect 21982 23826 22034 23838
rect 21982 23762 22034 23774
rect 22318 23826 22370 23838
rect 22318 23762 22370 23774
rect 22990 23826 23042 23838
rect 22990 23762 23042 23774
rect 23326 23826 23378 23838
rect 25118 23826 25170 23838
rect 24770 23774 24782 23826
rect 24834 23774 24846 23826
rect 23326 23762 23378 23774
rect 25118 23762 25170 23774
rect 25454 23826 25506 23838
rect 29150 23826 29202 23838
rect 28466 23774 28478 23826
rect 28530 23774 28542 23826
rect 25454 23762 25506 23774
rect 29150 23762 29202 23774
rect 29486 23826 29538 23838
rect 29486 23762 29538 23774
rect 37886 23826 37938 23838
rect 37886 23762 37938 23774
rect 1710 23714 1762 23726
rect 1710 23650 1762 23662
rect 10558 23714 10610 23726
rect 10558 23650 10610 23662
rect 12686 23714 12738 23726
rect 12686 23650 12738 23662
rect 18510 23714 18562 23726
rect 18510 23650 18562 23662
rect 22654 23714 22706 23726
rect 38222 23714 38274 23726
rect 27122 23662 27134 23714
rect 27186 23662 27198 23714
rect 22654 23650 22706 23662
rect 38222 23650 38274 23662
rect 1344 23546 38800 23580
rect 1344 23494 10538 23546
rect 10590 23494 10642 23546
rect 10694 23494 10746 23546
rect 10798 23494 19862 23546
rect 19914 23494 19966 23546
rect 20018 23494 20070 23546
rect 20122 23494 29186 23546
rect 29238 23494 29290 23546
rect 29342 23494 29394 23546
rect 29446 23494 38510 23546
rect 38562 23494 38614 23546
rect 38666 23494 38718 23546
rect 38770 23494 38800 23546
rect 1344 23460 38800 23494
rect 10110 23378 10162 23390
rect 10110 23314 10162 23326
rect 14030 23378 14082 23390
rect 14030 23314 14082 23326
rect 16494 23378 16546 23390
rect 16494 23314 16546 23326
rect 17726 23378 17778 23390
rect 17726 23314 17778 23326
rect 24110 23378 24162 23390
rect 24110 23314 24162 23326
rect 26462 23378 26514 23390
rect 26462 23314 26514 23326
rect 27582 23378 27634 23390
rect 27582 23314 27634 23326
rect 27918 23378 27970 23390
rect 27918 23314 27970 23326
rect 31278 23378 31330 23390
rect 31278 23314 31330 23326
rect 32398 23378 32450 23390
rect 32398 23314 32450 23326
rect 1710 23266 1762 23278
rect 1710 23202 1762 23214
rect 12238 23266 12290 23278
rect 12238 23202 12290 23214
rect 12574 23266 12626 23278
rect 12574 23202 12626 23214
rect 18174 23266 18226 23278
rect 18174 23202 18226 23214
rect 19966 23266 20018 23278
rect 19966 23202 20018 23214
rect 20302 23266 20354 23278
rect 20302 23202 20354 23214
rect 20638 23266 20690 23278
rect 20638 23202 20690 23214
rect 23774 23266 23826 23278
rect 23774 23202 23826 23214
rect 27246 23266 27298 23278
rect 27246 23202 27298 23214
rect 29374 23266 29426 23278
rect 29374 23202 29426 23214
rect 30606 23266 30658 23278
rect 30606 23202 30658 23214
rect 38222 23266 38274 23278
rect 38222 23202 38274 23214
rect 2046 23154 2098 23166
rect 2046 23090 2098 23102
rect 10446 23154 10498 23166
rect 10446 23090 10498 23102
rect 13694 23154 13746 23166
rect 13694 23090 13746 23102
rect 13918 23154 13970 23166
rect 17390 23154 17442 23166
rect 14130 23102 14142 23154
rect 14194 23102 14206 23154
rect 14802 23102 14814 23154
rect 14866 23102 14878 23154
rect 15026 23102 15038 23154
rect 15090 23102 15102 23154
rect 16706 23102 16718 23154
rect 16770 23102 16782 23154
rect 13918 23090 13970 23102
rect 17390 23090 17442 23102
rect 18846 23154 18898 23166
rect 18846 23090 18898 23102
rect 19406 23154 19458 23166
rect 19406 23090 19458 23102
rect 23438 23154 23490 23166
rect 23438 23090 23490 23102
rect 24446 23154 24498 23166
rect 24446 23090 24498 23102
rect 26126 23154 26178 23166
rect 26126 23090 26178 23102
rect 28254 23154 28306 23166
rect 28254 23090 28306 23102
rect 29038 23154 29090 23166
rect 29038 23090 29090 23102
rect 30270 23154 30322 23166
rect 32062 23154 32114 23166
rect 31042 23102 31054 23154
rect 31106 23102 31118 23154
rect 30270 23090 30322 23102
rect 32062 23090 32114 23102
rect 37886 23154 37938 23166
rect 37886 23090 37938 23102
rect 19182 23042 19234 23054
rect 14690 22990 14702 23042
rect 14754 22990 14766 23042
rect 19182 22978 19234 22990
rect 21310 23042 21362 23054
rect 21310 22978 21362 22990
rect 13470 22930 13522 22942
rect 18062 22930 18114 22942
rect 14578 22878 14590 22930
rect 14642 22878 14654 22930
rect 13470 22866 13522 22878
rect 18062 22866 18114 22878
rect 18958 22930 19010 22942
rect 18958 22866 19010 22878
rect 19518 22930 19570 22942
rect 19518 22866 19570 22878
rect 1344 22762 38640 22796
rect 1344 22710 5876 22762
rect 5928 22710 5980 22762
rect 6032 22710 6084 22762
rect 6136 22710 15200 22762
rect 15252 22710 15304 22762
rect 15356 22710 15408 22762
rect 15460 22710 24524 22762
rect 24576 22710 24628 22762
rect 24680 22710 24732 22762
rect 24784 22710 33848 22762
rect 33900 22710 33952 22762
rect 34004 22710 34056 22762
rect 34108 22710 38640 22762
rect 1344 22676 38640 22710
rect 9998 22594 10050 22606
rect 9998 22530 10050 22542
rect 10110 22594 10162 22606
rect 10110 22530 10162 22542
rect 10558 22594 10610 22606
rect 10558 22530 10610 22542
rect 12014 22594 12066 22606
rect 18622 22594 18674 22606
rect 17826 22542 17838 22594
rect 17890 22591 17902 22594
rect 18162 22591 18174 22594
rect 17890 22545 18174 22591
rect 17890 22542 17902 22545
rect 18162 22542 18174 22545
rect 18226 22542 18238 22594
rect 12014 22530 12066 22542
rect 18622 22530 18674 22542
rect 23326 22594 23378 22606
rect 30718 22594 30770 22606
rect 32510 22594 32562 22606
rect 30146 22542 30158 22594
rect 30210 22542 30222 22594
rect 31042 22542 31054 22594
rect 31106 22542 31118 22594
rect 31938 22542 31950 22594
rect 32002 22542 32014 22594
rect 23326 22530 23378 22542
rect 30718 22530 30770 22542
rect 32510 22530 32562 22542
rect 17838 22482 17890 22494
rect 17838 22418 17890 22430
rect 18286 22482 18338 22494
rect 18286 22418 18338 22430
rect 29598 22482 29650 22494
rect 29598 22418 29650 22430
rect 30494 22482 30546 22494
rect 30494 22418 30546 22430
rect 2718 22370 2770 22382
rect 2718 22306 2770 22318
rect 10334 22370 10386 22382
rect 10334 22306 10386 22318
rect 12126 22370 12178 22382
rect 12126 22306 12178 22318
rect 12350 22370 12402 22382
rect 12350 22306 12402 22318
rect 12574 22370 12626 22382
rect 16606 22370 16658 22382
rect 22430 22370 22482 22382
rect 14354 22318 14366 22370
rect 14418 22318 14430 22370
rect 15026 22318 15038 22370
rect 15090 22318 15102 22370
rect 19394 22318 19406 22370
rect 19458 22318 19470 22370
rect 21634 22318 21646 22370
rect 21698 22318 21710 22370
rect 12574 22306 12626 22318
rect 16606 22306 16658 22318
rect 22430 22306 22482 22318
rect 22654 22370 22706 22382
rect 23886 22370 23938 22382
rect 29822 22370 29874 22382
rect 22866 22318 22878 22370
rect 22930 22318 22942 22370
rect 25666 22318 25678 22370
rect 25730 22318 25742 22370
rect 22654 22306 22706 22318
rect 23886 22306 23938 22318
rect 29822 22306 29874 22318
rect 31390 22370 31442 22382
rect 31390 22306 31442 22318
rect 31614 22370 31666 22382
rect 31614 22306 31666 22318
rect 32286 22370 32338 22382
rect 32286 22306 32338 22318
rect 1710 22258 1762 22270
rect 1710 22194 1762 22206
rect 2046 22258 2098 22270
rect 2046 22194 2098 22206
rect 9214 22258 9266 22270
rect 9214 22194 9266 22206
rect 9550 22258 9602 22270
rect 9550 22194 9602 22206
rect 11566 22258 11618 22270
rect 11566 22194 11618 22206
rect 14142 22258 14194 22270
rect 16270 22258 16322 22270
rect 14802 22206 14814 22258
rect 14866 22206 14878 22258
rect 15474 22206 15486 22258
rect 15538 22206 15550 22258
rect 14142 22194 14194 22206
rect 16270 22194 16322 22206
rect 18734 22258 18786 22270
rect 18734 22194 18786 22206
rect 19630 22258 19682 22270
rect 19630 22194 19682 22206
rect 20414 22258 20466 22270
rect 20414 22194 20466 22206
rect 21870 22258 21922 22270
rect 21870 22194 21922 22206
rect 22542 22258 22594 22270
rect 22542 22194 22594 22206
rect 23550 22258 23602 22270
rect 23550 22194 23602 22206
rect 24334 22258 24386 22270
rect 24334 22194 24386 22206
rect 24670 22258 24722 22270
rect 24670 22194 24722 22206
rect 25902 22258 25954 22270
rect 25902 22194 25954 22206
rect 26014 22258 26066 22270
rect 26798 22258 26850 22270
rect 26450 22206 26462 22258
rect 26514 22206 26526 22258
rect 26014 22194 26066 22206
rect 26798 22194 26850 22206
rect 27134 22258 27186 22270
rect 27134 22194 27186 22206
rect 27470 22258 27522 22270
rect 27470 22194 27522 22206
rect 27806 22258 27858 22270
rect 27806 22194 27858 22206
rect 28254 22258 28306 22270
rect 28254 22194 28306 22206
rect 28590 22258 28642 22270
rect 28590 22194 28642 22206
rect 37214 22258 37266 22270
rect 37214 22194 37266 22206
rect 37886 22258 37938 22270
rect 37886 22194 37938 22206
rect 38222 22258 38274 22270
rect 38222 22194 38274 22206
rect 2382 22146 2434 22158
rect 2382 22082 2434 22094
rect 10446 22146 10498 22158
rect 10446 22082 10498 22094
rect 11230 22146 11282 22158
rect 11230 22082 11282 22094
rect 12014 22146 12066 22158
rect 12014 22082 12066 22094
rect 15822 22146 15874 22158
rect 15822 22082 15874 22094
rect 17278 22146 17330 22158
rect 17278 22082 17330 22094
rect 20078 22146 20130 22158
rect 20078 22082 20130 22094
rect 20750 22146 20802 22158
rect 37550 22146 37602 22158
rect 32834 22094 32846 22146
rect 32898 22094 32910 22146
rect 20750 22082 20802 22094
rect 37550 22082 37602 22094
rect 1344 21978 38800 22012
rect 1344 21926 10538 21978
rect 10590 21926 10642 21978
rect 10694 21926 10746 21978
rect 10798 21926 19862 21978
rect 19914 21926 19966 21978
rect 20018 21926 20070 21978
rect 20122 21926 29186 21978
rect 29238 21926 29290 21978
rect 29342 21926 29394 21978
rect 29446 21926 38510 21978
rect 38562 21926 38614 21978
rect 38666 21926 38718 21978
rect 38770 21926 38800 21978
rect 1344 21892 38800 21926
rect 9998 21810 10050 21822
rect 9998 21746 10050 21758
rect 13246 21810 13298 21822
rect 13246 21746 13298 21758
rect 16718 21810 16770 21822
rect 16718 21746 16770 21758
rect 17726 21810 17778 21822
rect 17726 21746 17778 21758
rect 19294 21810 19346 21822
rect 19294 21746 19346 21758
rect 21982 21810 22034 21822
rect 21982 21746 22034 21758
rect 24222 21810 24274 21822
rect 28926 21810 28978 21822
rect 27122 21758 27134 21810
rect 27186 21758 27198 21810
rect 24222 21746 24274 21758
rect 28926 21746 28978 21758
rect 1710 21698 1762 21710
rect 1710 21634 1762 21646
rect 11006 21698 11058 21710
rect 20302 21698 20354 21710
rect 18498 21646 18510 21698
rect 18562 21646 18574 21698
rect 11006 21634 11058 21646
rect 20302 21634 20354 21646
rect 21310 21698 21362 21710
rect 25566 21698 25618 21710
rect 23314 21646 23326 21698
rect 23378 21646 23390 21698
rect 23650 21646 23662 21698
rect 23714 21646 23726 21698
rect 21310 21634 21362 21646
rect 25566 21634 25618 21646
rect 26462 21698 26514 21710
rect 26462 21634 26514 21646
rect 26686 21698 26738 21710
rect 26686 21634 26738 21646
rect 27806 21698 27858 21710
rect 27806 21634 27858 21646
rect 30158 21698 30210 21710
rect 30158 21634 30210 21646
rect 32398 21698 32450 21710
rect 32398 21634 32450 21646
rect 37886 21698 37938 21710
rect 37886 21634 37938 21646
rect 38222 21698 38274 21710
rect 38222 21634 38274 21646
rect 2046 21586 2098 21598
rect 2046 21522 2098 21534
rect 9998 21586 10050 21598
rect 9998 21522 10050 21534
rect 10558 21586 10610 21598
rect 12350 21586 12402 21598
rect 11218 21534 11230 21586
rect 11282 21534 11294 21586
rect 10558 21522 10610 21534
rect 12350 21522 12402 21534
rect 12798 21586 12850 21598
rect 12798 21522 12850 21534
rect 12910 21586 12962 21598
rect 15262 21586 15314 21598
rect 17390 21586 17442 21598
rect 13458 21534 13470 21586
rect 13522 21534 13534 21586
rect 15474 21534 15486 21586
rect 15538 21534 15550 21586
rect 12910 21522 12962 21534
rect 15262 21522 15314 21534
rect 17390 21522 17442 21534
rect 18062 21586 18114 21598
rect 18062 21522 18114 21534
rect 18286 21586 18338 21598
rect 18286 21522 18338 21534
rect 18846 21586 18898 21598
rect 19966 21586 20018 21598
rect 19506 21534 19518 21586
rect 19570 21534 19582 21586
rect 18846 21522 18898 21534
rect 19966 21522 20018 21534
rect 20974 21586 21026 21598
rect 23214 21586 23266 21598
rect 21746 21534 21758 21586
rect 21810 21534 21822 21586
rect 20974 21522 21026 21534
rect 23214 21522 23266 21534
rect 23998 21586 24050 21598
rect 23998 21522 24050 21534
rect 25230 21586 25282 21598
rect 25230 21522 25282 21534
rect 26574 21586 26626 21598
rect 27694 21586 27746 21598
rect 28590 21586 28642 21598
rect 27458 21534 27470 21586
rect 27522 21534 27534 21586
rect 28242 21534 28254 21586
rect 28306 21534 28318 21586
rect 29922 21534 29934 21586
rect 29986 21534 29998 21586
rect 32162 21534 32174 21586
rect 32226 21534 32238 21586
rect 26574 21522 26626 21534
rect 27694 21522 27746 21534
rect 28590 21522 28642 21534
rect 12238 21474 12290 21486
rect 12238 21410 12290 21422
rect 15934 21474 15986 21486
rect 15934 21410 15986 21422
rect 16382 21474 16434 21486
rect 16382 21410 16434 21422
rect 16830 21474 16882 21486
rect 16830 21410 16882 21422
rect 19070 21474 19122 21486
rect 19070 21410 19122 21422
rect 22430 21474 22482 21486
rect 22430 21410 22482 21422
rect 22878 21474 22930 21486
rect 22878 21410 22930 21422
rect 10110 21362 10162 21374
rect 10110 21298 10162 21310
rect 10334 21362 10386 21374
rect 10334 21298 10386 21310
rect 12574 21362 12626 21374
rect 12574 21298 12626 21310
rect 14926 21362 14978 21374
rect 14926 21298 14978 21310
rect 15038 21362 15090 21374
rect 15038 21298 15090 21310
rect 1344 21194 38640 21228
rect 1344 21142 5876 21194
rect 5928 21142 5980 21194
rect 6032 21142 6084 21194
rect 6136 21142 15200 21194
rect 15252 21142 15304 21194
rect 15356 21142 15408 21194
rect 15460 21142 24524 21194
rect 24576 21142 24628 21194
rect 24680 21142 24732 21194
rect 24784 21142 33848 21194
rect 33900 21142 33952 21194
rect 34004 21142 34056 21194
rect 34108 21142 38640 21194
rect 1344 21108 38640 21142
rect 9998 21026 10050 21038
rect 9998 20962 10050 20974
rect 10110 21026 10162 21038
rect 10110 20962 10162 20974
rect 10670 21026 10722 21038
rect 10670 20962 10722 20974
rect 12238 21026 12290 21038
rect 12238 20962 12290 20974
rect 12350 21026 12402 21038
rect 12350 20962 12402 20974
rect 12798 21026 12850 21038
rect 12798 20962 12850 20974
rect 19406 21026 19458 21038
rect 19406 20962 19458 20974
rect 24334 21026 24386 21038
rect 24334 20962 24386 20974
rect 29486 21026 29538 21038
rect 31390 21026 31442 21038
rect 30146 20974 30158 21026
rect 30210 20974 30222 21026
rect 29486 20962 29538 20974
rect 31390 20962 31442 20974
rect 10334 20914 10386 20926
rect 10334 20850 10386 20862
rect 12574 20914 12626 20926
rect 12574 20850 12626 20862
rect 14366 20914 14418 20926
rect 17390 20914 17442 20926
rect 15586 20862 15598 20914
rect 15650 20862 15662 20914
rect 14366 20850 14418 20862
rect 17390 20850 17442 20862
rect 17726 20914 17778 20926
rect 17726 20850 17778 20862
rect 20750 20914 20802 20926
rect 20750 20850 20802 20862
rect 23326 20914 23378 20926
rect 23326 20850 23378 20862
rect 30494 20914 30546 20926
rect 30494 20850 30546 20862
rect 32286 20914 32338 20926
rect 32286 20850 32338 20862
rect 10558 20802 10610 20814
rect 10558 20738 10610 20750
rect 13470 20802 13522 20814
rect 14590 20802 14642 20814
rect 14130 20750 14142 20802
rect 14194 20750 14206 20802
rect 13470 20738 13522 20750
rect 14590 20738 14642 20750
rect 14926 20802 14978 20814
rect 15822 20802 15874 20814
rect 18398 20802 18450 20814
rect 15698 20750 15710 20802
rect 15762 20750 15774 20802
rect 16818 20750 16830 20802
rect 16882 20750 16894 20802
rect 14926 20738 14978 20750
rect 15822 20738 15874 20750
rect 18398 20738 18450 20750
rect 18734 20802 18786 20814
rect 24110 20802 24162 20814
rect 19058 20750 19070 20802
rect 19122 20750 19134 20802
rect 18734 20738 18786 20750
rect 24110 20738 24162 20750
rect 29262 20802 29314 20814
rect 29262 20738 29314 20750
rect 30718 20802 30770 20814
rect 30718 20738 30770 20750
rect 31166 20802 31218 20814
rect 31166 20738 31218 20750
rect 32062 20802 32114 20814
rect 32062 20738 32114 20750
rect 37886 20802 37938 20814
rect 37886 20738 37938 20750
rect 2046 20690 2098 20702
rect 2046 20626 2098 20638
rect 11006 20690 11058 20702
rect 11006 20626 11058 20638
rect 11342 20690 11394 20702
rect 11342 20626 11394 20638
rect 12910 20690 12962 20702
rect 17838 20690 17890 20702
rect 19854 20690 19906 20702
rect 13794 20638 13806 20690
rect 13858 20638 13870 20690
rect 16594 20638 16606 20690
rect 16658 20638 16670 20690
rect 18498 20638 18510 20690
rect 18562 20638 18574 20690
rect 12910 20626 12962 20638
rect 17838 20626 17890 20638
rect 19854 20626 19906 20638
rect 20190 20690 20242 20702
rect 20190 20626 20242 20638
rect 21310 20690 21362 20702
rect 21310 20626 21362 20638
rect 21982 20690 22034 20702
rect 21982 20626 22034 20638
rect 22766 20690 22818 20702
rect 22766 20626 22818 20638
rect 23550 20690 23602 20702
rect 24894 20690 24946 20702
rect 23762 20638 23774 20690
rect 23826 20638 23838 20690
rect 23550 20626 23602 20638
rect 24894 20626 24946 20638
rect 25230 20690 25282 20702
rect 25230 20626 25282 20638
rect 26014 20690 26066 20702
rect 26014 20626 26066 20638
rect 26350 20690 26402 20702
rect 26350 20626 26402 20638
rect 27694 20690 27746 20702
rect 27694 20626 27746 20638
rect 28030 20690 28082 20702
rect 32958 20690 33010 20702
rect 31714 20638 31726 20690
rect 31778 20638 31790 20690
rect 28030 20626 28082 20638
rect 32958 20626 33010 20638
rect 33294 20690 33346 20702
rect 33294 20626 33346 20638
rect 1710 20578 1762 20590
rect 1710 20514 1762 20526
rect 14254 20578 14306 20590
rect 14254 20514 14306 20526
rect 17278 20578 17330 20590
rect 17278 20514 17330 20526
rect 21646 20578 21698 20590
rect 21646 20514 21698 20526
rect 22318 20578 22370 20590
rect 38222 20578 38274 20590
rect 29810 20526 29822 20578
rect 29874 20526 29886 20578
rect 32610 20526 32622 20578
rect 32674 20526 32686 20578
rect 22318 20514 22370 20526
rect 38222 20514 38274 20526
rect 1344 20410 38800 20444
rect 1344 20358 10538 20410
rect 10590 20358 10642 20410
rect 10694 20358 10746 20410
rect 10798 20358 19862 20410
rect 19914 20358 19966 20410
rect 20018 20358 20070 20410
rect 20122 20358 29186 20410
rect 29238 20358 29290 20410
rect 29342 20358 29394 20410
rect 29446 20358 38510 20410
rect 38562 20358 38614 20410
rect 38666 20358 38718 20410
rect 38770 20358 38800 20410
rect 1344 20324 38800 20358
rect 10558 20242 10610 20254
rect 10558 20178 10610 20190
rect 12238 20242 12290 20254
rect 12238 20178 12290 20190
rect 19518 20242 19570 20254
rect 19518 20178 19570 20190
rect 19854 20242 19906 20254
rect 19854 20178 19906 20190
rect 24334 20242 24386 20254
rect 27570 20190 27582 20242
rect 27634 20190 27646 20242
rect 24334 20178 24386 20190
rect 9886 20130 9938 20142
rect 2034 20078 2046 20130
rect 2098 20078 2110 20130
rect 9886 20066 9938 20078
rect 11566 20130 11618 20142
rect 11566 20066 11618 20078
rect 12574 20130 12626 20142
rect 12574 20066 12626 20078
rect 12910 20130 12962 20142
rect 15038 20130 15090 20142
rect 13570 20078 13582 20130
rect 13634 20078 13646 20130
rect 14130 20078 14142 20130
rect 14194 20078 14206 20130
rect 12910 20066 12962 20078
rect 15038 20066 15090 20078
rect 17502 20130 17554 20142
rect 17502 20066 17554 20078
rect 17838 20130 17890 20142
rect 17838 20066 17890 20078
rect 18846 20130 18898 20142
rect 18846 20066 18898 20078
rect 21198 20130 21250 20142
rect 21198 20066 21250 20078
rect 21646 20130 21698 20142
rect 21646 20066 21698 20078
rect 22318 20130 22370 20142
rect 22318 20066 22370 20078
rect 22990 20130 23042 20142
rect 25566 20130 25618 20142
rect 23762 20078 23774 20130
rect 23826 20078 23838 20130
rect 22990 20066 23042 20078
rect 25566 20066 25618 20078
rect 27134 20130 27186 20142
rect 27134 20066 27186 20078
rect 28590 20130 28642 20142
rect 28590 20066 28642 20078
rect 29822 20130 29874 20142
rect 29822 20066 29874 20078
rect 30158 20130 30210 20142
rect 30158 20066 30210 20078
rect 32174 20130 32226 20142
rect 32174 20066 32226 20078
rect 38222 20130 38274 20142
rect 38222 20066 38274 20078
rect 1710 20018 1762 20030
rect 11230 20018 11282 20030
rect 13246 20018 13298 20030
rect 9650 19966 9662 20018
rect 9714 19966 9726 20018
rect 10322 19966 10334 20018
rect 10386 19966 10398 20018
rect 12002 19966 12014 20018
rect 12066 19966 12078 20018
rect 1710 19954 1762 19966
rect 11230 19954 11282 19966
rect 13246 19954 13298 19966
rect 14478 20018 14530 20030
rect 14478 19954 14530 19966
rect 15150 20018 15202 20030
rect 15150 19954 15202 19966
rect 15374 20018 15426 20030
rect 16382 20018 16434 20030
rect 15586 19966 15598 20018
rect 15650 19966 15662 20018
rect 15374 19954 15426 19966
rect 16382 19954 16434 19966
rect 16830 20018 16882 20030
rect 16830 19954 16882 19966
rect 18734 20018 18786 20030
rect 20862 20018 20914 20030
rect 19058 19966 19070 20018
rect 19122 19966 19134 20018
rect 18734 19954 18786 19966
rect 20862 19954 20914 19966
rect 21982 20018 22034 20030
rect 23326 20018 23378 20030
rect 22754 19966 22766 20018
rect 22818 19966 22830 20018
rect 21982 19954 22034 19966
rect 23326 19954 23378 19966
rect 23550 20018 23602 20030
rect 23550 19954 23602 19966
rect 24110 20018 24162 20030
rect 24110 19954 24162 19966
rect 25230 20018 25282 20030
rect 25230 19954 25282 19966
rect 26910 20018 26962 20030
rect 26910 19954 26962 19966
rect 27022 20018 27074 20030
rect 27022 19954 27074 19966
rect 28254 20018 28306 20030
rect 37886 20018 37938 20030
rect 31938 19966 31950 20018
rect 32002 19966 32014 20018
rect 28254 19954 28306 19966
rect 37886 19954 37938 19966
rect 2494 19906 2546 19918
rect 2494 19842 2546 19854
rect 18510 19906 18562 19918
rect 18510 19842 18562 19854
rect 20526 19906 20578 19918
rect 20526 19842 20578 19854
rect 1344 19626 38640 19660
rect 1344 19574 5876 19626
rect 5928 19574 5980 19626
rect 6032 19574 6084 19626
rect 6136 19574 15200 19626
rect 15252 19574 15304 19626
rect 15356 19574 15408 19626
rect 15460 19574 24524 19626
rect 24576 19574 24628 19626
rect 24680 19574 24732 19626
rect 24784 19574 33848 19626
rect 33900 19574 33952 19626
rect 34004 19574 34056 19626
rect 34108 19574 38640 19626
rect 1344 19540 38640 19574
rect 24782 19458 24834 19470
rect 24782 19394 24834 19406
rect 17838 19234 17890 19246
rect 10546 19182 10558 19234
rect 10610 19182 10622 19234
rect 12674 19182 12686 19234
rect 12738 19182 12750 19234
rect 17838 19170 17890 19182
rect 18510 19234 18562 19246
rect 18510 19170 18562 19182
rect 18846 19234 18898 19246
rect 23774 19234 23826 19246
rect 19058 19182 19070 19234
rect 19122 19182 19134 19234
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 22418 19182 22430 19234
rect 22482 19182 22494 19234
rect 23202 19182 23214 19234
rect 23266 19182 23278 19234
rect 18846 19170 18898 19182
rect 23774 19170 23826 19182
rect 23998 19234 24050 19246
rect 23998 19170 24050 19182
rect 24110 19234 24162 19246
rect 25902 19234 25954 19246
rect 24322 19182 24334 19234
rect 24386 19182 24398 19234
rect 24110 19170 24162 19182
rect 25902 19170 25954 19182
rect 26574 19234 26626 19246
rect 27582 19234 27634 19246
rect 27346 19182 27358 19234
rect 27410 19182 27422 19234
rect 30370 19182 30382 19234
rect 30434 19182 30446 19234
rect 31938 19182 31950 19234
rect 32002 19182 32014 19234
rect 26574 19170 26626 19182
rect 27582 19170 27634 19182
rect 11454 19122 11506 19134
rect 10770 19070 10782 19122
rect 10834 19070 10846 19122
rect 11454 19058 11506 19070
rect 14702 19122 14754 19134
rect 14702 19058 14754 19070
rect 15038 19122 15090 19134
rect 15038 19058 15090 19070
rect 15598 19122 15650 19134
rect 15598 19058 15650 19070
rect 15934 19122 15986 19134
rect 15934 19058 15986 19070
rect 16270 19122 16322 19134
rect 16270 19058 16322 19070
rect 16606 19122 16658 19134
rect 16606 19058 16658 19070
rect 16942 19122 16994 19134
rect 16942 19058 16994 19070
rect 17278 19122 17330 19134
rect 17278 19058 17330 19070
rect 18174 19122 18226 19134
rect 18174 19058 18226 19070
rect 18734 19122 18786 19134
rect 18734 19058 18786 19070
rect 19518 19122 19570 19134
rect 19518 19058 19570 19070
rect 19742 19122 19794 19134
rect 19742 19058 19794 19070
rect 20526 19122 20578 19134
rect 20526 19058 20578 19070
rect 22654 19122 22706 19134
rect 22654 19058 22706 19070
rect 23438 19122 23490 19134
rect 23438 19058 23490 19070
rect 26910 19122 26962 19134
rect 26910 19058 26962 19070
rect 27694 19122 27746 19134
rect 29150 19122 29202 19134
rect 28130 19070 28142 19122
rect 28194 19070 28206 19122
rect 27694 19058 27746 19070
rect 29150 19058 29202 19070
rect 30942 19122 30994 19134
rect 30942 19058 30994 19070
rect 37886 19122 37938 19134
rect 37886 19058 37938 19070
rect 1710 19010 1762 19022
rect 2494 19010 2546 19022
rect 2034 18958 2046 19010
rect 2098 18958 2110 19010
rect 1710 18946 1762 18958
rect 2494 18946 2546 18958
rect 11118 19010 11170 19022
rect 11118 18946 11170 18958
rect 12910 19010 12962 19022
rect 12910 18946 12962 18958
rect 14366 19010 14418 19022
rect 14366 18946 14418 18958
rect 20078 19010 20130 19022
rect 20078 18946 20130 18958
rect 21310 19010 21362 19022
rect 21310 18946 21362 18958
rect 25230 19010 25282 19022
rect 25230 18946 25282 18958
rect 26238 19010 26290 19022
rect 26238 18946 26290 18958
rect 29486 19010 29538 19022
rect 29486 18946 29538 18958
rect 30606 19010 30658 19022
rect 30606 18946 30658 18958
rect 31278 19010 31330 19022
rect 31278 18946 31330 18958
rect 32174 19010 32226 19022
rect 32174 18946 32226 18958
rect 38222 19010 38274 19022
rect 38222 18946 38274 18958
rect 1344 18842 38800 18876
rect 1344 18790 10538 18842
rect 10590 18790 10642 18842
rect 10694 18790 10746 18842
rect 10798 18790 19862 18842
rect 19914 18790 19966 18842
rect 20018 18790 20070 18842
rect 20122 18790 29186 18842
rect 29238 18790 29290 18842
rect 29342 18790 29394 18842
rect 29446 18790 38510 18842
rect 38562 18790 38614 18842
rect 38666 18790 38718 18842
rect 38770 18790 38800 18842
rect 1344 18756 38800 18790
rect 16830 18674 16882 18686
rect 16830 18610 16882 18622
rect 18062 18674 18114 18686
rect 22430 18674 22482 18686
rect 20178 18622 20190 18674
rect 20242 18622 20254 18674
rect 18062 18610 18114 18622
rect 22430 18610 22482 18622
rect 23662 18674 23714 18686
rect 28018 18622 28030 18674
rect 28082 18622 28094 18674
rect 30482 18622 30494 18674
rect 30546 18622 30558 18674
rect 31938 18622 31950 18674
rect 32002 18622 32014 18674
rect 23662 18610 23714 18622
rect 1710 18562 1762 18574
rect 1710 18498 1762 18510
rect 10894 18562 10946 18574
rect 10894 18498 10946 18510
rect 11566 18562 11618 18574
rect 11566 18498 11618 18510
rect 13358 18562 13410 18574
rect 13358 18498 13410 18510
rect 14814 18562 14866 18574
rect 14814 18498 14866 18510
rect 18734 18562 18786 18574
rect 18734 18498 18786 18510
rect 21646 18562 21698 18574
rect 21646 18498 21698 18510
rect 22654 18562 22706 18574
rect 22654 18498 22706 18510
rect 24334 18562 24386 18574
rect 24334 18498 24386 18510
rect 25790 18562 25842 18574
rect 25790 18498 25842 18510
rect 26126 18562 26178 18574
rect 26126 18498 26178 18510
rect 26462 18562 26514 18574
rect 26462 18498 26514 18510
rect 27358 18562 27410 18574
rect 27358 18498 27410 18510
rect 27582 18562 27634 18574
rect 27582 18498 27634 18510
rect 38222 18562 38274 18574
rect 38222 18498 38274 18510
rect 2046 18450 2098 18462
rect 2046 18386 2098 18398
rect 10446 18450 10498 18462
rect 11902 18450 11954 18462
rect 12910 18450 12962 18462
rect 11106 18398 11118 18450
rect 11170 18398 11182 18450
rect 12226 18398 12238 18450
rect 12290 18398 12302 18450
rect 10446 18386 10498 18398
rect 11902 18386 11954 18398
rect 12910 18386 12962 18398
rect 13022 18450 13074 18462
rect 13022 18386 13074 18398
rect 13694 18450 13746 18462
rect 13694 18386 13746 18398
rect 14478 18450 14530 18462
rect 14478 18386 14530 18398
rect 15374 18450 15426 18462
rect 15374 18386 15426 18398
rect 17614 18450 17666 18462
rect 17614 18386 17666 18398
rect 18398 18450 18450 18462
rect 19854 18450 19906 18462
rect 18946 18398 18958 18450
rect 19010 18398 19022 18450
rect 18398 18386 18450 18398
rect 19854 18386 19906 18398
rect 21422 18450 21474 18462
rect 21422 18386 21474 18398
rect 21758 18450 21810 18462
rect 21758 18386 21810 18398
rect 22206 18450 22258 18462
rect 23326 18450 23378 18462
rect 25454 18450 25506 18462
rect 22866 18398 22878 18450
rect 22930 18398 22942 18450
rect 24098 18398 24110 18450
rect 24162 18398 24174 18450
rect 22206 18386 22258 18398
rect 23326 18386 23378 18398
rect 25454 18386 25506 18398
rect 27470 18450 27522 18462
rect 27470 18386 27522 18398
rect 29598 18450 29650 18462
rect 31054 18450 31106 18462
rect 30146 18398 30158 18450
rect 30210 18398 30222 18450
rect 29598 18386 29650 18398
rect 31054 18386 31106 18398
rect 37886 18450 37938 18462
rect 37886 18386 37938 18398
rect 14254 18338 14306 18350
rect 14254 18274 14306 18286
rect 16158 18338 16210 18350
rect 16158 18274 16210 18286
rect 19518 18338 19570 18350
rect 19518 18274 19570 18286
rect 21086 18338 21138 18350
rect 21086 18274 21138 18286
rect 31390 18338 31442 18350
rect 31390 18274 31442 18286
rect 9886 18226 9938 18238
rect 9886 18162 9938 18174
rect 9998 18226 10050 18238
rect 9998 18162 10050 18174
rect 10222 18226 10274 18238
rect 10222 18162 10274 18174
rect 10558 18226 10610 18238
rect 10558 18162 10610 18174
rect 12462 18226 12514 18238
rect 12462 18162 12514 18174
rect 12686 18226 12738 18238
rect 12686 18162 12738 18174
rect 15262 18226 15314 18238
rect 15262 18162 15314 18174
rect 16046 18226 16098 18238
rect 16046 18162 16098 18174
rect 29822 18226 29874 18238
rect 29822 18162 29874 18174
rect 30830 18226 30882 18238
rect 30830 18162 30882 18174
rect 31614 18226 31666 18238
rect 31614 18162 31666 18174
rect 1344 18058 38640 18092
rect 1344 18006 5876 18058
rect 5928 18006 5980 18058
rect 6032 18006 6084 18058
rect 6136 18006 15200 18058
rect 15252 18006 15304 18058
rect 15356 18006 15408 18058
rect 15460 18006 24524 18058
rect 24576 18006 24628 18058
rect 24680 18006 24732 18058
rect 24784 18006 33848 18058
rect 33900 18006 33952 18058
rect 34004 18006 34056 18058
rect 34108 18006 38640 18058
rect 1344 17972 38640 18006
rect 10222 17890 10274 17902
rect 10222 17826 10274 17838
rect 10446 17890 10498 17902
rect 10446 17826 10498 17838
rect 10670 17890 10722 17902
rect 10670 17826 10722 17838
rect 10782 17890 10834 17902
rect 10782 17826 10834 17838
rect 12238 17890 12290 17902
rect 12238 17826 12290 17838
rect 12910 17890 12962 17902
rect 12910 17826 12962 17838
rect 14702 17890 14754 17902
rect 14702 17826 14754 17838
rect 15710 17890 15762 17902
rect 15710 17826 15762 17838
rect 25342 17890 25394 17902
rect 25342 17826 25394 17838
rect 19406 17778 19458 17790
rect 19406 17714 19458 17726
rect 24222 17778 24274 17790
rect 24222 17714 24274 17726
rect 26350 17778 26402 17790
rect 26350 17714 26402 17726
rect 2718 17666 2770 17678
rect 2718 17602 2770 17614
rect 8766 17666 8818 17678
rect 8766 17602 8818 17614
rect 10110 17666 10162 17678
rect 12350 17666 12402 17678
rect 11330 17614 11342 17666
rect 11394 17614 11406 17666
rect 10110 17602 10162 17614
rect 12350 17602 12402 17614
rect 12574 17666 12626 17678
rect 12574 17602 12626 17614
rect 12798 17666 12850 17678
rect 12798 17602 12850 17614
rect 14814 17666 14866 17678
rect 14814 17602 14866 17614
rect 15038 17666 15090 17678
rect 15934 17666 15986 17678
rect 15474 17614 15486 17666
rect 15538 17614 15550 17666
rect 15038 17602 15090 17614
rect 15934 17602 15986 17614
rect 16606 17666 16658 17678
rect 16606 17602 16658 17614
rect 18174 17666 18226 17678
rect 18174 17602 18226 17614
rect 18286 17666 18338 17678
rect 21758 17666 21810 17678
rect 18610 17614 18622 17666
rect 18674 17614 18686 17666
rect 18286 17602 18338 17614
rect 21758 17602 21810 17614
rect 22766 17666 22818 17678
rect 25566 17666 25618 17678
rect 24882 17614 24894 17666
rect 24946 17614 24958 17666
rect 22766 17602 22818 17614
rect 25566 17602 25618 17614
rect 27246 17666 27298 17678
rect 27246 17602 27298 17614
rect 27470 17666 27522 17678
rect 27470 17602 27522 17614
rect 31166 17666 31218 17678
rect 31166 17602 31218 17614
rect 31390 17666 31442 17678
rect 31390 17602 31442 17614
rect 37214 17666 37266 17678
rect 37214 17602 37266 17614
rect 1710 17554 1762 17566
rect 1710 17490 1762 17502
rect 2046 17554 2098 17566
rect 2046 17490 2098 17502
rect 8430 17554 8482 17566
rect 8430 17490 8482 17502
rect 15150 17554 15202 17566
rect 15150 17490 15202 17502
rect 17726 17554 17778 17566
rect 17726 17490 17778 17502
rect 18398 17554 18450 17566
rect 18398 17490 18450 17502
rect 19742 17554 19794 17566
rect 19742 17490 19794 17502
rect 20078 17554 20130 17566
rect 20078 17490 20130 17502
rect 23438 17554 23490 17566
rect 23438 17490 23490 17502
rect 23774 17554 23826 17566
rect 26126 17554 26178 17566
rect 24322 17502 24334 17554
rect 24386 17502 24398 17554
rect 24658 17502 24670 17554
rect 24722 17502 24734 17554
rect 25890 17502 25902 17554
rect 25954 17502 25966 17554
rect 23774 17490 23826 17502
rect 26126 17490 26178 17502
rect 27358 17554 27410 17566
rect 28254 17554 28306 17566
rect 27906 17502 27918 17554
rect 27970 17502 27982 17554
rect 27358 17490 27410 17502
rect 28254 17490 28306 17502
rect 28590 17554 28642 17566
rect 28590 17490 28642 17502
rect 29150 17554 29202 17566
rect 29150 17490 29202 17502
rect 29486 17554 29538 17566
rect 32062 17554 32114 17566
rect 31714 17502 31726 17554
rect 31778 17502 31790 17554
rect 29486 17490 29538 17502
rect 32062 17490 32114 17502
rect 32398 17554 32450 17566
rect 32398 17490 32450 17502
rect 37886 17554 37938 17566
rect 37886 17490 37938 17502
rect 38222 17554 38274 17566
rect 38222 17490 38274 17502
rect 2382 17442 2434 17454
rect 2382 17378 2434 17390
rect 11118 17442 11170 17454
rect 11118 17378 11170 17390
rect 15598 17442 15650 17454
rect 15598 17378 15650 17390
rect 16942 17442 16994 17454
rect 16942 17378 16994 17390
rect 17390 17442 17442 17454
rect 17390 17378 17442 17390
rect 19070 17442 19122 17454
rect 19070 17378 19122 17390
rect 22094 17442 22146 17454
rect 22094 17378 22146 17390
rect 23102 17442 23154 17454
rect 23102 17378 23154 17390
rect 25230 17442 25282 17454
rect 25230 17378 25282 17390
rect 37550 17442 37602 17454
rect 37550 17378 37602 17390
rect 1344 17274 38800 17308
rect 1344 17222 10538 17274
rect 10590 17222 10642 17274
rect 10694 17222 10746 17274
rect 10798 17222 19862 17274
rect 19914 17222 19966 17274
rect 20018 17222 20070 17274
rect 20122 17222 29186 17274
rect 29238 17222 29290 17274
rect 29342 17222 29394 17274
rect 29446 17222 38510 17274
rect 38562 17222 38614 17274
rect 38666 17222 38718 17274
rect 38770 17222 38800 17274
rect 1344 17188 38800 17222
rect 18398 17106 18450 17118
rect 18398 17042 18450 17054
rect 21646 17106 21698 17118
rect 21646 17042 21698 17054
rect 23662 17106 23714 17118
rect 23662 17042 23714 17054
rect 25678 17106 25730 17118
rect 25678 17042 25730 17054
rect 1710 16994 1762 17006
rect 1710 16930 1762 16942
rect 2046 16994 2098 17006
rect 2046 16930 2098 16942
rect 10782 16994 10834 17006
rect 10782 16930 10834 16942
rect 13358 16994 13410 17006
rect 13358 16930 13410 16942
rect 16494 16994 16546 17006
rect 16494 16930 16546 16942
rect 17614 16994 17666 17006
rect 19070 16994 19122 17006
rect 17826 16942 17838 16994
rect 17890 16942 17902 16994
rect 17614 16930 17666 16942
rect 19070 16930 19122 16942
rect 19406 16994 19458 17006
rect 19406 16930 19458 16942
rect 19966 16994 20018 17006
rect 21982 16994 22034 17006
rect 20626 16942 20638 16994
rect 20690 16942 20702 16994
rect 19966 16930 20018 16942
rect 21982 16930 22034 16942
rect 22318 16994 22370 17006
rect 22318 16930 22370 16942
rect 22878 16994 22930 17006
rect 22878 16930 22930 16942
rect 23214 16994 23266 17006
rect 23214 16930 23266 16942
rect 25342 16994 25394 17006
rect 25342 16930 25394 16942
rect 26574 16994 26626 17006
rect 26574 16930 26626 16942
rect 27246 16994 27298 17006
rect 27246 16930 27298 16942
rect 28366 16994 28418 17006
rect 28366 16930 28418 16942
rect 29150 16994 29202 17006
rect 29150 16930 29202 16942
rect 30718 16994 30770 17006
rect 30718 16930 30770 16942
rect 32510 16994 32562 17006
rect 32510 16930 32562 16942
rect 38222 16994 38274 17006
rect 38222 16930 38274 16942
rect 10222 16882 10274 16894
rect 13022 16882 13074 16894
rect 14702 16882 14754 16894
rect 12226 16830 12238 16882
rect 12290 16830 12302 16882
rect 13570 16830 13582 16882
rect 13634 16830 13646 16882
rect 10222 16818 10274 16830
rect 13022 16818 13074 16830
rect 14702 16818 14754 16830
rect 15038 16882 15090 16894
rect 15934 16882 15986 16894
rect 15474 16830 15486 16882
rect 15538 16830 15550 16882
rect 15038 16818 15090 16830
rect 15934 16818 15986 16830
rect 17390 16882 17442 16894
rect 17390 16818 17442 16830
rect 18174 16882 18226 16894
rect 20974 16882 21026 16894
rect 26238 16882 26290 16894
rect 27134 16882 27186 16894
rect 28030 16882 28082 16894
rect 29486 16882 29538 16894
rect 30382 16882 30434 16894
rect 20178 16830 20190 16882
rect 20242 16830 20254 16882
rect 21410 16830 21422 16882
rect 21474 16830 21486 16882
rect 26898 16830 26910 16882
rect 26962 16830 26974 16882
rect 27682 16830 27694 16882
rect 27746 16830 27758 16882
rect 28914 16830 28926 16882
rect 28978 16830 28990 16882
rect 30034 16830 30046 16882
rect 30098 16830 30110 16882
rect 18174 16818 18226 16830
rect 20974 16818 21026 16830
rect 26238 16818 26290 16830
rect 27134 16818 27186 16830
rect 28030 16818 28082 16830
rect 29486 16818 29538 16830
rect 30382 16818 30434 16830
rect 31278 16882 31330 16894
rect 32174 16882 32226 16894
rect 31826 16830 31838 16882
rect 31890 16830 31902 16882
rect 31278 16818 31330 16830
rect 32174 16818 32226 16830
rect 37886 16882 37938 16894
rect 37886 16818 37938 16830
rect 10446 16770 10498 16782
rect 10446 16706 10498 16718
rect 15150 16770 15202 16782
rect 15150 16706 15202 16718
rect 29710 16770 29762 16782
rect 29710 16706 29762 16718
rect 31502 16770 31554 16782
rect 31502 16706 31554 16718
rect 10110 16658 10162 16670
rect 10110 16594 10162 16606
rect 10670 16658 10722 16670
rect 10670 16594 10722 16606
rect 12462 16658 12514 16670
rect 12462 16594 12514 16606
rect 12686 16658 12738 16670
rect 12686 16594 12738 16606
rect 12910 16658 12962 16670
rect 12910 16594 12962 16606
rect 14814 16658 14866 16670
rect 14814 16594 14866 16606
rect 15710 16658 15762 16670
rect 15710 16594 15762 16606
rect 16046 16658 16098 16670
rect 16046 16594 16098 16606
rect 16382 16658 16434 16670
rect 16382 16594 16434 16606
rect 1344 16490 38640 16524
rect 1344 16438 5876 16490
rect 5928 16438 5980 16490
rect 6032 16438 6084 16490
rect 6136 16438 15200 16490
rect 15252 16438 15304 16490
rect 15356 16438 15408 16490
rect 15460 16438 24524 16490
rect 24576 16438 24628 16490
rect 24680 16438 24732 16490
rect 24784 16438 33848 16490
rect 33900 16438 33952 16490
rect 34004 16438 34056 16490
rect 34108 16438 38640 16490
rect 1344 16404 38640 16438
rect 10334 16322 10386 16334
rect 10334 16258 10386 16270
rect 10782 16322 10834 16334
rect 10782 16258 10834 16270
rect 12238 16322 12290 16334
rect 12238 16258 12290 16270
rect 15486 16322 15538 16334
rect 15486 16258 15538 16270
rect 29822 16322 29874 16334
rect 29822 16258 29874 16270
rect 31502 16322 31554 16334
rect 31502 16258 31554 16270
rect 10558 16210 10610 16222
rect 10558 16146 10610 16158
rect 12574 16210 12626 16222
rect 12574 16146 12626 16158
rect 17390 16210 17442 16222
rect 17390 16146 17442 16158
rect 17726 16210 17778 16222
rect 17726 16146 17778 16158
rect 22990 16210 23042 16222
rect 22990 16146 23042 16158
rect 24446 16210 24498 16222
rect 24446 16146 24498 16158
rect 29598 16210 29650 16222
rect 29598 16146 29650 16158
rect 31278 16210 31330 16222
rect 31278 16146 31330 16158
rect 2046 16098 2098 16110
rect 2046 16034 2098 16046
rect 8542 16098 8594 16110
rect 12350 16098 12402 16110
rect 8866 16046 8878 16098
rect 8930 16046 8942 16098
rect 9538 16046 9550 16098
rect 9602 16046 9614 16098
rect 10098 16046 10110 16098
rect 10162 16046 10174 16098
rect 8542 16034 8594 16046
rect 12350 16034 12402 16046
rect 12798 16098 12850 16110
rect 18062 16098 18114 16110
rect 18734 16098 18786 16110
rect 19742 16098 19794 16110
rect 14914 16046 14926 16098
rect 14978 16046 14990 16098
rect 16706 16046 16718 16098
rect 16770 16046 16782 16098
rect 18274 16046 18286 16098
rect 18338 16046 18350 16098
rect 19170 16046 19182 16098
rect 19234 16046 19246 16098
rect 12798 16034 12850 16046
rect 18062 16034 18114 16046
rect 18734 16034 18786 16046
rect 19742 16034 19794 16046
rect 23326 16098 23378 16110
rect 23326 16034 23378 16046
rect 23774 16098 23826 16110
rect 23774 16034 23826 16046
rect 24670 16098 24722 16110
rect 24994 16046 25006 16098
rect 25058 16046 25070 16098
rect 24670 16034 24722 16046
rect 9102 15986 9154 15998
rect 9102 15922 9154 15934
rect 9774 15986 9826 15998
rect 9774 15922 9826 15934
rect 10894 15986 10946 15998
rect 10894 15922 10946 15934
rect 11454 15986 11506 15998
rect 11454 15922 11506 15934
rect 11790 15986 11842 15998
rect 11790 15922 11842 15934
rect 12910 15986 12962 15998
rect 12910 15922 12962 15934
rect 13470 15986 13522 15998
rect 13470 15922 13522 15934
rect 13806 15986 13858 15998
rect 13806 15922 13858 15934
rect 15150 15986 15202 15998
rect 15150 15922 15202 15934
rect 15598 15986 15650 15998
rect 15598 15922 15650 15934
rect 15934 15986 15986 15998
rect 15934 15922 15986 15934
rect 16942 15986 16994 15998
rect 16942 15922 16994 15934
rect 17950 15986 18002 15998
rect 17950 15922 18002 15934
rect 21310 15986 21362 15998
rect 21310 15922 21362 15934
rect 21646 15986 21698 15998
rect 21646 15922 21698 15934
rect 22094 15986 22146 15998
rect 25454 15986 25506 15998
rect 23090 15934 23102 15986
rect 23154 15934 23166 15986
rect 24882 15934 24894 15986
rect 24946 15934 24958 15986
rect 22094 15922 22146 15934
rect 25454 15922 25506 15934
rect 25678 15986 25730 15998
rect 30494 15986 30546 15998
rect 30146 15934 30158 15986
rect 30210 15934 30222 15986
rect 25678 15922 25730 15934
rect 30494 15922 30546 15934
rect 30830 15986 30882 15998
rect 32174 15986 32226 15998
rect 31826 15934 31838 15986
rect 31890 15934 31902 15986
rect 30830 15922 30882 15934
rect 32174 15922 32226 15934
rect 37886 15986 37938 15998
rect 37886 15922 37938 15934
rect 1710 15874 1762 15886
rect 1710 15810 1762 15822
rect 14478 15874 14530 15886
rect 14478 15810 14530 15822
rect 16270 15874 16322 15886
rect 16270 15810 16322 15822
rect 18958 15874 19010 15886
rect 21982 15874 22034 15886
rect 20066 15822 20078 15874
rect 20130 15822 20142 15874
rect 18958 15810 19010 15822
rect 21982 15810 22034 15822
rect 23998 15874 24050 15886
rect 23998 15810 24050 15822
rect 26014 15874 26066 15886
rect 26014 15810 26066 15822
rect 32510 15874 32562 15886
rect 32510 15810 32562 15822
rect 38222 15874 38274 15886
rect 38222 15810 38274 15822
rect 1344 15706 38800 15740
rect 1344 15654 10538 15706
rect 10590 15654 10642 15706
rect 10694 15654 10746 15706
rect 10798 15654 19862 15706
rect 19914 15654 19966 15706
rect 20018 15654 20070 15706
rect 20122 15654 29186 15706
rect 29238 15654 29290 15706
rect 29342 15654 29394 15706
rect 29446 15654 38510 15706
rect 38562 15654 38614 15706
rect 38666 15654 38718 15706
rect 38770 15654 38800 15706
rect 1344 15620 38800 15654
rect 12462 15538 12514 15550
rect 12462 15474 12514 15486
rect 14030 15538 14082 15550
rect 14030 15474 14082 15486
rect 16046 15538 16098 15550
rect 16046 15474 16098 15486
rect 16830 15538 16882 15550
rect 23886 15538 23938 15550
rect 19394 15486 19406 15538
rect 19458 15486 19470 15538
rect 16830 15474 16882 15486
rect 23886 15474 23938 15486
rect 24558 15538 24610 15550
rect 24558 15474 24610 15486
rect 28814 15538 28866 15550
rect 28814 15474 28866 15486
rect 1710 15426 1762 15438
rect 1710 15362 1762 15374
rect 2046 15426 2098 15438
rect 2046 15362 2098 15374
rect 9998 15426 10050 15438
rect 9998 15362 10050 15374
rect 10334 15426 10386 15438
rect 10334 15362 10386 15374
rect 10670 15426 10722 15438
rect 10670 15362 10722 15374
rect 11006 15426 11058 15438
rect 11006 15362 11058 15374
rect 11342 15426 11394 15438
rect 11342 15362 11394 15374
rect 12798 15426 12850 15438
rect 12798 15362 12850 15374
rect 14926 15426 14978 15438
rect 14926 15362 14978 15374
rect 15262 15426 15314 15438
rect 15262 15362 15314 15374
rect 17614 15426 17666 15438
rect 18622 15426 18674 15438
rect 17826 15374 17838 15426
rect 17890 15374 17902 15426
rect 17614 15362 17666 15374
rect 18622 15362 18674 15374
rect 22990 15426 23042 15438
rect 22990 15362 23042 15374
rect 24222 15426 24274 15438
rect 24222 15362 24274 15374
rect 25566 15426 25618 15438
rect 25566 15362 25618 15374
rect 25902 15426 25954 15438
rect 25902 15362 25954 15374
rect 26350 15426 26402 15438
rect 26350 15362 26402 15374
rect 37886 15426 37938 15438
rect 37886 15362 37938 15374
rect 38222 15426 38274 15438
rect 38222 15362 38274 15374
rect 14590 15314 14642 15326
rect 13010 15262 13022 15314
rect 13074 15262 13086 15314
rect 14590 15250 14642 15262
rect 17502 15314 17554 15326
rect 17502 15250 17554 15262
rect 18174 15314 18226 15326
rect 18174 15250 18226 15262
rect 18398 15314 18450 15326
rect 20974 15314 21026 15326
rect 18834 15262 18846 15314
rect 18898 15262 18910 15314
rect 19618 15262 19630 15314
rect 19682 15262 19694 15314
rect 18398 15250 18450 15262
rect 20974 15250 21026 15262
rect 21086 15314 21138 15326
rect 21086 15250 21138 15262
rect 21198 15314 21250 15326
rect 21198 15250 21250 15262
rect 22318 15314 22370 15326
rect 22318 15250 22370 15262
rect 22654 15314 22706 15326
rect 26462 15314 26514 15326
rect 23650 15262 23662 15314
rect 23714 15262 23726 15314
rect 22654 15250 22706 15262
rect 26462 15250 26514 15262
rect 26574 15314 26626 15326
rect 27582 15314 27634 15326
rect 27346 15262 27358 15314
rect 27410 15262 27422 15314
rect 26574 15250 26626 15262
rect 27582 15250 27634 15262
rect 27694 15314 27746 15326
rect 28478 15314 28530 15326
rect 28130 15262 28142 15314
rect 28194 15262 28206 15314
rect 27694 15250 27746 15262
rect 28478 15250 28530 15262
rect 12014 15202 12066 15214
rect 14242 15150 14254 15202
rect 14306 15199 14318 15202
rect 14466 15199 14478 15202
rect 14306 15153 14478 15199
rect 14306 15150 14318 15153
rect 14466 15150 14478 15153
rect 14530 15150 14542 15202
rect 21634 15150 21646 15202
rect 21698 15150 21710 15202
rect 12014 15138 12066 15150
rect 27010 15038 27022 15090
rect 27074 15038 27086 15090
rect 1344 14922 38640 14956
rect 1344 14870 5876 14922
rect 5928 14870 5980 14922
rect 6032 14870 6084 14922
rect 6136 14870 15200 14922
rect 15252 14870 15304 14922
rect 15356 14870 15408 14922
rect 15460 14870 24524 14922
rect 24576 14870 24628 14922
rect 24680 14870 24732 14922
rect 24784 14870 33848 14922
rect 33900 14870 33952 14922
rect 34004 14870 34056 14922
rect 34108 14870 38640 14922
rect 1344 14836 38640 14870
rect 10446 14754 10498 14766
rect 10446 14690 10498 14702
rect 10894 14754 10946 14766
rect 10894 14690 10946 14702
rect 14142 14754 14194 14766
rect 20626 14702 20638 14754
rect 20690 14702 20702 14754
rect 14142 14690 14194 14702
rect 8542 14642 8594 14654
rect 8542 14578 8594 14590
rect 11678 14642 11730 14654
rect 11678 14578 11730 14590
rect 24222 14642 24274 14654
rect 24222 14578 24274 14590
rect 24558 14642 24610 14654
rect 24558 14578 24610 14590
rect 29150 14642 29202 14654
rect 29150 14578 29202 14590
rect 8878 14530 8930 14542
rect 10670 14530 10722 14542
rect 10210 14478 10222 14530
rect 10274 14478 10286 14530
rect 8878 14466 8930 14478
rect 10670 14466 10722 14478
rect 12238 14530 12290 14542
rect 13694 14530 13746 14542
rect 12786 14478 12798 14530
rect 12850 14478 12862 14530
rect 13458 14478 13470 14530
rect 13522 14478 13534 14530
rect 12238 14466 12290 14478
rect 13694 14466 13746 14478
rect 13918 14530 13970 14542
rect 13918 14466 13970 14478
rect 14814 14530 14866 14542
rect 14814 14466 14866 14478
rect 14926 14530 14978 14542
rect 14926 14466 14978 14478
rect 15150 14530 15202 14542
rect 15150 14466 15202 14478
rect 15598 14530 15650 14542
rect 19630 14530 19682 14542
rect 20526 14530 20578 14542
rect 18498 14478 18510 14530
rect 18562 14478 18574 14530
rect 19170 14478 19182 14530
rect 19234 14478 19246 14530
rect 20178 14478 20190 14530
rect 20242 14478 20254 14530
rect 15598 14466 15650 14478
rect 19630 14466 19682 14478
rect 20526 14466 20578 14478
rect 21310 14530 21362 14542
rect 21310 14466 21362 14478
rect 22878 14530 22930 14542
rect 22878 14466 22930 14478
rect 23102 14530 23154 14542
rect 24782 14530 24834 14542
rect 29374 14530 29426 14542
rect 23426 14478 23438 14530
rect 23490 14478 23502 14530
rect 25666 14478 25678 14530
rect 25730 14478 25742 14530
rect 27010 14478 27022 14530
rect 27074 14478 27086 14530
rect 23102 14466 23154 14478
rect 24782 14466 24834 14478
rect 29374 14466 29426 14478
rect 2046 14418 2098 14430
rect 2046 14354 2098 14366
rect 9214 14418 9266 14430
rect 9214 14354 9266 14366
rect 9886 14418 9938 14430
rect 9886 14354 9938 14366
rect 11902 14418 11954 14430
rect 11902 14354 11954 14366
rect 15262 14418 15314 14430
rect 15262 14354 15314 14366
rect 15710 14418 15762 14430
rect 15710 14354 15762 14366
rect 16718 14418 16770 14430
rect 16718 14354 16770 14366
rect 17054 14418 17106 14430
rect 17054 14354 17106 14366
rect 17726 14418 17778 14430
rect 17726 14354 17778 14366
rect 17950 14418 18002 14430
rect 17950 14354 18002 14366
rect 18062 14418 18114 14430
rect 23214 14418 23266 14430
rect 18722 14366 18734 14418
rect 18786 14366 18798 14418
rect 18062 14354 18114 14366
rect 23214 14354 23266 14366
rect 25454 14418 25506 14430
rect 25454 14354 25506 14366
rect 28254 14418 28306 14430
rect 28254 14354 28306 14366
rect 28590 14418 28642 14430
rect 30046 14418 30098 14430
rect 29698 14366 29710 14418
rect 29762 14366 29774 14418
rect 28590 14354 28642 14366
rect 30046 14354 30098 14366
rect 37886 14418 37938 14430
rect 37886 14354 37938 14366
rect 1710 14306 1762 14318
rect 1710 14242 1762 14254
rect 9550 14306 9602 14318
rect 9550 14242 9602 14254
rect 10334 14306 10386 14318
rect 10334 14242 10386 14254
rect 12574 14306 12626 14318
rect 12574 14242 12626 14254
rect 13582 14306 13634 14318
rect 16382 14306 16434 14318
rect 16034 14254 16046 14306
rect 16098 14254 16110 14306
rect 13582 14242 13634 14254
rect 16382 14242 16434 14254
rect 17502 14306 17554 14318
rect 17502 14242 17554 14254
rect 21870 14306 21922 14318
rect 21870 14242 21922 14254
rect 23886 14306 23938 14318
rect 27246 14306 27298 14318
rect 25106 14254 25118 14306
rect 25170 14254 25182 14306
rect 23886 14242 23938 14254
rect 27246 14242 27298 14254
rect 30382 14306 30434 14318
rect 30382 14242 30434 14254
rect 38222 14306 38274 14318
rect 38222 14242 38274 14254
rect 1344 14138 38800 14172
rect 1344 14086 10538 14138
rect 10590 14086 10642 14138
rect 10694 14086 10746 14138
rect 10798 14086 19862 14138
rect 19914 14086 19966 14138
rect 20018 14086 20070 14138
rect 20122 14086 29186 14138
rect 29238 14086 29290 14138
rect 29342 14086 29394 14138
rect 29446 14086 38510 14138
rect 38562 14086 38614 14138
rect 38666 14086 38718 14138
rect 38770 14086 38800 14138
rect 1344 14052 38800 14086
rect 13246 13970 13298 13982
rect 13246 13906 13298 13918
rect 18846 13970 18898 13982
rect 18846 13906 18898 13918
rect 19518 13970 19570 13982
rect 19518 13906 19570 13918
rect 22318 13970 22370 13982
rect 22318 13906 22370 13918
rect 1710 13858 1762 13870
rect 1710 13794 1762 13806
rect 2046 13858 2098 13870
rect 2046 13794 2098 13806
rect 11454 13858 11506 13870
rect 11454 13794 11506 13806
rect 12686 13858 12738 13870
rect 12686 13794 12738 13806
rect 14590 13858 14642 13870
rect 14590 13794 14642 13806
rect 14926 13858 14978 13870
rect 14926 13794 14978 13806
rect 16830 13858 16882 13870
rect 19630 13858 19682 13870
rect 17714 13806 17726 13858
rect 17778 13806 17790 13858
rect 16830 13794 16882 13806
rect 19630 13794 19682 13806
rect 20526 13858 20578 13870
rect 20526 13794 20578 13806
rect 23214 13858 23266 13870
rect 23214 13794 23266 13806
rect 24110 13858 24162 13870
rect 24110 13794 24162 13806
rect 24446 13858 24498 13870
rect 24446 13794 24498 13806
rect 25566 13858 25618 13870
rect 25566 13794 25618 13806
rect 26798 13858 26850 13870
rect 26798 13794 26850 13806
rect 27918 13858 27970 13870
rect 27918 13794 27970 13806
rect 29038 13858 29090 13870
rect 29038 13794 29090 13806
rect 38222 13858 38274 13870
rect 38222 13794 38274 13806
rect 10558 13746 10610 13758
rect 10322 13694 10334 13746
rect 10386 13694 10398 13746
rect 10558 13682 10610 13694
rect 11006 13746 11058 13758
rect 16158 13746 16210 13758
rect 17614 13746 17666 13758
rect 11666 13694 11678 13746
rect 11730 13694 11742 13746
rect 12450 13694 12462 13746
rect 12514 13694 12526 13746
rect 16594 13694 16606 13746
rect 16658 13694 16670 13746
rect 11006 13682 11058 13694
rect 16158 13682 16210 13694
rect 17614 13682 17666 13694
rect 17950 13746 18002 13758
rect 20078 13746 20130 13758
rect 18162 13694 18174 13746
rect 18226 13694 18238 13746
rect 19058 13694 19070 13746
rect 19122 13694 19134 13746
rect 17950 13682 18002 13694
rect 20078 13682 20130 13694
rect 21758 13746 21810 13758
rect 21758 13682 21810 13694
rect 23102 13746 23154 13758
rect 25230 13746 25282 13758
rect 23538 13694 23550 13746
rect 23602 13694 23614 13746
rect 23102 13682 23154 13694
rect 25230 13682 25282 13694
rect 26574 13746 26626 13758
rect 26574 13682 26626 13694
rect 26686 13746 26738 13758
rect 27806 13746 27858 13758
rect 28702 13746 28754 13758
rect 27570 13694 27582 13746
rect 27634 13694 27646 13746
rect 28354 13694 28366 13746
rect 28418 13694 28430 13746
rect 26686 13682 26738 13694
rect 27806 13682 27858 13694
rect 28702 13682 28754 13694
rect 37886 13746 37938 13758
rect 37886 13682 37938 13694
rect 14366 13634 14418 13646
rect 14366 13570 14418 13582
rect 15710 13634 15762 13646
rect 15710 13570 15762 13582
rect 18622 13634 18674 13646
rect 18622 13570 18674 13582
rect 22878 13634 22930 13646
rect 22878 13570 22930 13582
rect 10782 13522 10834 13534
rect 10782 13458 10834 13470
rect 11118 13522 11170 13534
rect 11118 13458 11170 13470
rect 15598 13522 15650 13534
rect 15598 13458 15650 13470
rect 23886 13522 23938 13534
rect 27234 13470 27246 13522
rect 27298 13470 27310 13522
rect 23886 13458 23938 13470
rect 1344 13354 38640 13388
rect 1344 13302 5876 13354
rect 5928 13302 5980 13354
rect 6032 13302 6084 13354
rect 6136 13302 15200 13354
rect 15252 13302 15304 13354
rect 15356 13302 15408 13354
rect 15460 13302 24524 13354
rect 24576 13302 24628 13354
rect 24680 13302 24732 13354
rect 24784 13302 33848 13354
rect 33900 13302 33952 13354
rect 34004 13302 34056 13354
rect 34108 13302 38640 13354
rect 1344 13268 38640 13302
rect 10222 13186 10274 13198
rect 10222 13122 10274 13134
rect 10334 13186 10386 13198
rect 10334 13122 10386 13134
rect 10782 13186 10834 13198
rect 13694 13186 13746 13198
rect 11106 13134 11118 13186
rect 11170 13183 11182 13186
rect 11442 13183 11454 13186
rect 11170 13137 11454 13183
rect 11170 13134 11182 13137
rect 11442 13134 11454 13137
rect 11506 13134 11518 13186
rect 10782 13122 10834 13134
rect 13694 13122 13746 13134
rect 14142 13186 14194 13198
rect 14142 13122 14194 13134
rect 15262 13186 15314 13198
rect 15262 13122 15314 13134
rect 16158 13186 16210 13198
rect 16158 13122 16210 13134
rect 24782 13186 24834 13198
rect 25106 13134 25118 13186
rect 25170 13134 25182 13186
rect 24782 13122 24834 13134
rect 11454 13074 11506 13086
rect 11454 13010 11506 13022
rect 16046 13074 16098 13086
rect 16046 13010 16098 13022
rect 17502 13074 17554 13086
rect 17502 13010 17554 13022
rect 21422 13074 21474 13086
rect 21422 13010 21474 13022
rect 2046 12962 2098 12974
rect 2046 12898 2098 12910
rect 2718 12962 2770 12974
rect 2718 12898 2770 12910
rect 10558 12962 10610 12974
rect 13918 12962 13970 12974
rect 12786 12910 12798 12962
rect 12850 12910 12862 12962
rect 13458 12910 13470 12962
rect 13522 12910 13534 12962
rect 10558 12898 10610 12910
rect 13918 12898 13970 12910
rect 14926 12962 14978 12974
rect 14926 12898 14978 12910
rect 15150 12962 15202 12974
rect 15150 12898 15202 12910
rect 15822 12962 15874 12974
rect 17726 12962 17778 12974
rect 18510 12962 18562 12974
rect 20414 12962 20466 12974
rect 17042 12910 17054 12962
rect 17106 12910 17118 12962
rect 18050 12910 18062 12962
rect 18114 12910 18126 12962
rect 19058 12910 19070 12962
rect 19122 12910 19134 12962
rect 15822 12898 15874 12910
rect 17726 12898 17778 12910
rect 18510 12898 18562 12910
rect 20414 12898 20466 12910
rect 21982 12962 22034 12974
rect 21982 12898 22034 12910
rect 22094 12962 22146 12974
rect 22094 12898 22146 12910
rect 22206 12962 22258 12974
rect 22206 12898 22258 12910
rect 22654 12962 22706 12974
rect 24558 12962 24610 12974
rect 23874 12910 23886 12962
rect 23938 12910 23950 12962
rect 22654 12898 22706 12910
rect 24558 12898 24610 12910
rect 25454 12962 25506 12974
rect 25454 12898 25506 12910
rect 27470 12962 27522 12974
rect 27470 12898 27522 12910
rect 37886 12962 37938 12974
rect 37886 12898 37938 12910
rect 1710 12850 1762 12862
rect 1710 12786 1762 12798
rect 10894 12850 10946 12862
rect 10894 12786 10946 12798
rect 14814 12850 14866 12862
rect 14814 12786 14866 12798
rect 15710 12850 15762 12862
rect 15710 12786 15762 12798
rect 16830 12850 16882 12862
rect 20750 12850 20802 12862
rect 17938 12798 17950 12850
rect 18002 12798 18014 12850
rect 16830 12786 16882 12798
rect 20750 12786 20802 12798
rect 22878 12850 22930 12862
rect 22878 12786 22930 12798
rect 23102 12850 23154 12862
rect 23102 12786 23154 12798
rect 25790 12850 25842 12862
rect 25790 12786 25842 12798
rect 26462 12850 26514 12862
rect 26462 12786 26514 12798
rect 26798 12850 26850 12862
rect 26798 12786 26850 12798
rect 37214 12850 37266 12862
rect 37214 12786 37266 12798
rect 38222 12850 38274 12862
rect 38222 12786 38274 12798
rect 2382 12738 2434 12750
rect 2382 12674 2434 12686
rect 12574 12738 12626 12750
rect 12574 12674 12626 12686
rect 13582 12738 13634 12750
rect 13582 12674 13634 12686
rect 18846 12738 18898 12750
rect 20078 12738 20130 12750
rect 19730 12686 19742 12738
rect 19794 12686 19806 12738
rect 18846 12674 18898 12686
rect 20078 12674 20130 12686
rect 23438 12738 23490 12750
rect 23438 12674 23490 12686
rect 24110 12738 24162 12750
rect 24110 12674 24162 12686
rect 26126 12738 26178 12750
rect 26126 12674 26178 12686
rect 27134 12738 27186 12750
rect 27134 12674 27186 12686
rect 27806 12738 27858 12750
rect 27806 12674 27858 12686
rect 37550 12738 37602 12750
rect 37550 12674 37602 12686
rect 1344 12570 38800 12604
rect 1344 12518 10538 12570
rect 10590 12518 10642 12570
rect 10694 12518 10746 12570
rect 10798 12518 19862 12570
rect 19914 12518 19966 12570
rect 20018 12518 20070 12570
rect 20122 12518 29186 12570
rect 29238 12518 29290 12570
rect 29342 12518 29394 12570
rect 29446 12518 38510 12570
rect 38562 12518 38614 12570
rect 38666 12518 38718 12570
rect 38770 12518 38800 12570
rect 1344 12484 38800 12518
rect 10670 12402 10722 12414
rect 10670 12338 10722 12350
rect 16270 12402 16322 12414
rect 16270 12338 16322 12350
rect 17502 12402 17554 12414
rect 25778 12350 25790 12402
rect 25842 12350 25854 12402
rect 17502 12338 17554 12350
rect 1710 12290 1762 12302
rect 1710 12226 1762 12238
rect 2046 12290 2098 12302
rect 2046 12226 2098 12238
rect 13806 12290 13858 12302
rect 27358 12290 27410 12302
rect 24546 12238 24558 12290
rect 24610 12238 24622 12290
rect 13806 12226 13858 12238
rect 27358 12226 27410 12238
rect 29038 12290 29090 12302
rect 29038 12226 29090 12238
rect 37886 12290 37938 12302
rect 37886 12226 37938 12238
rect 38222 12290 38274 12302
rect 38222 12226 38274 12238
rect 10222 12178 10274 12190
rect 10222 12114 10274 12126
rect 10334 12178 10386 12190
rect 10334 12114 10386 12126
rect 11790 12178 11842 12190
rect 11790 12114 11842 12126
rect 12238 12178 12290 12190
rect 12910 12178 12962 12190
rect 12674 12126 12686 12178
rect 12738 12126 12750 12178
rect 12238 12114 12290 12126
rect 12910 12114 12962 12126
rect 13134 12178 13186 12190
rect 13134 12114 13186 12126
rect 13358 12178 13410 12190
rect 13358 12114 13410 12126
rect 13470 12178 13522 12190
rect 24222 12178 24274 12190
rect 14018 12126 14030 12178
rect 14082 12126 14094 12178
rect 15474 12126 15486 12178
rect 15538 12126 15550 12178
rect 23426 12126 23438 12178
rect 23490 12126 23502 12178
rect 13470 12114 13522 12126
rect 24222 12114 24274 12126
rect 25230 12178 25282 12190
rect 25230 12114 25282 12126
rect 25454 12178 25506 12190
rect 25454 12114 25506 12126
rect 26126 12178 26178 12190
rect 26126 12114 26178 12126
rect 27022 12178 27074 12190
rect 27022 12114 27074 12126
rect 27806 12178 27858 12190
rect 27806 12114 27858 12126
rect 28030 12178 28082 12190
rect 28702 12178 28754 12190
rect 28354 12126 28366 12178
rect 28418 12126 28430 12178
rect 28030 12114 28082 12126
rect 28702 12114 28754 12126
rect 10558 12066 10610 12078
rect 10558 12002 10610 12014
rect 12014 12066 12066 12078
rect 12014 12002 12066 12014
rect 15262 12066 15314 12078
rect 15262 12002 15314 12014
rect 15822 12066 15874 12078
rect 15822 12002 15874 12014
rect 15934 12066 15986 12078
rect 15934 12002 15986 12014
rect 16382 12066 16434 12078
rect 26350 12066 26402 12078
rect 21298 12014 21310 12066
rect 21362 12014 21374 12066
rect 26674 12014 26686 12066
rect 26738 12014 26750 12066
rect 16382 12002 16434 12014
rect 26350 12002 26402 12014
rect 10782 11954 10834 11966
rect 10782 11890 10834 11902
rect 11678 11954 11730 11966
rect 11678 11890 11730 11902
rect 12350 11954 12402 11966
rect 12350 11890 12402 11902
rect 14926 11954 14978 11966
rect 14926 11890 14978 11902
rect 15038 11954 15090 11966
rect 15038 11890 15090 11902
rect 1344 11786 38640 11820
rect 1344 11734 5876 11786
rect 5928 11734 5980 11786
rect 6032 11734 6084 11786
rect 6136 11734 15200 11786
rect 15252 11734 15304 11786
rect 15356 11734 15408 11786
rect 15460 11734 24524 11786
rect 24576 11734 24628 11786
rect 24680 11734 24732 11786
rect 24784 11734 33848 11786
rect 33900 11734 33952 11786
rect 34004 11734 34056 11786
rect 34108 11734 38640 11786
rect 1344 11700 38640 11734
rect 27806 11618 27858 11630
rect 27806 11554 27858 11566
rect 25678 11506 25730 11518
rect 24210 11454 24222 11506
rect 24274 11454 24286 11506
rect 25678 11442 25730 11454
rect 26238 11506 26290 11518
rect 26238 11442 26290 11454
rect 26686 11506 26738 11518
rect 26686 11442 26738 11454
rect 26910 11506 26962 11518
rect 26910 11442 26962 11454
rect 27582 11506 27634 11518
rect 27582 11442 27634 11454
rect 2046 11394 2098 11406
rect 2046 11330 2098 11342
rect 10670 11394 10722 11406
rect 10670 11330 10722 11342
rect 11342 11394 11394 11406
rect 16046 11394 16098 11406
rect 13682 11342 13694 11394
rect 13746 11342 13758 11394
rect 11342 11330 11394 11342
rect 16046 11330 16098 11342
rect 16718 11394 16770 11406
rect 16718 11330 16770 11342
rect 17278 11394 17330 11406
rect 17714 11342 17726 11394
rect 17778 11342 17790 11394
rect 21298 11342 21310 11394
rect 21362 11342 21374 11394
rect 22082 11342 22094 11394
rect 22146 11342 22158 11394
rect 25554 11342 25566 11394
rect 25618 11342 25630 11394
rect 37986 11342 37998 11394
rect 38050 11342 38062 11394
rect 17278 11330 17330 11342
rect 16158 11282 16210 11294
rect 17390 11282 17442 11294
rect 18398 11282 18450 11294
rect 16370 11230 16382 11282
rect 16434 11230 16446 11282
rect 17602 11230 17614 11282
rect 17666 11230 17678 11282
rect 16158 11218 16210 11230
rect 17390 11218 17442 11230
rect 18398 11218 18450 11230
rect 19070 11282 19122 11294
rect 19070 11218 19122 11230
rect 19406 11282 19458 11294
rect 19406 11218 19458 11230
rect 19742 11282 19794 11294
rect 19742 11218 19794 11230
rect 20078 11282 20130 11294
rect 20078 11218 20130 11230
rect 20414 11282 20466 11294
rect 20414 11218 20466 11230
rect 20750 11282 20802 11294
rect 20750 11218 20802 11230
rect 24558 11282 24610 11294
rect 24558 11218 24610 11230
rect 25006 11282 25058 11294
rect 25006 11218 25058 11230
rect 25342 11282 25394 11294
rect 25342 11218 25394 11230
rect 25790 11282 25842 11294
rect 29150 11282 29202 11294
rect 28130 11230 28142 11282
rect 28194 11230 28206 11282
rect 25790 11218 25842 11230
rect 29150 11218 29202 11230
rect 1710 11170 1762 11182
rect 1710 11106 1762 11118
rect 10334 11170 10386 11182
rect 10334 11106 10386 11118
rect 11006 11170 11058 11182
rect 11006 11106 11058 11118
rect 13470 11170 13522 11182
rect 13470 11106 13522 11118
rect 15038 11170 15090 11182
rect 15038 11106 15090 11118
rect 15486 11170 15538 11182
rect 15486 11106 15538 11118
rect 16942 11170 16994 11182
rect 16942 11106 16994 11118
rect 18174 11170 18226 11182
rect 18174 11106 18226 11118
rect 18734 11170 18786 11182
rect 18734 11106 18786 11118
rect 24782 11170 24834 11182
rect 24782 11106 24834 11118
rect 25118 11170 25170 11182
rect 25118 11106 25170 11118
rect 26126 11170 26178 11182
rect 29486 11170 29538 11182
rect 27234 11118 27246 11170
rect 27298 11118 27310 11170
rect 26126 11106 26178 11118
rect 29486 11106 29538 11118
rect 38222 11170 38274 11182
rect 38222 11106 38274 11118
rect 1344 11002 38800 11036
rect 1344 10950 10538 11002
rect 10590 10950 10642 11002
rect 10694 10950 10746 11002
rect 10798 10950 19862 11002
rect 19914 10950 19966 11002
rect 20018 10950 20070 11002
rect 20122 10950 29186 11002
rect 29238 10950 29290 11002
rect 29342 10950 29394 11002
rect 29446 10950 38510 11002
rect 38562 10950 38614 11002
rect 38666 10950 38718 11002
rect 38770 10950 38800 11002
rect 1344 10916 38800 10950
rect 1710 10722 1762 10734
rect 1710 10658 1762 10670
rect 2046 10722 2098 10734
rect 2046 10658 2098 10670
rect 18062 10722 18114 10734
rect 18062 10658 18114 10670
rect 18734 10722 18786 10734
rect 37886 10722 37938 10734
rect 21746 10670 21758 10722
rect 21810 10670 21822 10722
rect 18734 10658 18786 10670
rect 37886 10658 37938 10670
rect 38222 10722 38274 10734
rect 38222 10658 38274 10670
rect 18274 10558 18286 10610
rect 18338 10558 18350 10610
rect 18946 10558 18958 10610
rect 19010 10558 19022 10610
rect 24658 10558 24670 10610
rect 24722 10558 24734 10610
rect 25330 10558 25342 10610
rect 25394 10558 25406 10610
rect 27234 10446 27246 10498
rect 27298 10446 27310 10498
rect 1344 10218 38640 10252
rect 1344 10166 5876 10218
rect 5928 10166 5980 10218
rect 6032 10166 6084 10218
rect 6136 10166 15200 10218
rect 15252 10166 15304 10218
rect 15356 10166 15408 10218
rect 15460 10166 24524 10218
rect 24576 10166 24628 10218
rect 24680 10166 24732 10218
rect 24784 10166 33848 10218
rect 33900 10166 33952 10218
rect 34004 10166 34056 10218
rect 34108 10166 38640 10218
rect 1344 10132 38640 10166
rect 19406 9938 19458 9950
rect 19406 9874 19458 9886
rect 27582 9938 27634 9950
rect 27582 9874 27634 9886
rect 2046 9826 2098 9838
rect 27806 9826 27858 9838
rect 26786 9774 26798 9826
rect 26850 9774 26862 9826
rect 2046 9762 2098 9774
rect 27806 9762 27858 9774
rect 28030 9826 28082 9838
rect 37886 9826 37938 9838
rect 29138 9774 29150 9826
rect 29202 9774 29214 9826
rect 28030 9762 28082 9774
rect 37886 9762 37938 9774
rect 20526 9714 20578 9726
rect 20526 9650 20578 9662
rect 20638 9714 20690 9726
rect 24882 9662 24894 9714
rect 24946 9662 24958 9714
rect 31154 9662 31166 9714
rect 31218 9662 31230 9714
rect 20638 9650 20690 9662
rect 1710 9602 1762 9614
rect 1710 9538 1762 9550
rect 20862 9602 20914 9614
rect 20862 9538 20914 9550
rect 27246 9602 27298 9614
rect 27246 9538 27298 9550
rect 27470 9602 27522 9614
rect 27470 9538 27522 9550
rect 28366 9602 28418 9614
rect 28366 9538 28418 9550
rect 38222 9602 38274 9614
rect 38222 9538 38274 9550
rect 1344 9434 38800 9468
rect 1344 9382 10538 9434
rect 10590 9382 10642 9434
rect 10694 9382 10746 9434
rect 10798 9382 19862 9434
rect 19914 9382 19966 9434
rect 20018 9382 20070 9434
rect 20122 9382 29186 9434
rect 29238 9382 29290 9434
rect 29342 9382 29394 9434
rect 29446 9382 38510 9434
rect 38562 9382 38614 9434
rect 38666 9382 38718 9434
rect 38770 9382 38800 9434
rect 1344 9348 38800 9382
rect 24334 9266 24386 9278
rect 24334 9202 24386 9214
rect 1710 9154 1762 9166
rect 1710 9090 1762 9102
rect 2046 9154 2098 9166
rect 22878 9154 22930 9166
rect 19730 9102 19742 9154
rect 19794 9102 19806 9154
rect 2046 9090 2098 9102
rect 22878 9090 22930 9102
rect 23214 9154 23266 9166
rect 23214 9090 23266 9102
rect 23326 9154 23378 9166
rect 23326 9090 23378 9102
rect 24558 9154 24610 9166
rect 24558 9090 24610 9102
rect 38222 9154 38274 9166
rect 38222 9090 38274 9102
rect 22318 9042 22370 9054
rect 23998 9042 24050 9054
rect 18946 8990 18958 9042
rect 19010 8990 19022 9042
rect 22642 8990 22654 9042
rect 22706 8990 22718 9042
rect 23538 8990 23550 9042
rect 23602 8990 23614 9042
rect 22318 8978 22370 8990
rect 23998 8978 24050 8990
rect 24110 9042 24162 9054
rect 25218 8990 25230 9042
rect 25282 8990 25294 9042
rect 37986 8990 37998 9042
rect 38050 8990 38062 9042
rect 24110 8978 24162 8990
rect 24670 8930 24722 8942
rect 21858 8878 21870 8930
rect 21922 8878 21934 8930
rect 27234 8878 27246 8930
rect 27298 8878 27310 8930
rect 24670 8866 24722 8878
rect 22990 8818 23042 8830
rect 22990 8754 23042 8766
rect 1344 8650 38640 8684
rect 1344 8598 5876 8650
rect 5928 8598 5980 8650
rect 6032 8598 6084 8650
rect 6136 8598 15200 8650
rect 15252 8598 15304 8650
rect 15356 8598 15408 8650
rect 15460 8598 24524 8650
rect 24576 8598 24628 8650
rect 24680 8598 24732 8650
rect 24784 8598 33848 8650
rect 33900 8598 33952 8650
rect 34004 8598 34056 8650
rect 34108 8598 38640 8650
rect 1344 8564 38640 8598
rect 3166 8370 3218 8382
rect 22866 8318 22878 8370
rect 22930 8318 22942 8370
rect 3166 8306 3218 8318
rect 23886 8258 23938 8270
rect 2594 8206 2606 8258
rect 2658 8206 2670 8258
rect 23886 8194 23938 8206
rect 24222 8258 24274 8270
rect 24222 8194 24274 8206
rect 24446 8258 24498 8270
rect 24446 8194 24498 8206
rect 24782 8258 24834 8270
rect 24782 8194 24834 8206
rect 25230 8258 25282 8270
rect 25230 8194 25282 8206
rect 25454 8258 25506 8270
rect 25454 8194 25506 8206
rect 25790 8258 25842 8270
rect 25790 8194 25842 8206
rect 25902 8258 25954 8270
rect 25902 8194 25954 8206
rect 36430 8258 36482 8270
rect 36430 8194 36482 8206
rect 37214 8258 37266 8270
rect 37214 8194 37266 8206
rect 37886 8258 37938 8270
rect 37886 8194 37938 8206
rect 1710 8146 1762 8158
rect 1710 8082 1762 8094
rect 2046 8146 2098 8158
rect 2046 8082 2098 8094
rect 22094 8146 22146 8158
rect 22094 8082 22146 8094
rect 22430 8146 22482 8158
rect 22430 8082 22482 8094
rect 23102 8146 23154 8158
rect 23102 8082 23154 8094
rect 38222 8146 38274 8158
rect 38222 8082 38274 8094
rect 2382 8034 2434 8046
rect 2382 7970 2434 7982
rect 22878 8034 22930 8046
rect 22878 7970 22930 7982
rect 23998 8034 24050 8046
rect 23998 7970 24050 7982
rect 24558 8034 24610 8046
rect 24558 7970 24610 7982
rect 25006 8034 25058 8046
rect 25006 7970 25058 7982
rect 25566 8034 25618 8046
rect 25566 7970 25618 7982
rect 27134 8034 27186 8046
rect 27134 7970 27186 7982
rect 37550 8034 37602 8046
rect 37550 7970 37602 7982
rect 1344 7866 38800 7900
rect 1344 7814 10538 7866
rect 10590 7814 10642 7866
rect 10694 7814 10746 7866
rect 10798 7814 19862 7866
rect 19914 7814 19966 7866
rect 20018 7814 20070 7866
rect 20122 7814 29186 7866
rect 29238 7814 29290 7866
rect 29342 7814 29394 7866
rect 29446 7814 38510 7866
rect 38562 7814 38614 7866
rect 38666 7814 38718 7866
rect 38770 7814 38800 7866
rect 1344 7780 38800 7814
rect 22878 7698 22930 7710
rect 22878 7634 22930 7646
rect 23550 7698 23602 7710
rect 23550 7634 23602 7646
rect 24110 7698 24162 7710
rect 24110 7634 24162 7646
rect 23438 7586 23490 7598
rect 19618 7534 19630 7586
rect 19682 7534 19694 7586
rect 23438 7522 23490 7534
rect 24222 7586 24274 7598
rect 24222 7522 24274 7534
rect 24670 7586 24722 7598
rect 24670 7522 24722 7534
rect 37886 7586 37938 7598
rect 37886 7522 37938 7534
rect 38222 7586 38274 7598
rect 38222 7522 38274 7534
rect 22990 7474 23042 7486
rect 18946 7422 18958 7474
rect 19010 7422 19022 7474
rect 22990 7410 23042 7422
rect 2382 7362 2434 7374
rect 21746 7310 21758 7362
rect 21810 7310 21822 7362
rect 2382 7298 2434 7310
rect 24558 7250 24610 7262
rect 24558 7186 24610 7198
rect 1344 7082 38640 7116
rect 1344 7030 5876 7082
rect 5928 7030 5980 7082
rect 6032 7030 6084 7082
rect 6136 7030 15200 7082
rect 15252 7030 15304 7082
rect 15356 7030 15408 7082
rect 15460 7030 24524 7082
rect 24576 7030 24628 7082
rect 24680 7030 24732 7082
rect 24784 7030 33848 7082
rect 33900 7030 33952 7082
rect 34004 7030 34056 7082
rect 34108 7030 38640 7082
rect 1344 6996 38640 7030
rect 37550 6690 37602 6702
rect 37986 6638 37998 6690
rect 38050 6638 38062 6690
rect 37550 6626 37602 6638
rect 38222 6466 38274 6478
rect 38222 6402 38274 6414
rect 1344 6298 38800 6332
rect 1344 6246 10538 6298
rect 10590 6246 10642 6298
rect 10694 6246 10746 6298
rect 10798 6246 19862 6298
rect 19914 6246 19966 6298
rect 20018 6246 20070 6298
rect 20122 6246 29186 6298
rect 29238 6246 29290 6298
rect 29342 6246 29394 6298
rect 29446 6246 38510 6298
rect 38562 6246 38614 6298
rect 38666 6246 38718 6298
rect 38770 6246 38800 6298
rect 1344 6212 38800 6246
rect 37662 6130 37714 6142
rect 37662 6066 37714 6078
rect 37886 6018 37938 6030
rect 37886 5954 37938 5966
rect 38222 6018 38274 6030
rect 38222 5954 38274 5966
rect 1344 5514 38640 5548
rect 1344 5462 5876 5514
rect 5928 5462 5980 5514
rect 6032 5462 6084 5514
rect 6136 5462 15200 5514
rect 15252 5462 15304 5514
rect 15356 5462 15408 5514
rect 15460 5462 24524 5514
rect 24576 5462 24628 5514
rect 24680 5462 24732 5514
rect 24784 5462 33848 5514
rect 33900 5462 33952 5514
rect 34004 5462 34056 5514
rect 34108 5462 38640 5514
rect 1344 5428 38640 5462
rect 37550 5234 37602 5246
rect 37550 5170 37602 5182
rect 37986 5070 37998 5122
rect 38050 5070 38062 5122
rect 38222 4898 38274 4910
rect 38222 4834 38274 4846
rect 1344 4730 38800 4764
rect 1344 4678 10538 4730
rect 10590 4678 10642 4730
rect 10694 4678 10746 4730
rect 10798 4678 19862 4730
rect 19914 4678 19966 4730
rect 20018 4678 20070 4730
rect 20122 4678 29186 4730
rect 29238 4678 29290 4730
rect 29342 4678 29394 4730
rect 29446 4678 38510 4730
rect 38562 4678 38614 4730
rect 38666 4678 38718 4730
rect 38770 4678 38800 4730
rect 1344 4644 38800 4678
rect 6414 4562 6466 4574
rect 5954 4510 5966 4562
rect 6018 4510 6030 4562
rect 6414 4498 6466 4510
rect 7646 4562 7698 4574
rect 7646 4498 7698 4510
rect 9998 4562 10050 4574
rect 9998 4498 10050 4510
rect 33854 4562 33906 4574
rect 33854 4498 33906 4510
rect 37662 4562 37714 4574
rect 37662 4498 37714 4510
rect 16382 4450 16434 4462
rect 16382 4386 16434 4398
rect 16718 4450 16770 4462
rect 16718 4386 16770 4398
rect 27134 4450 27186 4462
rect 27134 4386 27186 4398
rect 37886 4450 37938 4462
rect 37886 4386 37938 4398
rect 38222 4450 38274 4462
rect 38222 4386 38274 4398
rect 5630 4338 5682 4350
rect 5630 4274 5682 4286
rect 9102 4338 9154 4350
rect 9102 4274 9154 4286
rect 9662 4338 9714 4350
rect 27346 4286 27358 4338
rect 27410 4286 27422 4338
rect 9662 4274 9714 4286
rect 5406 4226 5458 4238
rect 5406 4162 5458 4174
rect 6974 4226 7026 4238
rect 6974 4162 7026 4174
rect 8094 4226 8146 4238
rect 8094 4162 8146 4174
rect 8654 4226 8706 4238
rect 8654 4162 8706 4174
rect 10446 4226 10498 4238
rect 10446 4162 10498 4174
rect 15934 4226 15986 4238
rect 15934 4162 15986 4174
rect 20414 4226 20466 4238
rect 20414 4162 20466 4174
rect 21534 4226 21586 4238
rect 21534 4162 21586 4174
rect 22206 4226 22258 4238
rect 22206 4162 22258 4174
rect 34638 4226 34690 4238
rect 34638 4162 34690 4174
rect 1344 3946 38640 3980
rect 1344 3894 5876 3946
rect 5928 3894 5980 3946
rect 6032 3894 6084 3946
rect 6136 3894 15200 3946
rect 15252 3894 15304 3946
rect 15356 3894 15408 3946
rect 15460 3894 24524 3946
rect 24576 3894 24628 3946
rect 24680 3894 24732 3946
rect 24784 3894 33848 3946
rect 33900 3894 33952 3946
rect 34004 3894 34056 3946
rect 34108 3894 38640 3946
rect 1344 3860 38640 3894
rect 37550 3666 37602 3678
rect 37550 3602 37602 3614
rect 10222 3554 10274 3566
rect 5842 3502 5854 3554
rect 5906 3502 5918 3554
rect 7186 3502 7198 3554
rect 7250 3502 7262 3554
rect 7858 3502 7870 3554
rect 7922 3502 7934 3554
rect 8530 3502 8542 3554
rect 8594 3502 8606 3554
rect 10222 3490 10274 3502
rect 10894 3554 10946 3566
rect 10894 3490 10946 3502
rect 11566 3554 11618 3566
rect 13694 3554 13746 3566
rect 16046 3554 16098 3566
rect 18510 3554 18562 3566
rect 20190 3554 20242 3566
rect 24894 3554 24946 3566
rect 12338 3502 12350 3554
rect 12402 3502 12414 3554
rect 14914 3502 14926 3554
rect 14978 3502 14990 3554
rect 15474 3502 15486 3554
rect 15538 3502 15550 3554
rect 17266 3502 17278 3554
rect 17330 3502 17342 3554
rect 17938 3502 17950 3554
rect 18002 3502 18014 3554
rect 19282 3502 19294 3554
rect 19346 3502 19358 3554
rect 21298 3502 21310 3554
rect 21362 3502 21374 3554
rect 21970 3502 21982 3554
rect 22034 3502 22046 3554
rect 22642 3502 22654 3554
rect 22706 3502 22718 3554
rect 23314 3502 23326 3554
rect 23378 3502 23390 3554
rect 11566 3490 11618 3502
rect 13694 3490 13746 3502
rect 16046 3490 16098 3502
rect 18510 3490 18562 3502
rect 20190 3490 20242 3502
rect 24894 3490 24946 3502
rect 25566 3554 25618 3566
rect 29374 3554 29426 3566
rect 26114 3502 26126 3554
rect 26178 3502 26190 3554
rect 26786 3502 26798 3554
rect 26850 3502 26862 3554
rect 27458 3502 27470 3554
rect 27522 3502 27534 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 29922 3502 29934 3554
rect 29986 3502 29998 3554
rect 30594 3502 30606 3554
rect 30658 3502 30670 3554
rect 31266 3502 31278 3554
rect 31330 3502 31342 3554
rect 32386 3502 32398 3554
rect 32450 3502 32462 3554
rect 33730 3502 33742 3554
rect 33794 3502 33806 3554
rect 34402 3502 34414 3554
rect 34466 3502 34478 3554
rect 35074 3502 35086 3554
rect 35138 3502 35150 3554
rect 37986 3502 37998 3554
rect 38050 3502 38062 3554
rect 25566 3490 25618 3502
rect 29374 3490 29426 3502
rect 6414 3442 6466 3454
rect 8766 3442 8818 3454
rect 6738 3390 6750 3442
rect 6802 3390 6814 3442
rect 8082 3390 8094 3442
rect 8146 3390 8158 3442
rect 6414 3378 6466 3390
rect 8766 3378 8818 3390
rect 9550 3442 9602 3454
rect 13358 3442 13410 3454
rect 9874 3390 9886 3442
rect 9938 3390 9950 3442
rect 9550 3378 9602 3390
rect 13358 3378 13410 3390
rect 14366 3442 14418 3454
rect 14366 3378 14418 3390
rect 15710 3442 15762 3454
rect 15710 3378 15762 3390
rect 16382 3442 16434 3454
rect 16382 3378 16434 3390
rect 19854 3442 19906 3454
rect 19854 3378 19906 3390
rect 22430 3442 22482 3454
rect 22430 3378 22482 3390
rect 25230 3442 25282 3454
rect 29038 3442 29090 3454
rect 32846 3442 32898 3454
rect 25890 3390 25902 3442
rect 25954 3390 25966 3442
rect 27234 3390 27246 3442
rect 27298 3390 27310 3442
rect 30370 3390 30382 3442
rect 30434 3390 30446 3442
rect 32162 3390 32174 3442
rect 32226 3390 32238 3442
rect 25230 3378 25282 3390
rect 29038 3378 29090 3390
rect 32846 3378 32898 3390
rect 33182 3442 33234 3454
rect 38222 3442 38274 3454
rect 34178 3390 34190 3442
rect 34242 3390 34254 3442
rect 34850 3390 34862 3442
rect 34914 3390 34926 3442
rect 33182 3378 33234 3390
rect 38222 3378 38274 3390
rect 6078 3330 6130 3342
rect 6078 3266 6130 3278
rect 7422 3330 7474 3342
rect 7422 3266 7474 3278
rect 10558 3330 10610 3342
rect 10558 3266 10610 3278
rect 11230 3330 11282 3342
rect 11230 3266 11282 3278
rect 11902 3330 11954 3342
rect 11902 3266 11954 3278
rect 12574 3330 12626 3342
rect 12574 3266 12626 3278
rect 14030 3330 14082 3342
rect 14030 3266 14082 3278
rect 14702 3330 14754 3342
rect 14702 3266 14754 3278
rect 17502 3330 17554 3342
rect 17502 3266 17554 3278
rect 18174 3330 18226 3342
rect 18174 3266 18226 3278
rect 18846 3330 18898 3342
rect 18846 3266 18898 3278
rect 19518 3330 19570 3342
rect 19518 3266 19570 3278
rect 21086 3330 21138 3342
rect 21086 3266 21138 3278
rect 21758 3330 21810 3342
rect 24558 3330 24610 3342
rect 23090 3278 23102 3330
rect 23154 3278 23166 3330
rect 21758 3266 21810 3278
rect 24558 3266 24610 3278
rect 26574 3330 26626 3342
rect 26574 3266 26626 3278
rect 28366 3330 28418 3342
rect 31054 3330 31106 3342
rect 29698 3278 29710 3330
rect 29762 3278 29774 3330
rect 33506 3278 33518 3330
rect 33570 3278 33582 3330
rect 28366 3266 28418 3278
rect 31054 3266 31106 3278
rect 1344 3162 38800 3196
rect 1344 3110 10538 3162
rect 10590 3110 10642 3162
rect 10694 3110 10746 3162
rect 10798 3110 19862 3162
rect 19914 3110 19966 3162
rect 20018 3110 20070 3162
rect 20122 3110 29186 3162
rect 29238 3110 29290 3162
rect 29342 3110 29394 3162
rect 29446 3110 38510 3162
rect 38562 3110 38614 3162
rect 38666 3110 38718 3162
rect 38770 3110 38800 3162
rect 1344 3076 38800 3110
rect 33618 2494 33630 2546
rect 33682 2543 33694 2546
rect 34626 2543 34638 2546
rect 33682 2497 34638 2543
rect 33682 2494 33694 2497
rect 34626 2494 34638 2497
rect 34690 2543 34702 2546
rect 35074 2543 35086 2546
rect 34690 2497 35086 2543
rect 34690 2494 34702 2497
rect 35074 2494 35086 2497
rect 35138 2494 35150 2546
rect 30258 926 30270 978
rect 30322 975 30334 978
rect 31042 975 31054 978
rect 30322 929 31054 975
rect 30322 926 30334 929
rect 31042 926 31054 929
rect 31106 926 31118 978
<< via1 >>
rect 32286 37774 32338 37826
rect 33518 37774 33570 37826
rect 33630 37662 33682 37714
rect 34862 37662 34914 37714
rect 5876 36822 5928 36874
rect 5980 36822 6032 36874
rect 6084 36822 6136 36874
rect 15200 36822 15252 36874
rect 15304 36822 15356 36874
rect 15408 36822 15460 36874
rect 24524 36822 24576 36874
rect 24628 36822 24680 36874
rect 24732 36822 24784 36874
rect 33848 36822 33900 36874
rect 33952 36822 34004 36874
rect 34056 36822 34108 36874
rect 2718 36430 2770 36482
rect 4062 36430 4114 36482
rect 4846 36430 4898 36482
rect 5742 36430 5794 36482
rect 6526 36430 6578 36482
rect 7870 36430 7922 36482
rect 9662 36430 9714 36482
rect 10334 36430 10386 36482
rect 11006 36430 11058 36482
rect 11678 36430 11730 36482
rect 14814 36430 14866 36482
rect 15486 36430 15538 36482
rect 17278 36430 17330 36482
rect 17950 36430 18002 36482
rect 19294 36430 19346 36482
rect 22654 36430 22706 36482
rect 23326 36430 23378 36482
rect 25454 36430 25506 36482
rect 26798 36430 26850 36482
rect 27470 36430 27522 36482
rect 29262 36430 29314 36482
rect 32398 36430 32450 36482
rect 33070 36430 33122 36482
rect 34414 36430 34466 36482
rect 36206 36430 36258 36482
rect 36878 36430 36930 36482
rect 37550 36430 37602 36482
rect 3278 36318 3330 36370
rect 3614 36318 3666 36370
rect 4622 36318 4674 36370
rect 7086 36318 7138 36370
rect 7422 36318 7474 36370
rect 8094 36318 8146 36370
rect 8430 36318 8482 36370
rect 8766 36318 8818 36370
rect 9886 36318 9938 36370
rect 10558 36318 10610 36370
rect 11230 36318 11282 36370
rect 11902 36318 11954 36370
rect 12238 36318 12290 36370
rect 12574 36318 12626 36370
rect 13358 36318 13410 36370
rect 13694 36318 13746 36370
rect 14030 36318 14082 36370
rect 14366 36318 14418 36370
rect 16046 36318 16098 36370
rect 16382 36318 16434 36370
rect 17502 36318 17554 36370
rect 18174 36318 18226 36370
rect 18510 36318 18562 36370
rect 18846 36318 18898 36370
rect 19518 36318 19570 36370
rect 19854 36318 19906 36370
rect 20190 36318 20242 36370
rect 21086 36318 21138 36370
rect 21422 36318 21474 36370
rect 21758 36318 21810 36370
rect 22094 36318 22146 36370
rect 22430 36318 22482 36370
rect 23102 36318 23154 36370
rect 24558 36318 24610 36370
rect 24894 36318 24946 36370
rect 25230 36318 25282 36370
rect 25902 36318 25954 36370
rect 26238 36318 26290 36370
rect 26574 36318 26626 36370
rect 27246 36318 27298 36370
rect 28366 36318 28418 36370
rect 28702 36318 28754 36370
rect 29710 36318 29762 36370
rect 30046 36318 30098 36370
rect 30718 36318 30770 36370
rect 31054 36318 31106 36370
rect 31390 36318 31442 36370
rect 32174 36318 32226 36370
rect 32846 36318 32898 36370
rect 33518 36318 33570 36370
rect 33854 36318 33906 36370
rect 34190 36318 34242 36370
rect 34862 36318 34914 36370
rect 35198 36318 35250 36370
rect 35982 36318 36034 36370
rect 36654 36318 36706 36370
rect 37326 36318 37378 36370
rect 2942 36206 2994 36258
rect 4286 36206 4338 36258
rect 6078 36206 6130 36258
rect 6750 36206 6802 36258
rect 15038 36206 15090 36258
rect 15710 36206 15762 36258
rect 29038 36206 29090 36258
rect 30382 36206 30434 36258
rect 38110 36206 38162 36258
rect 10538 36038 10590 36090
rect 10642 36038 10694 36090
rect 10746 36038 10798 36090
rect 19862 36038 19914 36090
rect 19966 36038 20018 36090
rect 20070 36038 20122 36090
rect 29186 36038 29238 36090
rect 29290 36038 29342 36090
rect 29394 36038 29446 36090
rect 38510 36038 38562 36090
rect 38614 36038 38666 36090
rect 38718 36038 38770 36090
rect 3166 35870 3218 35922
rect 4510 35870 4562 35922
rect 5406 35870 5458 35922
rect 5630 35870 5682 35922
rect 6974 35870 7026 35922
rect 9102 35870 9154 35922
rect 9662 35870 9714 35922
rect 15262 35870 15314 35922
rect 15934 35870 15986 35922
rect 16382 35870 16434 35922
rect 27134 35870 27186 35922
rect 33742 35870 33794 35922
rect 34526 35870 34578 35922
rect 5966 35758 6018 35810
rect 9998 35758 10050 35810
rect 37550 35758 37602 35810
rect 38222 35758 38274 35810
rect 16606 35646 16658 35698
rect 27358 35646 27410 35698
rect 34750 35646 34802 35698
rect 37214 35646 37266 35698
rect 37886 35646 37938 35698
rect 3614 35534 3666 35586
rect 4174 35534 4226 35586
rect 6414 35534 6466 35586
rect 10446 35534 10498 35586
rect 32510 35534 32562 35586
rect 33182 35534 33234 35586
rect 34190 35534 34242 35586
rect 35310 35534 35362 35586
rect 35758 35534 35810 35586
rect 36318 35534 36370 35586
rect 36878 35534 36930 35586
rect 4174 35422 4226 35474
rect 4622 35422 4674 35474
rect 5876 35254 5928 35306
rect 5980 35254 6032 35306
rect 6084 35254 6136 35306
rect 15200 35254 15252 35306
rect 15304 35254 15356 35306
rect 15408 35254 15460 35306
rect 24524 35254 24576 35306
rect 24628 35254 24680 35306
rect 24732 35254 24784 35306
rect 33848 35254 33900 35306
rect 33952 35254 34004 35306
rect 34056 35254 34108 35306
rect 37662 34750 37714 34802
rect 37886 34750 37938 34802
rect 37102 34638 37154 34690
rect 38222 34638 38274 34690
rect 10538 34470 10590 34522
rect 10642 34470 10694 34522
rect 10746 34470 10798 34522
rect 19862 34470 19914 34522
rect 19966 34470 20018 34522
rect 20070 34470 20122 34522
rect 29186 34470 29238 34522
rect 29290 34470 29342 34522
rect 29394 34470 29446 34522
rect 38510 34470 38562 34522
rect 38614 34470 38666 34522
rect 38718 34470 38770 34522
rect 38222 34190 38274 34242
rect 37998 34078 38050 34130
rect 37550 33966 37602 34018
rect 5876 33686 5928 33738
rect 5980 33686 6032 33738
rect 6084 33686 6136 33738
rect 15200 33686 15252 33738
rect 15304 33686 15356 33738
rect 15408 33686 15460 33738
rect 24524 33686 24576 33738
rect 24628 33686 24680 33738
rect 24732 33686 24784 33738
rect 33848 33686 33900 33738
rect 33952 33686 34004 33738
rect 34056 33686 34108 33738
rect 37886 33182 37938 33234
rect 1710 33070 1762 33122
rect 2046 33070 2098 33122
rect 2494 33070 2546 33122
rect 37662 33070 37714 33122
rect 38222 33070 38274 33122
rect 10538 32902 10590 32954
rect 10642 32902 10694 32954
rect 10746 32902 10798 32954
rect 19862 32902 19914 32954
rect 19966 32902 20018 32954
rect 20070 32902 20122 32954
rect 29186 32902 29238 32954
rect 29290 32902 29342 32954
rect 29394 32902 29446 32954
rect 38510 32902 38562 32954
rect 38614 32902 38666 32954
rect 38718 32902 38770 32954
rect 1710 32622 1762 32674
rect 38222 32622 38274 32674
rect 2046 32510 2098 32562
rect 37550 32510 37602 32562
rect 37998 32510 38050 32562
rect 2606 32398 2658 32450
rect 2942 32398 2994 32450
rect 2270 32286 2322 32338
rect 2942 32286 2994 32338
rect 5876 32118 5928 32170
rect 5980 32118 6032 32170
rect 6084 32118 6136 32170
rect 15200 32118 15252 32170
rect 15304 32118 15356 32170
rect 15408 32118 15460 32170
rect 24524 32118 24576 32170
rect 24628 32118 24680 32170
rect 24732 32118 24784 32170
rect 33848 32118 33900 32170
rect 33952 32118 34004 32170
rect 34056 32118 34108 32170
rect 2046 31614 2098 31666
rect 2382 31614 2434 31666
rect 2718 31614 2770 31666
rect 37214 31614 37266 31666
rect 37550 31614 37602 31666
rect 37886 31614 37938 31666
rect 1710 31502 1762 31554
rect 3278 31502 3330 31554
rect 38222 31502 38274 31554
rect 10538 31334 10590 31386
rect 10642 31334 10694 31386
rect 10746 31334 10798 31386
rect 19862 31334 19914 31386
rect 19966 31334 20018 31386
rect 20070 31334 20122 31386
rect 29186 31334 29238 31386
rect 29290 31334 29342 31386
rect 29394 31334 29446 31386
rect 38510 31334 38562 31386
rect 38614 31334 38666 31386
rect 38718 31334 38770 31386
rect 1710 31054 1762 31106
rect 38222 31054 38274 31106
rect 1934 30942 1986 30994
rect 37886 30942 37938 30994
rect 2494 30830 2546 30882
rect 5876 30550 5928 30602
rect 5980 30550 6032 30602
rect 6084 30550 6136 30602
rect 15200 30550 15252 30602
rect 15304 30550 15356 30602
rect 15408 30550 15460 30602
rect 24524 30550 24576 30602
rect 24628 30550 24680 30602
rect 24732 30550 24784 30602
rect 33848 30550 33900 30602
rect 33952 30550 34004 30602
rect 34056 30550 34108 30602
rect 18958 30158 19010 30210
rect 21534 30158 21586 30210
rect 24110 30158 24162 30210
rect 25566 30158 25618 30210
rect 28030 30158 28082 30210
rect 2046 30046 2098 30098
rect 13694 30046 13746 30098
rect 14030 30046 14082 30098
rect 18734 30046 18786 30098
rect 21758 30046 21810 30098
rect 22094 30046 22146 30098
rect 22430 30046 22482 30098
rect 23326 30046 23378 30098
rect 23662 30046 23714 30098
rect 24334 30046 24386 30098
rect 25790 30046 25842 30098
rect 26126 30046 26178 30098
rect 26462 30046 26514 30098
rect 27246 30046 27298 30098
rect 27582 30046 27634 30098
rect 28254 30046 28306 30098
rect 37886 30046 37938 30098
rect 1710 29934 1762 29986
rect 2606 29934 2658 29986
rect 17390 29934 17442 29986
rect 18398 29934 18450 29986
rect 19630 29934 19682 29986
rect 38222 29934 38274 29986
rect 10538 29766 10590 29818
rect 10642 29766 10694 29818
rect 10746 29766 10798 29818
rect 19862 29766 19914 29818
rect 19966 29766 20018 29818
rect 20070 29766 20122 29818
rect 29186 29766 29238 29818
rect 29290 29766 29342 29818
rect 29394 29766 29446 29818
rect 38510 29766 38562 29818
rect 38614 29766 38666 29818
rect 38718 29766 38770 29818
rect 14366 29598 14418 29650
rect 18734 29598 18786 29650
rect 19630 29598 19682 29650
rect 21534 29598 21586 29650
rect 21870 29598 21922 29650
rect 23326 29598 23378 29650
rect 24222 29598 24274 29650
rect 25790 29598 25842 29650
rect 27134 29598 27186 29650
rect 28030 29598 28082 29650
rect 1710 29486 1762 29538
rect 14030 29486 14082 29538
rect 19294 29486 19346 29538
rect 19966 29486 20018 29538
rect 20302 29486 20354 29538
rect 38222 29486 38274 29538
rect 2046 29374 2098 29426
rect 13246 29374 13298 29426
rect 14590 29374 14642 29426
rect 15822 29374 15874 29426
rect 16718 29374 16770 29426
rect 17838 29374 17890 29426
rect 17950 29374 18002 29426
rect 18062 29374 18114 29426
rect 18286 29374 18338 29426
rect 22430 29374 22482 29426
rect 37886 29374 37938 29426
rect 2494 29262 2546 29314
rect 15374 29262 15426 29314
rect 16270 29262 16322 29314
rect 20974 29262 21026 29314
rect 22766 29262 22818 29314
rect 23662 29262 23714 29314
rect 25230 29262 25282 29314
rect 26574 29262 26626 29314
rect 27470 29262 27522 29314
rect 13470 29150 13522 29202
rect 13694 29150 13746 29202
rect 13918 29150 13970 29202
rect 16158 29150 16210 29202
rect 16606 29150 16658 29202
rect 21198 29150 21250 29202
rect 22206 29150 22258 29202
rect 22990 29150 23042 29202
rect 23886 29150 23938 29202
rect 25454 29150 25506 29202
rect 26798 29150 26850 29202
rect 27694 29150 27746 29202
rect 5876 28982 5928 29034
rect 5980 28982 6032 29034
rect 6084 28982 6136 29034
rect 15200 28982 15252 29034
rect 15304 28982 15356 29034
rect 15408 28982 15460 29034
rect 24524 28982 24576 29034
rect 24628 28982 24680 29034
rect 24732 28982 24784 29034
rect 33848 28982 33900 29034
rect 33952 28982 34004 29034
rect 34056 28982 34108 29034
rect 14254 28814 14306 28866
rect 15486 28814 15538 28866
rect 15822 28814 15874 28866
rect 18734 28814 18786 28866
rect 25230 28814 25282 28866
rect 25566 28814 25618 28866
rect 13918 28702 13970 28754
rect 16494 28702 16546 28754
rect 16942 28702 16994 28754
rect 17390 28702 17442 28754
rect 13582 28590 13634 28642
rect 13694 28590 13746 28642
rect 14142 28590 14194 28642
rect 15598 28590 15650 28642
rect 16046 28590 16098 28642
rect 17838 28590 17890 28642
rect 17950 28590 18002 28642
rect 18062 28590 18114 28642
rect 18398 28590 18450 28642
rect 19182 28590 19234 28642
rect 19854 28590 19906 28642
rect 21758 28590 21810 28642
rect 21870 28590 21922 28642
rect 22430 28590 22482 28642
rect 25006 28590 25058 28642
rect 26014 28590 26066 28642
rect 2046 28478 2098 28530
rect 11454 28478 11506 28530
rect 11790 28478 11842 28530
rect 22094 28478 22146 28530
rect 23774 28478 23826 28530
rect 24110 28478 24162 28530
rect 26238 28478 26290 28530
rect 27358 28478 27410 28530
rect 27694 28478 27746 28530
rect 37886 28478 37938 28530
rect 1710 28366 1762 28418
rect 18958 28366 19010 28418
rect 22654 28366 22706 28418
rect 38222 28366 38274 28418
rect 10538 28198 10590 28250
rect 10642 28198 10694 28250
rect 10746 28198 10798 28250
rect 19862 28198 19914 28250
rect 19966 28198 20018 28250
rect 20070 28198 20122 28250
rect 29186 28198 29238 28250
rect 29290 28198 29342 28250
rect 29394 28198 29446 28250
rect 38510 28198 38562 28250
rect 38614 28198 38666 28250
rect 38718 28198 38770 28250
rect 12350 28030 12402 28082
rect 19854 28030 19906 28082
rect 23550 28030 23602 28082
rect 24222 28030 24274 28082
rect 26014 28030 26066 28082
rect 28926 28030 28978 28082
rect 1710 27918 1762 27970
rect 14702 27918 14754 27970
rect 15598 27918 15650 27970
rect 18398 27918 18450 27970
rect 20190 27918 20242 27970
rect 20526 27918 20578 27970
rect 22094 27918 22146 27970
rect 22206 27918 22258 27970
rect 25454 27918 25506 27970
rect 26574 27918 26626 27970
rect 27694 27918 27746 27970
rect 38222 27918 38274 27970
rect 2046 27806 2098 27858
rect 12574 27806 12626 27858
rect 13134 27806 13186 27858
rect 14814 27806 14866 27858
rect 15262 27806 15314 27858
rect 15710 27806 15762 27858
rect 16046 27806 16098 27858
rect 18286 27806 18338 27858
rect 18622 27806 18674 27858
rect 19070 27806 19122 27858
rect 19518 27806 19570 27858
rect 21870 27806 21922 27858
rect 22430 27806 22482 27858
rect 22878 27806 22930 27858
rect 23214 27806 23266 27858
rect 23886 27806 23938 27858
rect 25342 27806 25394 27858
rect 25566 27806 25618 27858
rect 26462 27806 26514 27858
rect 26686 27806 26738 27858
rect 27470 27806 27522 27858
rect 27806 27806 27858 27858
rect 28254 27806 28306 27858
rect 28590 27806 28642 27858
rect 37998 27806 38050 27858
rect 12014 27694 12066 27746
rect 16942 27694 16994 27746
rect 17502 27694 17554 27746
rect 18062 27694 18114 27746
rect 37550 27694 37602 27746
rect 11342 27582 11394 27634
rect 11454 27582 11506 27634
rect 11678 27582 11730 27634
rect 11902 27582 11954 27634
rect 13358 27582 13410 27634
rect 13582 27582 13634 27634
rect 13806 27582 13858 27634
rect 13918 27582 13970 27634
rect 15038 27582 15090 27634
rect 15934 27582 15986 27634
rect 17390 27582 17442 27634
rect 27134 27582 27186 27634
rect 5876 27414 5928 27466
rect 5980 27414 6032 27466
rect 6084 27414 6136 27466
rect 15200 27414 15252 27466
rect 15304 27414 15356 27466
rect 15408 27414 15460 27466
rect 24524 27414 24576 27466
rect 24628 27414 24680 27466
rect 24732 27414 24784 27466
rect 33848 27414 33900 27466
rect 33952 27414 34004 27466
rect 34056 27414 34108 27466
rect 10446 27246 10498 27298
rect 10670 27246 10722 27298
rect 15934 27134 15986 27186
rect 20190 27134 20242 27186
rect 21758 27134 21810 27186
rect 10222 27022 10274 27074
rect 10894 27022 10946 27074
rect 11230 27022 11282 27074
rect 12350 27022 12402 27074
rect 13918 27022 13970 27074
rect 14926 27022 14978 27074
rect 15374 27022 15426 27074
rect 15710 27022 15762 27074
rect 16158 27022 16210 27074
rect 17390 27022 17442 27074
rect 17950 27022 18002 27074
rect 18174 27022 18226 27074
rect 18510 27022 18562 27074
rect 21982 27022 22034 27074
rect 22318 27022 22370 27074
rect 22990 27022 23042 27074
rect 24670 27022 24722 27074
rect 24894 27022 24946 27074
rect 25006 27022 25058 27074
rect 26910 27022 26962 27074
rect 37214 27022 37266 27074
rect 2046 26910 2098 26962
rect 2382 26910 2434 26962
rect 2718 26910 2770 26962
rect 9438 26910 9490 26962
rect 9774 26910 9826 26962
rect 10110 26910 10162 26962
rect 11342 26910 11394 26962
rect 12798 26910 12850 26962
rect 13582 26910 13634 26962
rect 15150 26910 15202 26962
rect 17614 26910 17666 26962
rect 18398 26910 18450 26962
rect 18958 26910 19010 26962
rect 19406 26910 19458 26962
rect 19742 26910 19794 26962
rect 22206 26910 22258 26962
rect 22766 26910 22818 26962
rect 23326 26910 23378 26962
rect 25454 26910 25506 26962
rect 25790 26910 25842 26962
rect 26126 26910 26178 26962
rect 27134 26910 27186 26962
rect 28254 26910 28306 26962
rect 28590 26910 28642 26962
rect 37550 26910 37602 26962
rect 37886 26910 37938 26962
rect 38222 26910 38274 26962
rect 1710 26798 1762 26850
rect 11902 26798 11954 26850
rect 10538 26630 10590 26682
rect 10642 26630 10694 26682
rect 10746 26630 10798 26682
rect 19862 26630 19914 26682
rect 19966 26630 20018 26682
rect 20070 26630 20122 26682
rect 29186 26630 29238 26682
rect 29290 26630 29342 26682
rect 29394 26630 29446 26682
rect 38510 26630 38562 26682
rect 38614 26630 38666 26682
rect 38718 26630 38770 26682
rect 10110 26462 10162 26514
rect 11678 26462 11730 26514
rect 13022 26462 13074 26514
rect 14478 26462 14530 26514
rect 15934 26462 15986 26514
rect 16606 26462 16658 26514
rect 17838 26462 17890 26514
rect 18174 26462 18226 26514
rect 21534 26462 21586 26514
rect 23438 26462 23490 26514
rect 26462 26462 26514 26514
rect 28142 26462 28194 26514
rect 1710 26350 1762 26402
rect 10446 26350 10498 26402
rect 15598 26350 15650 26402
rect 17502 26350 17554 26402
rect 19182 26350 19234 26402
rect 21982 26350 22034 26402
rect 24110 26350 24162 26402
rect 38222 26350 38274 26402
rect 2046 26238 2098 26290
rect 9774 26238 9826 26290
rect 10670 26238 10722 26290
rect 11118 26238 11170 26290
rect 11342 26238 11394 26290
rect 12686 26238 12738 26290
rect 13582 26238 13634 26290
rect 14142 26238 14194 26290
rect 14702 26238 14754 26290
rect 16270 26238 16322 26290
rect 18398 26238 18450 26290
rect 18846 26238 18898 26290
rect 19742 26238 19794 26290
rect 19854 26238 19906 26290
rect 20078 26238 20130 26290
rect 21310 26238 21362 26290
rect 21870 26238 21922 26290
rect 22206 26238 22258 26290
rect 22430 26238 22482 26290
rect 22878 26238 22930 26290
rect 23102 26238 23154 26290
rect 23774 26238 23826 26290
rect 26798 26238 26850 26290
rect 27806 26238 27858 26290
rect 37886 26238 37938 26290
rect 11566 26126 11618 26178
rect 13806 26126 13858 26178
rect 16718 26126 16770 26178
rect 19518 26126 19570 26178
rect 27582 26126 27634 26178
rect 11790 26014 11842 26066
rect 13470 26014 13522 26066
rect 14030 26014 14082 26066
rect 20526 26014 20578 26066
rect 5876 25846 5928 25898
rect 5980 25846 6032 25898
rect 6084 25846 6136 25898
rect 15200 25846 15252 25898
rect 15304 25846 15356 25898
rect 15408 25846 15460 25898
rect 24524 25846 24576 25898
rect 24628 25846 24680 25898
rect 24732 25846 24784 25898
rect 33848 25846 33900 25898
rect 33952 25846 34004 25898
rect 34056 25846 34108 25898
rect 15262 25678 15314 25730
rect 18398 25678 18450 25730
rect 18958 25678 19010 25730
rect 22766 25678 22818 25730
rect 23326 25678 23378 25730
rect 24670 25678 24722 25730
rect 14926 25566 14978 25618
rect 16158 25566 16210 25618
rect 18846 25566 18898 25618
rect 11678 25454 11730 25506
rect 15150 25454 15202 25506
rect 16830 25454 16882 25506
rect 17390 25454 17442 25506
rect 17950 25454 18002 25506
rect 20526 25454 20578 25506
rect 22878 25454 22930 25506
rect 23102 25454 23154 25506
rect 24446 25454 24498 25506
rect 26574 25454 26626 25506
rect 26798 25454 26850 25506
rect 26910 25454 26962 25506
rect 2046 25342 2098 25394
rect 12462 25342 12514 25394
rect 12798 25342 12850 25394
rect 16382 25342 16434 25394
rect 16494 25342 16546 25394
rect 17614 25342 17666 25394
rect 17726 25342 17778 25394
rect 20750 25342 20802 25394
rect 21310 25342 21362 25394
rect 21646 25342 21698 25394
rect 23438 25342 23490 25394
rect 23774 25342 23826 25394
rect 24110 25342 24162 25394
rect 25006 25342 25058 25394
rect 25342 25342 25394 25394
rect 25678 25342 25730 25394
rect 27358 25342 27410 25394
rect 27694 25342 27746 25394
rect 28030 25342 28082 25394
rect 37886 25342 37938 25394
rect 1710 25230 1762 25282
rect 11454 25230 11506 25282
rect 15262 25230 15314 25282
rect 15822 25230 15874 25282
rect 17166 25230 17218 25282
rect 19406 25230 19458 25282
rect 20078 25230 20130 25282
rect 38222 25230 38274 25282
rect 10538 25062 10590 25114
rect 10642 25062 10694 25114
rect 10746 25062 10798 25114
rect 19862 25062 19914 25114
rect 19966 25062 20018 25114
rect 20070 25062 20122 25114
rect 29186 25062 29238 25114
rect 29290 25062 29342 25114
rect 29394 25062 29446 25114
rect 38510 25062 38562 25114
rect 38614 25062 38666 25114
rect 38718 25062 38770 25114
rect 13022 24894 13074 24946
rect 14814 24894 14866 24946
rect 17390 24894 17442 24946
rect 22430 24894 22482 24946
rect 29374 24894 29426 24946
rect 1710 24782 1762 24834
rect 2046 24782 2098 24834
rect 9886 24782 9938 24834
rect 10222 24782 10274 24834
rect 11678 24782 11730 24834
rect 12014 24782 12066 24834
rect 12350 24782 12402 24834
rect 20526 24782 20578 24834
rect 20974 24782 21026 24834
rect 21198 24782 21250 24834
rect 24670 24782 24722 24834
rect 26686 24782 26738 24834
rect 27806 24782 27858 24834
rect 38222 24782 38274 24834
rect 9662 24670 9714 24722
rect 10558 24670 10610 24722
rect 11454 24670 11506 24722
rect 13358 24670 13410 24722
rect 13694 24670 13746 24722
rect 13806 24670 13858 24722
rect 14254 24670 14306 24722
rect 15150 24670 15202 24722
rect 15486 24670 15538 24722
rect 16046 24670 16098 24722
rect 17614 24670 17666 24722
rect 18958 24670 19010 24722
rect 20190 24670 20242 24722
rect 21422 24670 21474 24722
rect 21870 24670 21922 24722
rect 22094 24670 22146 24722
rect 24446 24670 24498 24722
rect 25230 24670 25282 24722
rect 26350 24670 26402 24722
rect 26574 24670 26626 24722
rect 27134 24670 27186 24722
rect 27470 24670 27522 24722
rect 28366 24670 28418 24722
rect 28702 24670 28754 24722
rect 29038 24670 29090 24722
rect 37886 24670 37938 24722
rect 16830 24558 16882 24610
rect 18398 24558 18450 24610
rect 19406 24558 19458 24610
rect 20862 24558 20914 24610
rect 25790 24558 25842 24610
rect 28142 24558 28194 24610
rect 14030 24446 14082 24498
rect 14366 24446 14418 24498
rect 15598 24446 15650 24498
rect 15822 24446 15874 24498
rect 16158 24446 16210 24498
rect 18286 24446 18338 24498
rect 18846 24446 18898 24498
rect 19182 24446 19234 24498
rect 19518 24446 19570 24498
rect 25566 24446 25618 24498
rect 5876 24278 5928 24330
rect 5980 24278 6032 24330
rect 6084 24278 6136 24330
rect 15200 24278 15252 24330
rect 15304 24278 15356 24330
rect 15408 24278 15460 24330
rect 24524 24278 24576 24330
rect 24628 24278 24680 24330
rect 24732 24278 24784 24330
rect 33848 24278 33900 24330
rect 33952 24278 34004 24330
rect 34056 24278 34108 24330
rect 10222 24110 10274 24162
rect 10670 24110 10722 24162
rect 14478 24110 14530 24162
rect 14702 24110 14754 24162
rect 14814 24110 14866 24162
rect 24446 24110 24498 24162
rect 28142 24110 28194 24162
rect 12350 23998 12402 24050
rect 9438 23886 9490 23938
rect 9998 23886 10050 23938
rect 10446 23886 10498 23938
rect 11566 23886 11618 23938
rect 12126 23886 12178 23938
rect 12574 23886 12626 23938
rect 12798 23886 12850 23938
rect 16606 23886 16658 23938
rect 17278 23886 17330 23938
rect 17838 23886 17890 23938
rect 18286 23886 18338 23938
rect 18734 23886 18786 23938
rect 19518 23886 19570 23938
rect 23550 23886 23602 23938
rect 24222 23886 24274 23938
rect 26350 23886 26402 23938
rect 26574 23886 26626 23938
rect 26686 23886 26738 23938
rect 27918 23886 27970 23938
rect 2046 23774 2098 23826
rect 9662 23774 9714 23826
rect 11790 23774 11842 23826
rect 14366 23774 14418 23826
rect 15374 23774 15426 23826
rect 16270 23774 16322 23826
rect 17390 23774 17442 23826
rect 17726 23774 17778 23826
rect 19182 23774 19234 23826
rect 21310 23774 21362 23826
rect 21646 23774 21698 23826
rect 21982 23774 22034 23826
rect 22318 23774 22370 23826
rect 22990 23774 23042 23826
rect 23326 23774 23378 23826
rect 24782 23774 24834 23826
rect 25118 23774 25170 23826
rect 25454 23774 25506 23826
rect 28478 23774 28530 23826
rect 29150 23774 29202 23826
rect 29486 23774 29538 23826
rect 37886 23774 37938 23826
rect 1710 23662 1762 23714
rect 10558 23662 10610 23714
rect 12686 23662 12738 23714
rect 18510 23662 18562 23714
rect 22654 23662 22706 23714
rect 27134 23662 27186 23714
rect 38222 23662 38274 23714
rect 10538 23494 10590 23546
rect 10642 23494 10694 23546
rect 10746 23494 10798 23546
rect 19862 23494 19914 23546
rect 19966 23494 20018 23546
rect 20070 23494 20122 23546
rect 29186 23494 29238 23546
rect 29290 23494 29342 23546
rect 29394 23494 29446 23546
rect 38510 23494 38562 23546
rect 38614 23494 38666 23546
rect 38718 23494 38770 23546
rect 10110 23326 10162 23378
rect 14030 23326 14082 23378
rect 16494 23326 16546 23378
rect 17726 23326 17778 23378
rect 24110 23326 24162 23378
rect 26462 23326 26514 23378
rect 27582 23326 27634 23378
rect 27918 23326 27970 23378
rect 31278 23326 31330 23378
rect 32398 23326 32450 23378
rect 1710 23214 1762 23266
rect 12238 23214 12290 23266
rect 12574 23214 12626 23266
rect 18174 23214 18226 23266
rect 19966 23214 20018 23266
rect 20302 23214 20354 23266
rect 20638 23214 20690 23266
rect 23774 23214 23826 23266
rect 27246 23214 27298 23266
rect 29374 23214 29426 23266
rect 30606 23214 30658 23266
rect 38222 23214 38274 23266
rect 2046 23102 2098 23154
rect 10446 23102 10498 23154
rect 13694 23102 13746 23154
rect 13918 23102 13970 23154
rect 14142 23102 14194 23154
rect 14814 23102 14866 23154
rect 15038 23102 15090 23154
rect 16718 23102 16770 23154
rect 17390 23102 17442 23154
rect 18846 23102 18898 23154
rect 19406 23102 19458 23154
rect 23438 23102 23490 23154
rect 24446 23102 24498 23154
rect 26126 23102 26178 23154
rect 28254 23102 28306 23154
rect 29038 23102 29090 23154
rect 30270 23102 30322 23154
rect 31054 23102 31106 23154
rect 32062 23102 32114 23154
rect 37886 23102 37938 23154
rect 14702 22990 14754 23042
rect 19182 22990 19234 23042
rect 21310 22990 21362 23042
rect 13470 22878 13522 22930
rect 14590 22878 14642 22930
rect 18062 22878 18114 22930
rect 18958 22878 19010 22930
rect 19518 22878 19570 22930
rect 5876 22710 5928 22762
rect 5980 22710 6032 22762
rect 6084 22710 6136 22762
rect 15200 22710 15252 22762
rect 15304 22710 15356 22762
rect 15408 22710 15460 22762
rect 24524 22710 24576 22762
rect 24628 22710 24680 22762
rect 24732 22710 24784 22762
rect 33848 22710 33900 22762
rect 33952 22710 34004 22762
rect 34056 22710 34108 22762
rect 9998 22542 10050 22594
rect 10110 22542 10162 22594
rect 10558 22542 10610 22594
rect 12014 22542 12066 22594
rect 17838 22542 17890 22594
rect 18174 22542 18226 22594
rect 18622 22542 18674 22594
rect 23326 22542 23378 22594
rect 30158 22542 30210 22594
rect 30718 22542 30770 22594
rect 31054 22542 31106 22594
rect 31950 22542 32002 22594
rect 32510 22542 32562 22594
rect 17838 22430 17890 22482
rect 18286 22430 18338 22482
rect 29598 22430 29650 22482
rect 30494 22430 30546 22482
rect 2718 22318 2770 22370
rect 10334 22318 10386 22370
rect 12126 22318 12178 22370
rect 12350 22318 12402 22370
rect 12574 22318 12626 22370
rect 14366 22318 14418 22370
rect 15038 22318 15090 22370
rect 16606 22318 16658 22370
rect 19406 22318 19458 22370
rect 21646 22318 21698 22370
rect 22430 22318 22482 22370
rect 22654 22318 22706 22370
rect 22878 22318 22930 22370
rect 23886 22318 23938 22370
rect 25678 22318 25730 22370
rect 29822 22318 29874 22370
rect 31390 22318 31442 22370
rect 31614 22318 31666 22370
rect 32286 22318 32338 22370
rect 1710 22206 1762 22258
rect 2046 22206 2098 22258
rect 9214 22206 9266 22258
rect 9550 22206 9602 22258
rect 11566 22206 11618 22258
rect 14142 22206 14194 22258
rect 14814 22206 14866 22258
rect 15486 22206 15538 22258
rect 16270 22206 16322 22258
rect 18734 22206 18786 22258
rect 19630 22206 19682 22258
rect 20414 22206 20466 22258
rect 21870 22206 21922 22258
rect 22542 22206 22594 22258
rect 23550 22206 23602 22258
rect 24334 22206 24386 22258
rect 24670 22206 24722 22258
rect 25902 22206 25954 22258
rect 26014 22206 26066 22258
rect 26462 22206 26514 22258
rect 26798 22206 26850 22258
rect 27134 22206 27186 22258
rect 27470 22206 27522 22258
rect 27806 22206 27858 22258
rect 28254 22206 28306 22258
rect 28590 22206 28642 22258
rect 37214 22206 37266 22258
rect 37886 22206 37938 22258
rect 38222 22206 38274 22258
rect 2382 22094 2434 22146
rect 10446 22094 10498 22146
rect 11230 22094 11282 22146
rect 12014 22094 12066 22146
rect 15822 22094 15874 22146
rect 17278 22094 17330 22146
rect 20078 22094 20130 22146
rect 20750 22094 20802 22146
rect 32846 22094 32898 22146
rect 37550 22094 37602 22146
rect 10538 21926 10590 21978
rect 10642 21926 10694 21978
rect 10746 21926 10798 21978
rect 19862 21926 19914 21978
rect 19966 21926 20018 21978
rect 20070 21926 20122 21978
rect 29186 21926 29238 21978
rect 29290 21926 29342 21978
rect 29394 21926 29446 21978
rect 38510 21926 38562 21978
rect 38614 21926 38666 21978
rect 38718 21926 38770 21978
rect 9998 21758 10050 21810
rect 13246 21758 13298 21810
rect 16718 21758 16770 21810
rect 17726 21758 17778 21810
rect 19294 21758 19346 21810
rect 21982 21758 22034 21810
rect 24222 21758 24274 21810
rect 27134 21758 27186 21810
rect 28926 21758 28978 21810
rect 1710 21646 1762 21698
rect 11006 21646 11058 21698
rect 18510 21646 18562 21698
rect 20302 21646 20354 21698
rect 21310 21646 21362 21698
rect 23326 21646 23378 21698
rect 23662 21646 23714 21698
rect 25566 21646 25618 21698
rect 26462 21646 26514 21698
rect 26686 21646 26738 21698
rect 27806 21646 27858 21698
rect 30158 21646 30210 21698
rect 32398 21646 32450 21698
rect 37886 21646 37938 21698
rect 38222 21646 38274 21698
rect 2046 21534 2098 21586
rect 9998 21534 10050 21586
rect 10558 21534 10610 21586
rect 11230 21534 11282 21586
rect 12350 21534 12402 21586
rect 12798 21534 12850 21586
rect 12910 21534 12962 21586
rect 13470 21534 13522 21586
rect 15262 21534 15314 21586
rect 15486 21534 15538 21586
rect 17390 21534 17442 21586
rect 18062 21534 18114 21586
rect 18286 21534 18338 21586
rect 18846 21534 18898 21586
rect 19518 21534 19570 21586
rect 19966 21534 20018 21586
rect 20974 21534 21026 21586
rect 21758 21534 21810 21586
rect 23214 21534 23266 21586
rect 23998 21534 24050 21586
rect 25230 21534 25282 21586
rect 26574 21534 26626 21586
rect 27470 21534 27522 21586
rect 27694 21534 27746 21586
rect 28254 21534 28306 21586
rect 28590 21534 28642 21586
rect 29934 21534 29986 21586
rect 32174 21534 32226 21586
rect 12238 21422 12290 21474
rect 15934 21422 15986 21474
rect 16382 21422 16434 21474
rect 16830 21422 16882 21474
rect 19070 21422 19122 21474
rect 22430 21422 22482 21474
rect 22878 21422 22930 21474
rect 10110 21310 10162 21362
rect 10334 21310 10386 21362
rect 12574 21310 12626 21362
rect 14926 21310 14978 21362
rect 15038 21310 15090 21362
rect 5876 21142 5928 21194
rect 5980 21142 6032 21194
rect 6084 21142 6136 21194
rect 15200 21142 15252 21194
rect 15304 21142 15356 21194
rect 15408 21142 15460 21194
rect 24524 21142 24576 21194
rect 24628 21142 24680 21194
rect 24732 21142 24784 21194
rect 33848 21142 33900 21194
rect 33952 21142 34004 21194
rect 34056 21142 34108 21194
rect 9998 20974 10050 21026
rect 10110 20974 10162 21026
rect 10670 20974 10722 21026
rect 12238 20974 12290 21026
rect 12350 20974 12402 21026
rect 12798 20974 12850 21026
rect 19406 20974 19458 21026
rect 24334 20974 24386 21026
rect 29486 20974 29538 21026
rect 30158 20974 30210 21026
rect 31390 20974 31442 21026
rect 10334 20862 10386 20914
rect 12574 20862 12626 20914
rect 14366 20862 14418 20914
rect 15598 20862 15650 20914
rect 17390 20862 17442 20914
rect 17726 20862 17778 20914
rect 20750 20862 20802 20914
rect 23326 20862 23378 20914
rect 30494 20862 30546 20914
rect 32286 20862 32338 20914
rect 10558 20750 10610 20802
rect 13470 20750 13522 20802
rect 14142 20750 14194 20802
rect 14590 20750 14642 20802
rect 14926 20750 14978 20802
rect 15710 20750 15762 20802
rect 15822 20750 15874 20802
rect 16830 20750 16882 20802
rect 18398 20750 18450 20802
rect 18734 20750 18786 20802
rect 19070 20750 19122 20802
rect 24110 20750 24162 20802
rect 29262 20750 29314 20802
rect 30718 20750 30770 20802
rect 31166 20750 31218 20802
rect 32062 20750 32114 20802
rect 37886 20750 37938 20802
rect 2046 20638 2098 20690
rect 11006 20638 11058 20690
rect 11342 20638 11394 20690
rect 12910 20638 12962 20690
rect 13806 20638 13858 20690
rect 16606 20638 16658 20690
rect 17838 20638 17890 20690
rect 18510 20638 18562 20690
rect 19854 20638 19906 20690
rect 20190 20638 20242 20690
rect 21310 20638 21362 20690
rect 21982 20638 22034 20690
rect 22766 20638 22818 20690
rect 23550 20638 23602 20690
rect 23774 20638 23826 20690
rect 24894 20638 24946 20690
rect 25230 20638 25282 20690
rect 26014 20638 26066 20690
rect 26350 20638 26402 20690
rect 27694 20638 27746 20690
rect 28030 20638 28082 20690
rect 31726 20638 31778 20690
rect 32958 20638 33010 20690
rect 33294 20638 33346 20690
rect 1710 20526 1762 20578
rect 14254 20526 14306 20578
rect 17278 20526 17330 20578
rect 21646 20526 21698 20578
rect 22318 20526 22370 20578
rect 29822 20526 29874 20578
rect 32622 20526 32674 20578
rect 38222 20526 38274 20578
rect 10538 20358 10590 20410
rect 10642 20358 10694 20410
rect 10746 20358 10798 20410
rect 19862 20358 19914 20410
rect 19966 20358 20018 20410
rect 20070 20358 20122 20410
rect 29186 20358 29238 20410
rect 29290 20358 29342 20410
rect 29394 20358 29446 20410
rect 38510 20358 38562 20410
rect 38614 20358 38666 20410
rect 38718 20358 38770 20410
rect 10558 20190 10610 20242
rect 12238 20190 12290 20242
rect 19518 20190 19570 20242
rect 19854 20190 19906 20242
rect 24334 20190 24386 20242
rect 27582 20190 27634 20242
rect 2046 20078 2098 20130
rect 9886 20078 9938 20130
rect 11566 20078 11618 20130
rect 12574 20078 12626 20130
rect 12910 20078 12962 20130
rect 13582 20078 13634 20130
rect 14142 20078 14194 20130
rect 15038 20078 15090 20130
rect 17502 20078 17554 20130
rect 17838 20078 17890 20130
rect 18846 20078 18898 20130
rect 21198 20078 21250 20130
rect 21646 20078 21698 20130
rect 22318 20078 22370 20130
rect 22990 20078 23042 20130
rect 23774 20078 23826 20130
rect 25566 20078 25618 20130
rect 27134 20078 27186 20130
rect 28590 20078 28642 20130
rect 29822 20078 29874 20130
rect 30158 20078 30210 20130
rect 32174 20078 32226 20130
rect 38222 20078 38274 20130
rect 1710 19966 1762 20018
rect 9662 19966 9714 20018
rect 10334 19966 10386 20018
rect 11230 19966 11282 20018
rect 12014 19966 12066 20018
rect 13246 19966 13298 20018
rect 14478 19966 14530 20018
rect 15150 19966 15202 20018
rect 15374 19966 15426 20018
rect 15598 19966 15650 20018
rect 16382 19966 16434 20018
rect 16830 19966 16882 20018
rect 18734 19966 18786 20018
rect 19070 19966 19122 20018
rect 20862 19966 20914 20018
rect 21982 19966 22034 20018
rect 22766 19966 22818 20018
rect 23326 19966 23378 20018
rect 23550 19966 23602 20018
rect 24110 19966 24162 20018
rect 25230 19966 25282 20018
rect 26910 19966 26962 20018
rect 27022 19966 27074 20018
rect 28254 19966 28306 20018
rect 31950 19966 32002 20018
rect 37886 19966 37938 20018
rect 2494 19854 2546 19906
rect 18510 19854 18562 19906
rect 20526 19854 20578 19906
rect 5876 19574 5928 19626
rect 5980 19574 6032 19626
rect 6084 19574 6136 19626
rect 15200 19574 15252 19626
rect 15304 19574 15356 19626
rect 15408 19574 15460 19626
rect 24524 19574 24576 19626
rect 24628 19574 24680 19626
rect 24732 19574 24784 19626
rect 33848 19574 33900 19626
rect 33952 19574 34004 19626
rect 34056 19574 34108 19626
rect 24782 19406 24834 19458
rect 10558 19182 10610 19234
rect 12686 19182 12738 19234
rect 17838 19182 17890 19234
rect 18510 19182 18562 19234
rect 18846 19182 18898 19234
rect 19070 19182 19122 19234
rect 21534 19182 21586 19234
rect 22430 19182 22482 19234
rect 23214 19182 23266 19234
rect 23774 19182 23826 19234
rect 23998 19182 24050 19234
rect 24110 19182 24162 19234
rect 24334 19182 24386 19234
rect 25902 19182 25954 19234
rect 26574 19182 26626 19234
rect 27358 19182 27410 19234
rect 27582 19182 27634 19234
rect 30382 19182 30434 19234
rect 31950 19182 32002 19234
rect 10782 19070 10834 19122
rect 11454 19070 11506 19122
rect 14702 19070 14754 19122
rect 15038 19070 15090 19122
rect 15598 19070 15650 19122
rect 15934 19070 15986 19122
rect 16270 19070 16322 19122
rect 16606 19070 16658 19122
rect 16942 19070 16994 19122
rect 17278 19070 17330 19122
rect 18174 19070 18226 19122
rect 18734 19070 18786 19122
rect 19518 19070 19570 19122
rect 19742 19070 19794 19122
rect 20526 19070 20578 19122
rect 22654 19070 22706 19122
rect 23438 19070 23490 19122
rect 26910 19070 26962 19122
rect 27694 19070 27746 19122
rect 28142 19070 28194 19122
rect 29150 19070 29202 19122
rect 30942 19070 30994 19122
rect 37886 19070 37938 19122
rect 1710 18958 1762 19010
rect 2046 18958 2098 19010
rect 2494 18958 2546 19010
rect 11118 18958 11170 19010
rect 12910 18958 12962 19010
rect 14366 18958 14418 19010
rect 20078 18958 20130 19010
rect 21310 18958 21362 19010
rect 25230 18958 25282 19010
rect 26238 18958 26290 19010
rect 29486 18958 29538 19010
rect 30606 18958 30658 19010
rect 31278 18958 31330 19010
rect 32174 18958 32226 19010
rect 38222 18958 38274 19010
rect 10538 18790 10590 18842
rect 10642 18790 10694 18842
rect 10746 18790 10798 18842
rect 19862 18790 19914 18842
rect 19966 18790 20018 18842
rect 20070 18790 20122 18842
rect 29186 18790 29238 18842
rect 29290 18790 29342 18842
rect 29394 18790 29446 18842
rect 38510 18790 38562 18842
rect 38614 18790 38666 18842
rect 38718 18790 38770 18842
rect 16830 18622 16882 18674
rect 18062 18622 18114 18674
rect 20190 18622 20242 18674
rect 22430 18622 22482 18674
rect 23662 18622 23714 18674
rect 28030 18622 28082 18674
rect 30494 18622 30546 18674
rect 31950 18622 32002 18674
rect 1710 18510 1762 18562
rect 10894 18510 10946 18562
rect 11566 18510 11618 18562
rect 13358 18510 13410 18562
rect 14814 18510 14866 18562
rect 18734 18510 18786 18562
rect 21646 18510 21698 18562
rect 22654 18510 22706 18562
rect 24334 18510 24386 18562
rect 25790 18510 25842 18562
rect 26126 18510 26178 18562
rect 26462 18510 26514 18562
rect 27358 18510 27410 18562
rect 27582 18510 27634 18562
rect 38222 18510 38274 18562
rect 2046 18398 2098 18450
rect 10446 18398 10498 18450
rect 11118 18398 11170 18450
rect 11902 18398 11954 18450
rect 12238 18398 12290 18450
rect 12910 18398 12962 18450
rect 13022 18398 13074 18450
rect 13694 18398 13746 18450
rect 14478 18398 14530 18450
rect 15374 18398 15426 18450
rect 17614 18398 17666 18450
rect 18398 18398 18450 18450
rect 18958 18398 19010 18450
rect 19854 18398 19906 18450
rect 21422 18398 21474 18450
rect 21758 18398 21810 18450
rect 22206 18398 22258 18450
rect 22878 18398 22930 18450
rect 23326 18398 23378 18450
rect 24110 18398 24162 18450
rect 25454 18398 25506 18450
rect 27470 18398 27522 18450
rect 29598 18398 29650 18450
rect 30158 18398 30210 18450
rect 31054 18398 31106 18450
rect 37886 18398 37938 18450
rect 14254 18286 14306 18338
rect 16158 18286 16210 18338
rect 19518 18286 19570 18338
rect 21086 18286 21138 18338
rect 31390 18286 31442 18338
rect 9886 18174 9938 18226
rect 9998 18174 10050 18226
rect 10222 18174 10274 18226
rect 10558 18174 10610 18226
rect 12462 18174 12514 18226
rect 12686 18174 12738 18226
rect 15262 18174 15314 18226
rect 16046 18174 16098 18226
rect 29822 18174 29874 18226
rect 30830 18174 30882 18226
rect 31614 18174 31666 18226
rect 5876 18006 5928 18058
rect 5980 18006 6032 18058
rect 6084 18006 6136 18058
rect 15200 18006 15252 18058
rect 15304 18006 15356 18058
rect 15408 18006 15460 18058
rect 24524 18006 24576 18058
rect 24628 18006 24680 18058
rect 24732 18006 24784 18058
rect 33848 18006 33900 18058
rect 33952 18006 34004 18058
rect 34056 18006 34108 18058
rect 10222 17838 10274 17890
rect 10446 17838 10498 17890
rect 10670 17838 10722 17890
rect 10782 17838 10834 17890
rect 12238 17838 12290 17890
rect 12910 17838 12962 17890
rect 14702 17838 14754 17890
rect 15710 17838 15762 17890
rect 25342 17838 25394 17890
rect 19406 17726 19458 17778
rect 24222 17726 24274 17778
rect 26350 17726 26402 17778
rect 2718 17614 2770 17666
rect 8766 17614 8818 17666
rect 10110 17614 10162 17666
rect 11342 17614 11394 17666
rect 12350 17614 12402 17666
rect 12574 17614 12626 17666
rect 12798 17614 12850 17666
rect 14814 17614 14866 17666
rect 15038 17614 15090 17666
rect 15486 17614 15538 17666
rect 15934 17614 15986 17666
rect 16606 17614 16658 17666
rect 18174 17614 18226 17666
rect 18286 17614 18338 17666
rect 18622 17614 18674 17666
rect 21758 17614 21810 17666
rect 22766 17614 22818 17666
rect 24894 17614 24946 17666
rect 25566 17614 25618 17666
rect 27246 17614 27298 17666
rect 27470 17614 27522 17666
rect 31166 17614 31218 17666
rect 31390 17614 31442 17666
rect 37214 17614 37266 17666
rect 1710 17502 1762 17554
rect 2046 17502 2098 17554
rect 8430 17502 8482 17554
rect 15150 17502 15202 17554
rect 17726 17502 17778 17554
rect 18398 17502 18450 17554
rect 19742 17502 19794 17554
rect 20078 17502 20130 17554
rect 23438 17502 23490 17554
rect 23774 17502 23826 17554
rect 24334 17502 24386 17554
rect 24670 17502 24722 17554
rect 25902 17502 25954 17554
rect 26126 17502 26178 17554
rect 27358 17502 27410 17554
rect 27918 17502 27970 17554
rect 28254 17502 28306 17554
rect 28590 17502 28642 17554
rect 29150 17502 29202 17554
rect 29486 17502 29538 17554
rect 31726 17502 31778 17554
rect 32062 17502 32114 17554
rect 32398 17502 32450 17554
rect 37886 17502 37938 17554
rect 38222 17502 38274 17554
rect 2382 17390 2434 17442
rect 11118 17390 11170 17442
rect 15598 17390 15650 17442
rect 16942 17390 16994 17442
rect 17390 17390 17442 17442
rect 19070 17390 19122 17442
rect 22094 17390 22146 17442
rect 23102 17390 23154 17442
rect 25230 17390 25282 17442
rect 37550 17390 37602 17442
rect 10538 17222 10590 17274
rect 10642 17222 10694 17274
rect 10746 17222 10798 17274
rect 19862 17222 19914 17274
rect 19966 17222 20018 17274
rect 20070 17222 20122 17274
rect 29186 17222 29238 17274
rect 29290 17222 29342 17274
rect 29394 17222 29446 17274
rect 38510 17222 38562 17274
rect 38614 17222 38666 17274
rect 38718 17222 38770 17274
rect 18398 17054 18450 17106
rect 21646 17054 21698 17106
rect 23662 17054 23714 17106
rect 25678 17054 25730 17106
rect 1710 16942 1762 16994
rect 2046 16942 2098 16994
rect 10782 16942 10834 16994
rect 13358 16942 13410 16994
rect 16494 16942 16546 16994
rect 17614 16942 17666 16994
rect 17838 16942 17890 16994
rect 19070 16942 19122 16994
rect 19406 16942 19458 16994
rect 19966 16942 20018 16994
rect 20638 16942 20690 16994
rect 21982 16942 22034 16994
rect 22318 16942 22370 16994
rect 22878 16942 22930 16994
rect 23214 16942 23266 16994
rect 25342 16942 25394 16994
rect 26574 16942 26626 16994
rect 27246 16942 27298 16994
rect 28366 16942 28418 16994
rect 29150 16942 29202 16994
rect 30718 16942 30770 16994
rect 32510 16942 32562 16994
rect 38222 16942 38274 16994
rect 10222 16830 10274 16882
rect 12238 16830 12290 16882
rect 13022 16830 13074 16882
rect 13582 16830 13634 16882
rect 14702 16830 14754 16882
rect 15038 16830 15090 16882
rect 15486 16830 15538 16882
rect 15934 16830 15986 16882
rect 17390 16830 17442 16882
rect 18174 16830 18226 16882
rect 20190 16830 20242 16882
rect 20974 16830 21026 16882
rect 21422 16830 21474 16882
rect 26238 16830 26290 16882
rect 26910 16830 26962 16882
rect 27134 16830 27186 16882
rect 27694 16830 27746 16882
rect 28030 16830 28082 16882
rect 28926 16830 28978 16882
rect 29486 16830 29538 16882
rect 30046 16830 30098 16882
rect 30382 16830 30434 16882
rect 31278 16830 31330 16882
rect 31838 16830 31890 16882
rect 32174 16830 32226 16882
rect 37886 16830 37938 16882
rect 10446 16718 10498 16770
rect 15150 16718 15202 16770
rect 29710 16718 29762 16770
rect 31502 16718 31554 16770
rect 10110 16606 10162 16658
rect 10670 16606 10722 16658
rect 12462 16606 12514 16658
rect 12686 16606 12738 16658
rect 12910 16606 12962 16658
rect 14814 16606 14866 16658
rect 15710 16606 15762 16658
rect 16046 16606 16098 16658
rect 16382 16606 16434 16658
rect 5876 16438 5928 16490
rect 5980 16438 6032 16490
rect 6084 16438 6136 16490
rect 15200 16438 15252 16490
rect 15304 16438 15356 16490
rect 15408 16438 15460 16490
rect 24524 16438 24576 16490
rect 24628 16438 24680 16490
rect 24732 16438 24784 16490
rect 33848 16438 33900 16490
rect 33952 16438 34004 16490
rect 34056 16438 34108 16490
rect 10334 16270 10386 16322
rect 10782 16270 10834 16322
rect 12238 16270 12290 16322
rect 15486 16270 15538 16322
rect 29822 16270 29874 16322
rect 31502 16270 31554 16322
rect 10558 16158 10610 16210
rect 12574 16158 12626 16210
rect 17390 16158 17442 16210
rect 17726 16158 17778 16210
rect 22990 16158 23042 16210
rect 24446 16158 24498 16210
rect 29598 16158 29650 16210
rect 31278 16158 31330 16210
rect 2046 16046 2098 16098
rect 8542 16046 8594 16098
rect 8878 16046 8930 16098
rect 9550 16046 9602 16098
rect 10110 16046 10162 16098
rect 12350 16046 12402 16098
rect 12798 16046 12850 16098
rect 14926 16046 14978 16098
rect 16718 16046 16770 16098
rect 18062 16046 18114 16098
rect 18286 16046 18338 16098
rect 18734 16046 18786 16098
rect 19182 16046 19234 16098
rect 19742 16046 19794 16098
rect 23326 16046 23378 16098
rect 23774 16046 23826 16098
rect 24670 16046 24722 16098
rect 25006 16046 25058 16098
rect 9102 15934 9154 15986
rect 9774 15934 9826 15986
rect 10894 15934 10946 15986
rect 11454 15934 11506 15986
rect 11790 15934 11842 15986
rect 12910 15934 12962 15986
rect 13470 15934 13522 15986
rect 13806 15934 13858 15986
rect 15150 15934 15202 15986
rect 15598 15934 15650 15986
rect 15934 15934 15986 15986
rect 16942 15934 16994 15986
rect 17950 15934 18002 15986
rect 21310 15934 21362 15986
rect 21646 15934 21698 15986
rect 22094 15934 22146 15986
rect 23102 15934 23154 15986
rect 24894 15934 24946 15986
rect 25454 15934 25506 15986
rect 25678 15934 25730 15986
rect 30158 15934 30210 15986
rect 30494 15934 30546 15986
rect 30830 15934 30882 15986
rect 31838 15934 31890 15986
rect 32174 15934 32226 15986
rect 37886 15934 37938 15986
rect 1710 15822 1762 15874
rect 14478 15822 14530 15874
rect 16270 15822 16322 15874
rect 18958 15822 19010 15874
rect 20078 15822 20130 15874
rect 21982 15822 22034 15874
rect 23998 15822 24050 15874
rect 26014 15822 26066 15874
rect 32510 15822 32562 15874
rect 38222 15822 38274 15874
rect 10538 15654 10590 15706
rect 10642 15654 10694 15706
rect 10746 15654 10798 15706
rect 19862 15654 19914 15706
rect 19966 15654 20018 15706
rect 20070 15654 20122 15706
rect 29186 15654 29238 15706
rect 29290 15654 29342 15706
rect 29394 15654 29446 15706
rect 38510 15654 38562 15706
rect 38614 15654 38666 15706
rect 38718 15654 38770 15706
rect 12462 15486 12514 15538
rect 14030 15486 14082 15538
rect 16046 15486 16098 15538
rect 16830 15486 16882 15538
rect 19406 15486 19458 15538
rect 23886 15486 23938 15538
rect 24558 15486 24610 15538
rect 28814 15486 28866 15538
rect 1710 15374 1762 15426
rect 2046 15374 2098 15426
rect 9998 15374 10050 15426
rect 10334 15374 10386 15426
rect 10670 15374 10722 15426
rect 11006 15374 11058 15426
rect 11342 15374 11394 15426
rect 12798 15374 12850 15426
rect 14926 15374 14978 15426
rect 15262 15374 15314 15426
rect 17614 15374 17666 15426
rect 17838 15374 17890 15426
rect 18622 15374 18674 15426
rect 22990 15374 23042 15426
rect 24222 15374 24274 15426
rect 25566 15374 25618 15426
rect 25902 15374 25954 15426
rect 26350 15374 26402 15426
rect 37886 15374 37938 15426
rect 38222 15374 38274 15426
rect 13022 15262 13074 15314
rect 14590 15262 14642 15314
rect 17502 15262 17554 15314
rect 18174 15262 18226 15314
rect 18398 15262 18450 15314
rect 18846 15262 18898 15314
rect 19630 15262 19682 15314
rect 20974 15262 21026 15314
rect 21086 15262 21138 15314
rect 21198 15262 21250 15314
rect 22318 15262 22370 15314
rect 22654 15262 22706 15314
rect 23662 15262 23714 15314
rect 26462 15262 26514 15314
rect 26574 15262 26626 15314
rect 27358 15262 27410 15314
rect 27582 15262 27634 15314
rect 27694 15262 27746 15314
rect 28142 15262 28194 15314
rect 28478 15262 28530 15314
rect 12014 15150 12066 15202
rect 14254 15150 14306 15202
rect 14478 15150 14530 15202
rect 21646 15150 21698 15202
rect 27022 15038 27074 15090
rect 5876 14870 5928 14922
rect 5980 14870 6032 14922
rect 6084 14870 6136 14922
rect 15200 14870 15252 14922
rect 15304 14870 15356 14922
rect 15408 14870 15460 14922
rect 24524 14870 24576 14922
rect 24628 14870 24680 14922
rect 24732 14870 24784 14922
rect 33848 14870 33900 14922
rect 33952 14870 34004 14922
rect 34056 14870 34108 14922
rect 10446 14702 10498 14754
rect 10894 14702 10946 14754
rect 14142 14702 14194 14754
rect 20638 14702 20690 14754
rect 8542 14590 8594 14642
rect 11678 14590 11730 14642
rect 24222 14590 24274 14642
rect 24558 14590 24610 14642
rect 29150 14590 29202 14642
rect 8878 14478 8930 14530
rect 10222 14478 10274 14530
rect 10670 14478 10722 14530
rect 12238 14478 12290 14530
rect 12798 14478 12850 14530
rect 13470 14478 13522 14530
rect 13694 14478 13746 14530
rect 13918 14478 13970 14530
rect 14814 14478 14866 14530
rect 14926 14478 14978 14530
rect 15150 14478 15202 14530
rect 15598 14478 15650 14530
rect 18510 14478 18562 14530
rect 19182 14478 19234 14530
rect 19630 14478 19682 14530
rect 20190 14478 20242 14530
rect 20526 14478 20578 14530
rect 21310 14478 21362 14530
rect 22878 14478 22930 14530
rect 23102 14478 23154 14530
rect 23438 14478 23490 14530
rect 24782 14478 24834 14530
rect 25678 14478 25730 14530
rect 27022 14478 27074 14530
rect 29374 14478 29426 14530
rect 2046 14366 2098 14418
rect 9214 14366 9266 14418
rect 9886 14366 9938 14418
rect 11902 14366 11954 14418
rect 15262 14366 15314 14418
rect 15710 14366 15762 14418
rect 16718 14366 16770 14418
rect 17054 14366 17106 14418
rect 17726 14366 17778 14418
rect 17950 14366 18002 14418
rect 18062 14366 18114 14418
rect 18734 14366 18786 14418
rect 23214 14366 23266 14418
rect 25454 14366 25506 14418
rect 28254 14366 28306 14418
rect 28590 14366 28642 14418
rect 29710 14366 29762 14418
rect 30046 14366 30098 14418
rect 37886 14366 37938 14418
rect 1710 14254 1762 14306
rect 9550 14254 9602 14306
rect 10334 14254 10386 14306
rect 12574 14254 12626 14306
rect 13582 14254 13634 14306
rect 16046 14254 16098 14306
rect 16382 14254 16434 14306
rect 17502 14254 17554 14306
rect 21870 14254 21922 14306
rect 23886 14254 23938 14306
rect 25118 14254 25170 14306
rect 27246 14254 27298 14306
rect 30382 14254 30434 14306
rect 38222 14254 38274 14306
rect 10538 14086 10590 14138
rect 10642 14086 10694 14138
rect 10746 14086 10798 14138
rect 19862 14086 19914 14138
rect 19966 14086 20018 14138
rect 20070 14086 20122 14138
rect 29186 14086 29238 14138
rect 29290 14086 29342 14138
rect 29394 14086 29446 14138
rect 38510 14086 38562 14138
rect 38614 14086 38666 14138
rect 38718 14086 38770 14138
rect 13246 13918 13298 13970
rect 18846 13918 18898 13970
rect 19518 13918 19570 13970
rect 22318 13918 22370 13970
rect 1710 13806 1762 13858
rect 2046 13806 2098 13858
rect 11454 13806 11506 13858
rect 12686 13806 12738 13858
rect 14590 13806 14642 13858
rect 14926 13806 14978 13858
rect 16830 13806 16882 13858
rect 17726 13806 17778 13858
rect 19630 13806 19682 13858
rect 20526 13806 20578 13858
rect 23214 13806 23266 13858
rect 24110 13806 24162 13858
rect 24446 13806 24498 13858
rect 25566 13806 25618 13858
rect 26798 13806 26850 13858
rect 27918 13806 27970 13858
rect 29038 13806 29090 13858
rect 38222 13806 38274 13858
rect 10334 13694 10386 13746
rect 10558 13694 10610 13746
rect 11006 13694 11058 13746
rect 11678 13694 11730 13746
rect 12462 13694 12514 13746
rect 16158 13694 16210 13746
rect 16606 13694 16658 13746
rect 17614 13694 17666 13746
rect 17950 13694 18002 13746
rect 18174 13694 18226 13746
rect 19070 13694 19122 13746
rect 20078 13694 20130 13746
rect 21758 13694 21810 13746
rect 23102 13694 23154 13746
rect 23550 13694 23602 13746
rect 25230 13694 25282 13746
rect 26574 13694 26626 13746
rect 26686 13694 26738 13746
rect 27582 13694 27634 13746
rect 27806 13694 27858 13746
rect 28366 13694 28418 13746
rect 28702 13694 28754 13746
rect 37886 13694 37938 13746
rect 14366 13582 14418 13634
rect 15710 13582 15762 13634
rect 18622 13582 18674 13634
rect 22878 13582 22930 13634
rect 10782 13470 10834 13522
rect 11118 13470 11170 13522
rect 15598 13470 15650 13522
rect 23886 13470 23938 13522
rect 27246 13470 27298 13522
rect 5876 13302 5928 13354
rect 5980 13302 6032 13354
rect 6084 13302 6136 13354
rect 15200 13302 15252 13354
rect 15304 13302 15356 13354
rect 15408 13302 15460 13354
rect 24524 13302 24576 13354
rect 24628 13302 24680 13354
rect 24732 13302 24784 13354
rect 33848 13302 33900 13354
rect 33952 13302 34004 13354
rect 34056 13302 34108 13354
rect 10222 13134 10274 13186
rect 10334 13134 10386 13186
rect 10782 13134 10834 13186
rect 11118 13134 11170 13186
rect 11454 13134 11506 13186
rect 13694 13134 13746 13186
rect 14142 13134 14194 13186
rect 15262 13134 15314 13186
rect 16158 13134 16210 13186
rect 24782 13134 24834 13186
rect 25118 13134 25170 13186
rect 11454 13022 11506 13074
rect 16046 13022 16098 13074
rect 17502 13022 17554 13074
rect 21422 13022 21474 13074
rect 2046 12910 2098 12962
rect 2718 12910 2770 12962
rect 10558 12910 10610 12962
rect 12798 12910 12850 12962
rect 13470 12910 13522 12962
rect 13918 12910 13970 12962
rect 14926 12910 14978 12962
rect 15150 12910 15202 12962
rect 15822 12910 15874 12962
rect 17054 12910 17106 12962
rect 17726 12910 17778 12962
rect 18062 12910 18114 12962
rect 18510 12910 18562 12962
rect 19070 12910 19122 12962
rect 20414 12910 20466 12962
rect 21982 12910 22034 12962
rect 22094 12910 22146 12962
rect 22206 12910 22258 12962
rect 22654 12910 22706 12962
rect 23886 12910 23938 12962
rect 24558 12910 24610 12962
rect 25454 12910 25506 12962
rect 27470 12910 27522 12962
rect 37886 12910 37938 12962
rect 1710 12798 1762 12850
rect 10894 12798 10946 12850
rect 14814 12798 14866 12850
rect 15710 12798 15762 12850
rect 16830 12798 16882 12850
rect 17950 12798 18002 12850
rect 20750 12798 20802 12850
rect 22878 12798 22930 12850
rect 23102 12798 23154 12850
rect 25790 12798 25842 12850
rect 26462 12798 26514 12850
rect 26798 12798 26850 12850
rect 37214 12798 37266 12850
rect 38222 12798 38274 12850
rect 2382 12686 2434 12738
rect 12574 12686 12626 12738
rect 13582 12686 13634 12738
rect 18846 12686 18898 12738
rect 19742 12686 19794 12738
rect 20078 12686 20130 12738
rect 23438 12686 23490 12738
rect 24110 12686 24162 12738
rect 26126 12686 26178 12738
rect 27134 12686 27186 12738
rect 27806 12686 27858 12738
rect 37550 12686 37602 12738
rect 10538 12518 10590 12570
rect 10642 12518 10694 12570
rect 10746 12518 10798 12570
rect 19862 12518 19914 12570
rect 19966 12518 20018 12570
rect 20070 12518 20122 12570
rect 29186 12518 29238 12570
rect 29290 12518 29342 12570
rect 29394 12518 29446 12570
rect 38510 12518 38562 12570
rect 38614 12518 38666 12570
rect 38718 12518 38770 12570
rect 10670 12350 10722 12402
rect 16270 12350 16322 12402
rect 17502 12350 17554 12402
rect 25790 12350 25842 12402
rect 1710 12238 1762 12290
rect 2046 12238 2098 12290
rect 13806 12238 13858 12290
rect 24558 12238 24610 12290
rect 27358 12238 27410 12290
rect 29038 12238 29090 12290
rect 37886 12238 37938 12290
rect 38222 12238 38274 12290
rect 10222 12126 10274 12178
rect 10334 12126 10386 12178
rect 11790 12126 11842 12178
rect 12238 12126 12290 12178
rect 12686 12126 12738 12178
rect 12910 12126 12962 12178
rect 13134 12126 13186 12178
rect 13358 12126 13410 12178
rect 13470 12126 13522 12178
rect 14030 12126 14082 12178
rect 15486 12126 15538 12178
rect 23438 12126 23490 12178
rect 24222 12126 24274 12178
rect 25230 12126 25282 12178
rect 25454 12126 25506 12178
rect 26126 12126 26178 12178
rect 27022 12126 27074 12178
rect 27806 12126 27858 12178
rect 28030 12126 28082 12178
rect 28366 12126 28418 12178
rect 28702 12126 28754 12178
rect 10558 12014 10610 12066
rect 12014 12014 12066 12066
rect 15262 12014 15314 12066
rect 15822 12014 15874 12066
rect 15934 12014 15986 12066
rect 16382 12014 16434 12066
rect 21310 12014 21362 12066
rect 26350 12014 26402 12066
rect 26686 12014 26738 12066
rect 10782 11902 10834 11954
rect 11678 11902 11730 11954
rect 12350 11902 12402 11954
rect 14926 11902 14978 11954
rect 15038 11902 15090 11954
rect 5876 11734 5928 11786
rect 5980 11734 6032 11786
rect 6084 11734 6136 11786
rect 15200 11734 15252 11786
rect 15304 11734 15356 11786
rect 15408 11734 15460 11786
rect 24524 11734 24576 11786
rect 24628 11734 24680 11786
rect 24732 11734 24784 11786
rect 33848 11734 33900 11786
rect 33952 11734 34004 11786
rect 34056 11734 34108 11786
rect 27806 11566 27858 11618
rect 24222 11454 24274 11506
rect 25678 11454 25730 11506
rect 26238 11454 26290 11506
rect 26686 11454 26738 11506
rect 26910 11454 26962 11506
rect 27582 11454 27634 11506
rect 2046 11342 2098 11394
rect 10670 11342 10722 11394
rect 11342 11342 11394 11394
rect 13694 11342 13746 11394
rect 16046 11342 16098 11394
rect 16718 11342 16770 11394
rect 17278 11342 17330 11394
rect 17726 11342 17778 11394
rect 21310 11342 21362 11394
rect 22094 11342 22146 11394
rect 25566 11342 25618 11394
rect 37998 11342 38050 11394
rect 16158 11230 16210 11282
rect 16382 11230 16434 11282
rect 17390 11230 17442 11282
rect 17614 11230 17666 11282
rect 18398 11230 18450 11282
rect 19070 11230 19122 11282
rect 19406 11230 19458 11282
rect 19742 11230 19794 11282
rect 20078 11230 20130 11282
rect 20414 11230 20466 11282
rect 20750 11230 20802 11282
rect 24558 11230 24610 11282
rect 25006 11230 25058 11282
rect 25342 11230 25394 11282
rect 25790 11230 25842 11282
rect 28142 11230 28194 11282
rect 29150 11230 29202 11282
rect 1710 11118 1762 11170
rect 10334 11118 10386 11170
rect 11006 11118 11058 11170
rect 13470 11118 13522 11170
rect 15038 11118 15090 11170
rect 15486 11118 15538 11170
rect 16942 11118 16994 11170
rect 18174 11118 18226 11170
rect 18734 11118 18786 11170
rect 24782 11118 24834 11170
rect 25118 11118 25170 11170
rect 26126 11118 26178 11170
rect 27246 11118 27298 11170
rect 29486 11118 29538 11170
rect 38222 11118 38274 11170
rect 10538 10950 10590 11002
rect 10642 10950 10694 11002
rect 10746 10950 10798 11002
rect 19862 10950 19914 11002
rect 19966 10950 20018 11002
rect 20070 10950 20122 11002
rect 29186 10950 29238 11002
rect 29290 10950 29342 11002
rect 29394 10950 29446 11002
rect 38510 10950 38562 11002
rect 38614 10950 38666 11002
rect 38718 10950 38770 11002
rect 1710 10670 1762 10722
rect 2046 10670 2098 10722
rect 18062 10670 18114 10722
rect 18734 10670 18786 10722
rect 21758 10670 21810 10722
rect 37886 10670 37938 10722
rect 38222 10670 38274 10722
rect 18286 10558 18338 10610
rect 18958 10558 19010 10610
rect 24670 10558 24722 10610
rect 25342 10558 25394 10610
rect 27246 10446 27298 10498
rect 5876 10166 5928 10218
rect 5980 10166 6032 10218
rect 6084 10166 6136 10218
rect 15200 10166 15252 10218
rect 15304 10166 15356 10218
rect 15408 10166 15460 10218
rect 24524 10166 24576 10218
rect 24628 10166 24680 10218
rect 24732 10166 24784 10218
rect 33848 10166 33900 10218
rect 33952 10166 34004 10218
rect 34056 10166 34108 10218
rect 19406 9886 19458 9938
rect 27582 9886 27634 9938
rect 2046 9774 2098 9826
rect 26798 9774 26850 9826
rect 27806 9774 27858 9826
rect 28030 9774 28082 9826
rect 29150 9774 29202 9826
rect 37886 9774 37938 9826
rect 20526 9662 20578 9714
rect 20638 9662 20690 9714
rect 24894 9662 24946 9714
rect 31166 9662 31218 9714
rect 1710 9550 1762 9602
rect 20862 9550 20914 9602
rect 27246 9550 27298 9602
rect 27470 9550 27522 9602
rect 28366 9550 28418 9602
rect 38222 9550 38274 9602
rect 10538 9382 10590 9434
rect 10642 9382 10694 9434
rect 10746 9382 10798 9434
rect 19862 9382 19914 9434
rect 19966 9382 20018 9434
rect 20070 9382 20122 9434
rect 29186 9382 29238 9434
rect 29290 9382 29342 9434
rect 29394 9382 29446 9434
rect 38510 9382 38562 9434
rect 38614 9382 38666 9434
rect 38718 9382 38770 9434
rect 24334 9214 24386 9266
rect 1710 9102 1762 9154
rect 2046 9102 2098 9154
rect 19742 9102 19794 9154
rect 22878 9102 22930 9154
rect 23214 9102 23266 9154
rect 23326 9102 23378 9154
rect 24558 9102 24610 9154
rect 38222 9102 38274 9154
rect 18958 8990 19010 9042
rect 22318 8990 22370 9042
rect 22654 8990 22706 9042
rect 23550 8990 23602 9042
rect 23998 8990 24050 9042
rect 24110 8990 24162 9042
rect 25230 8990 25282 9042
rect 37998 8990 38050 9042
rect 21870 8878 21922 8930
rect 24670 8878 24722 8930
rect 27246 8878 27298 8930
rect 22990 8766 23042 8818
rect 5876 8598 5928 8650
rect 5980 8598 6032 8650
rect 6084 8598 6136 8650
rect 15200 8598 15252 8650
rect 15304 8598 15356 8650
rect 15408 8598 15460 8650
rect 24524 8598 24576 8650
rect 24628 8598 24680 8650
rect 24732 8598 24784 8650
rect 33848 8598 33900 8650
rect 33952 8598 34004 8650
rect 34056 8598 34108 8650
rect 3166 8318 3218 8370
rect 22878 8318 22930 8370
rect 2606 8206 2658 8258
rect 23886 8206 23938 8258
rect 24222 8206 24274 8258
rect 24446 8206 24498 8258
rect 24782 8206 24834 8258
rect 25230 8206 25282 8258
rect 25454 8206 25506 8258
rect 25790 8206 25842 8258
rect 25902 8206 25954 8258
rect 36430 8206 36482 8258
rect 37214 8206 37266 8258
rect 37886 8206 37938 8258
rect 1710 8094 1762 8146
rect 2046 8094 2098 8146
rect 22094 8094 22146 8146
rect 22430 8094 22482 8146
rect 23102 8094 23154 8146
rect 38222 8094 38274 8146
rect 2382 7982 2434 8034
rect 22878 7982 22930 8034
rect 23998 7982 24050 8034
rect 24558 7982 24610 8034
rect 25006 7982 25058 8034
rect 25566 7982 25618 8034
rect 27134 7982 27186 8034
rect 37550 7982 37602 8034
rect 10538 7814 10590 7866
rect 10642 7814 10694 7866
rect 10746 7814 10798 7866
rect 19862 7814 19914 7866
rect 19966 7814 20018 7866
rect 20070 7814 20122 7866
rect 29186 7814 29238 7866
rect 29290 7814 29342 7866
rect 29394 7814 29446 7866
rect 38510 7814 38562 7866
rect 38614 7814 38666 7866
rect 38718 7814 38770 7866
rect 22878 7646 22930 7698
rect 23550 7646 23602 7698
rect 24110 7646 24162 7698
rect 19630 7534 19682 7586
rect 23438 7534 23490 7586
rect 24222 7534 24274 7586
rect 24670 7534 24722 7586
rect 37886 7534 37938 7586
rect 38222 7534 38274 7586
rect 18958 7422 19010 7474
rect 22990 7422 23042 7474
rect 2382 7310 2434 7362
rect 21758 7310 21810 7362
rect 24558 7198 24610 7250
rect 5876 7030 5928 7082
rect 5980 7030 6032 7082
rect 6084 7030 6136 7082
rect 15200 7030 15252 7082
rect 15304 7030 15356 7082
rect 15408 7030 15460 7082
rect 24524 7030 24576 7082
rect 24628 7030 24680 7082
rect 24732 7030 24784 7082
rect 33848 7030 33900 7082
rect 33952 7030 34004 7082
rect 34056 7030 34108 7082
rect 37550 6638 37602 6690
rect 37998 6638 38050 6690
rect 38222 6414 38274 6466
rect 10538 6246 10590 6298
rect 10642 6246 10694 6298
rect 10746 6246 10798 6298
rect 19862 6246 19914 6298
rect 19966 6246 20018 6298
rect 20070 6246 20122 6298
rect 29186 6246 29238 6298
rect 29290 6246 29342 6298
rect 29394 6246 29446 6298
rect 38510 6246 38562 6298
rect 38614 6246 38666 6298
rect 38718 6246 38770 6298
rect 37662 6078 37714 6130
rect 37886 5966 37938 6018
rect 38222 5966 38274 6018
rect 5876 5462 5928 5514
rect 5980 5462 6032 5514
rect 6084 5462 6136 5514
rect 15200 5462 15252 5514
rect 15304 5462 15356 5514
rect 15408 5462 15460 5514
rect 24524 5462 24576 5514
rect 24628 5462 24680 5514
rect 24732 5462 24784 5514
rect 33848 5462 33900 5514
rect 33952 5462 34004 5514
rect 34056 5462 34108 5514
rect 37550 5182 37602 5234
rect 37998 5070 38050 5122
rect 38222 4846 38274 4898
rect 10538 4678 10590 4730
rect 10642 4678 10694 4730
rect 10746 4678 10798 4730
rect 19862 4678 19914 4730
rect 19966 4678 20018 4730
rect 20070 4678 20122 4730
rect 29186 4678 29238 4730
rect 29290 4678 29342 4730
rect 29394 4678 29446 4730
rect 38510 4678 38562 4730
rect 38614 4678 38666 4730
rect 38718 4678 38770 4730
rect 5966 4510 6018 4562
rect 6414 4510 6466 4562
rect 7646 4510 7698 4562
rect 9998 4510 10050 4562
rect 33854 4510 33906 4562
rect 37662 4510 37714 4562
rect 16382 4398 16434 4450
rect 16718 4398 16770 4450
rect 27134 4398 27186 4450
rect 37886 4398 37938 4450
rect 38222 4398 38274 4450
rect 5630 4286 5682 4338
rect 9102 4286 9154 4338
rect 9662 4286 9714 4338
rect 27358 4286 27410 4338
rect 5406 4174 5458 4226
rect 6974 4174 7026 4226
rect 8094 4174 8146 4226
rect 8654 4174 8706 4226
rect 10446 4174 10498 4226
rect 15934 4174 15986 4226
rect 20414 4174 20466 4226
rect 21534 4174 21586 4226
rect 22206 4174 22258 4226
rect 34638 4174 34690 4226
rect 5876 3894 5928 3946
rect 5980 3894 6032 3946
rect 6084 3894 6136 3946
rect 15200 3894 15252 3946
rect 15304 3894 15356 3946
rect 15408 3894 15460 3946
rect 24524 3894 24576 3946
rect 24628 3894 24680 3946
rect 24732 3894 24784 3946
rect 33848 3894 33900 3946
rect 33952 3894 34004 3946
rect 34056 3894 34108 3946
rect 37550 3614 37602 3666
rect 5854 3502 5906 3554
rect 7198 3502 7250 3554
rect 7870 3502 7922 3554
rect 8542 3502 8594 3554
rect 10222 3502 10274 3554
rect 10894 3502 10946 3554
rect 11566 3502 11618 3554
rect 12350 3502 12402 3554
rect 13694 3502 13746 3554
rect 14926 3502 14978 3554
rect 15486 3502 15538 3554
rect 16046 3502 16098 3554
rect 17278 3502 17330 3554
rect 17950 3502 18002 3554
rect 18510 3502 18562 3554
rect 19294 3502 19346 3554
rect 20190 3502 20242 3554
rect 21310 3502 21362 3554
rect 21982 3502 22034 3554
rect 22654 3502 22706 3554
rect 23326 3502 23378 3554
rect 24894 3502 24946 3554
rect 25566 3502 25618 3554
rect 26126 3502 26178 3554
rect 26798 3502 26850 3554
rect 27470 3502 27522 3554
rect 28590 3502 28642 3554
rect 29374 3502 29426 3554
rect 29934 3502 29986 3554
rect 30606 3502 30658 3554
rect 31278 3502 31330 3554
rect 32398 3502 32450 3554
rect 33742 3502 33794 3554
rect 34414 3502 34466 3554
rect 35086 3502 35138 3554
rect 37998 3502 38050 3554
rect 6414 3390 6466 3442
rect 6750 3390 6802 3442
rect 8094 3390 8146 3442
rect 8766 3390 8818 3442
rect 9550 3390 9602 3442
rect 9886 3390 9938 3442
rect 13358 3390 13410 3442
rect 14366 3390 14418 3442
rect 15710 3390 15762 3442
rect 16382 3390 16434 3442
rect 19854 3390 19906 3442
rect 22430 3390 22482 3442
rect 25230 3390 25282 3442
rect 25902 3390 25954 3442
rect 27246 3390 27298 3442
rect 29038 3390 29090 3442
rect 30382 3390 30434 3442
rect 32174 3390 32226 3442
rect 32846 3390 32898 3442
rect 33182 3390 33234 3442
rect 34190 3390 34242 3442
rect 34862 3390 34914 3442
rect 38222 3390 38274 3442
rect 6078 3278 6130 3330
rect 7422 3278 7474 3330
rect 10558 3278 10610 3330
rect 11230 3278 11282 3330
rect 11902 3278 11954 3330
rect 12574 3278 12626 3330
rect 14030 3278 14082 3330
rect 14702 3278 14754 3330
rect 17502 3278 17554 3330
rect 18174 3278 18226 3330
rect 18846 3278 18898 3330
rect 19518 3278 19570 3330
rect 21086 3278 21138 3330
rect 21758 3278 21810 3330
rect 23102 3278 23154 3330
rect 24558 3278 24610 3330
rect 26574 3278 26626 3330
rect 28366 3278 28418 3330
rect 29710 3278 29762 3330
rect 31054 3278 31106 3330
rect 33518 3278 33570 3330
rect 10538 3110 10590 3162
rect 10642 3110 10694 3162
rect 10746 3110 10798 3162
rect 19862 3110 19914 3162
rect 19966 3110 20018 3162
rect 20070 3110 20122 3162
rect 29186 3110 29238 3162
rect 29290 3110 29342 3162
rect 29394 3110 29446 3162
rect 38510 3110 38562 3162
rect 38614 3110 38666 3162
rect 38718 3110 38770 3162
rect 33630 2494 33682 2546
rect 34638 2494 34690 2546
rect 35086 2494 35138 2546
rect 30270 926 30322 978
rect 31054 926 31106 978
<< metal2 >>
rect 2688 39200 2800 40000
rect 3360 39200 3472 40000
rect 4032 39200 4144 40000
rect 4704 39200 4816 40000
rect 5376 39200 5488 40000
rect 6048 39200 6160 40000
rect 6720 39200 6832 40000
rect 7392 39200 7504 40000
rect 8064 39200 8176 40000
rect 8736 39200 8848 40000
rect 9408 39200 9520 40000
rect 10080 39200 10192 40000
rect 10752 39200 10864 40000
rect 11424 39200 11536 40000
rect 12096 39200 12208 40000
rect 12768 39200 12880 40000
rect 13440 39200 13552 40000
rect 14112 39200 14224 40000
rect 14784 39200 14896 40000
rect 15456 39200 15568 40000
rect 16128 39200 16240 40000
rect 16800 39200 16912 40000
rect 17472 39200 17584 40000
rect 18144 39200 18256 40000
rect 18816 39200 18928 40000
rect 19488 39200 19600 40000
rect 20160 39200 20272 40000
rect 20832 39200 20944 40000
rect 21504 39200 21616 40000
rect 22176 39200 22288 40000
rect 22848 39200 22960 40000
rect 23520 39200 23632 40000
rect 24192 39200 24304 40000
rect 24864 39200 24976 40000
rect 25536 39200 25648 40000
rect 26208 39200 26320 40000
rect 26880 39200 26992 40000
rect 27552 39200 27664 40000
rect 28224 39200 28336 40000
rect 28896 39200 29008 40000
rect 29568 39200 29680 40000
rect 30240 39200 30352 40000
rect 30912 39200 31024 40000
rect 31584 39200 31696 40000
rect 32256 39200 32368 40000
rect 32928 39200 33040 40000
rect 33600 39200 33712 40000
rect 34272 39200 34384 40000
rect 34944 39200 35056 40000
rect 35616 39200 35728 40000
rect 36288 39200 36400 40000
rect 2716 36484 2772 39200
rect 2716 36482 3220 36484
rect 2716 36430 2718 36482
rect 2770 36430 3220 36482
rect 2716 36428 3220 36430
rect 2716 36418 2772 36428
rect 2940 36260 2996 36270
rect 2940 36258 3108 36260
rect 2940 36206 2942 36258
rect 2994 36206 3108 36258
rect 2940 36204 3108 36206
rect 2940 36194 2996 36204
rect 1708 33122 1764 33134
rect 2044 33124 2100 33134
rect 1708 33070 1710 33122
rect 1762 33070 1764 33122
rect 1708 33012 1764 33070
rect 1708 32946 1764 32956
rect 1820 33122 2100 33124
rect 1820 33070 2046 33122
rect 2098 33070 2100 33122
rect 1820 33068 2100 33070
rect 1708 32674 1764 32686
rect 1708 32622 1710 32674
rect 1762 32622 1764 32674
rect 1708 32340 1764 32622
rect 1708 32274 1764 32284
rect 1708 31556 1764 31566
rect 1708 31462 1764 31500
rect 1708 31106 1764 31118
rect 1708 31054 1710 31106
rect 1762 31054 1764 31106
rect 1708 30324 1764 31054
rect 1708 30258 1764 30268
rect 1708 29988 1764 29998
rect 1820 29988 1876 33068
rect 2044 33058 2100 33068
rect 2492 33122 2548 33134
rect 2492 33070 2494 33122
rect 2546 33070 2548 33122
rect 2492 33012 2548 33070
rect 2492 32946 2548 32956
rect 2044 32562 2100 32574
rect 2044 32510 2046 32562
rect 2098 32510 2100 32562
rect 2044 32340 2100 32510
rect 2604 32450 2660 32462
rect 2604 32398 2606 32450
rect 2658 32398 2660 32450
rect 2268 32340 2324 32350
rect 2044 32338 2324 32340
rect 2044 32286 2270 32338
rect 2322 32286 2324 32338
rect 2044 32284 2324 32286
rect 2268 32274 2324 32284
rect 2044 31666 2100 31678
rect 2044 31614 2046 31666
rect 2098 31614 2100 31666
rect 1932 30994 1988 31006
rect 1932 30942 1934 30994
rect 1986 30942 1988 30994
rect 1932 30884 1988 30942
rect 1932 30818 1988 30828
rect 2044 30324 2100 31614
rect 2380 31668 2436 31678
rect 2380 31574 2436 31612
rect 2492 30884 2548 30894
rect 2492 30790 2548 30828
rect 2604 30324 2660 32398
rect 2940 32450 2996 32462
rect 2940 32398 2942 32450
rect 2994 32398 2996 32450
rect 2940 32338 2996 32398
rect 2940 32286 2942 32338
rect 2994 32286 2996 32338
rect 2716 31666 2772 31678
rect 2716 31614 2718 31666
rect 2770 31614 2772 31666
rect 2716 31556 2772 31614
rect 2716 31490 2772 31500
rect 2044 30268 2884 30324
rect 2044 30098 2100 30110
rect 2044 30046 2046 30098
rect 2098 30046 2100 30098
rect 2044 29988 2100 30046
rect 2604 29988 2660 29998
rect 1820 29932 1988 29988
rect 2044 29986 2660 29988
rect 2044 29934 2606 29986
rect 2658 29934 2660 29986
rect 2044 29932 2660 29934
rect 1708 29894 1764 29932
rect 1708 29538 1764 29550
rect 1708 29486 1710 29538
rect 1762 29486 1764 29538
rect 1708 28980 1764 29486
rect 1708 28914 1764 28924
rect 1708 28420 1764 28430
rect 1708 28326 1764 28364
rect 1708 27970 1764 27982
rect 1708 27918 1710 27970
rect 1762 27918 1764 27970
rect 1708 27636 1764 27918
rect 1708 27570 1764 27580
rect 1708 26852 1764 26862
rect 1708 26850 1876 26852
rect 1708 26798 1710 26850
rect 1762 26798 1876 26850
rect 1708 26796 1876 26798
rect 1708 26786 1764 26796
rect 1708 26402 1764 26414
rect 1708 26350 1710 26402
rect 1762 26350 1764 26402
rect 1708 25620 1764 26350
rect 1820 26292 1876 26796
rect 1820 26226 1876 26236
rect 1708 25554 1764 25564
rect 1708 25282 1764 25294
rect 1708 25230 1710 25282
rect 1762 25230 1764 25282
rect 1708 25060 1764 25230
rect 1708 24994 1764 25004
rect 1708 24834 1764 24846
rect 1708 24782 1710 24834
rect 1762 24782 1764 24834
rect 1708 24276 1764 24782
rect 1708 24210 1764 24220
rect 1708 23716 1764 23726
rect 1708 23622 1764 23660
rect 1708 23266 1764 23278
rect 1708 23214 1710 23266
rect 1762 23214 1764 23266
rect 1708 22932 1764 23214
rect 1708 22866 1764 22876
rect 1708 22260 1764 22270
rect 1708 22166 1764 22204
rect 1708 21698 1764 21710
rect 1708 21646 1710 21698
rect 1762 21646 1764 21698
rect 1708 20916 1764 21646
rect 1708 20850 1764 20860
rect 1932 20692 1988 29932
rect 2044 29426 2100 29438
rect 2044 29374 2046 29426
rect 2098 29374 2100 29426
rect 2044 29316 2100 29374
rect 2044 29250 2100 29260
rect 2492 29316 2548 29326
rect 2492 29222 2548 29260
rect 2044 28532 2100 28542
rect 2044 28438 2100 28476
rect 2044 27860 2100 27870
rect 2044 27766 2100 27804
rect 2044 26962 2100 26974
rect 2044 26910 2046 26962
rect 2098 26910 2100 26962
rect 2044 26908 2100 26910
rect 2380 26964 2436 27002
rect 2044 26852 2324 26908
rect 2380 26898 2436 26908
rect 2044 26290 2100 26302
rect 2044 26238 2046 26290
rect 2098 26238 2100 26290
rect 2044 25620 2100 26238
rect 2044 25554 2100 25564
rect 2044 25396 2100 25406
rect 2044 25394 2212 25396
rect 2044 25342 2046 25394
rect 2098 25342 2212 25394
rect 2044 25340 2212 25342
rect 2044 25330 2100 25340
rect 2044 24836 2100 24846
rect 2044 24742 2100 24780
rect 2044 23826 2100 23838
rect 2044 23774 2046 23826
rect 2098 23774 2100 23826
rect 2044 23380 2100 23774
rect 2156 23716 2212 25340
rect 2268 25284 2324 26852
rect 2268 25218 2324 25228
rect 2156 23650 2212 23660
rect 2044 23314 2100 23324
rect 2044 23156 2100 23166
rect 2044 23154 2212 23156
rect 2044 23102 2046 23154
rect 2098 23102 2212 23154
rect 2044 23100 2212 23102
rect 2044 23090 2100 23100
rect 2044 22260 2100 22270
rect 2044 22166 2100 22204
rect 2156 22148 2212 23100
rect 2156 22082 2212 22092
rect 2380 22146 2436 22158
rect 2380 22094 2382 22146
rect 2434 22094 2436 22146
rect 2380 21812 2436 22094
rect 2380 21746 2436 21756
rect 2604 21812 2660 29932
rect 2716 26964 2772 27002
rect 2716 26898 2772 26908
rect 2828 25172 2884 30268
rect 2828 25106 2884 25116
rect 2716 22484 2772 22494
rect 2716 22370 2772 22428
rect 2716 22318 2718 22370
rect 2770 22318 2772 22370
rect 2716 22306 2772 22318
rect 2604 21746 2660 21756
rect 2044 21588 2100 21598
rect 2044 21494 2100 21532
rect 1932 20626 1988 20636
rect 2044 20690 2100 20702
rect 2044 20638 2046 20690
rect 2098 20638 2100 20690
rect 1708 20578 1764 20590
rect 1708 20526 1710 20578
rect 1762 20526 1764 20578
rect 1708 20244 1764 20526
rect 2044 20356 2100 20638
rect 2044 20290 2100 20300
rect 1708 20178 1764 20188
rect 2044 20132 2100 20142
rect 2044 20038 2100 20076
rect 1708 20018 1764 20030
rect 1708 19966 1710 20018
rect 1762 19966 1764 20018
rect 1708 19572 1764 19966
rect 1708 19506 1764 19516
rect 2492 19906 2548 19918
rect 2492 19854 2494 19906
rect 2546 19854 2548 19906
rect 2492 19572 2548 19854
rect 2940 19796 2996 32286
rect 3052 26180 3108 36204
rect 3164 35922 3220 36428
rect 3276 36372 3332 36382
rect 3388 36372 3444 39200
rect 4060 36484 4116 39200
rect 4060 36482 4564 36484
rect 4060 36430 4062 36482
rect 4114 36430 4564 36482
rect 4060 36428 4564 36430
rect 4060 36418 4116 36428
rect 3276 36370 3444 36372
rect 3276 36318 3278 36370
rect 3330 36318 3444 36370
rect 3276 36316 3444 36318
rect 3612 36370 3668 36382
rect 3612 36318 3614 36370
rect 3666 36318 3668 36370
rect 3276 36306 3332 36316
rect 3164 35870 3166 35922
rect 3218 35870 3220 35922
rect 3164 35858 3220 35870
rect 3612 35586 3668 36318
rect 4284 36258 4340 36270
rect 4284 36206 4286 36258
rect 4338 36206 4340 36258
rect 3612 35534 3614 35586
rect 3666 35534 3668 35586
rect 3276 31556 3332 31566
rect 3276 31462 3332 31500
rect 3612 30100 3668 35534
rect 3612 30034 3668 30044
rect 4172 35586 4228 35598
rect 4172 35534 4174 35586
rect 4226 35534 4228 35586
rect 4172 35474 4228 35534
rect 4172 35422 4174 35474
rect 4226 35422 4228 35474
rect 3052 26114 3108 26124
rect 4060 29316 4116 29326
rect 4060 22596 4116 29260
rect 4172 27076 4228 35422
rect 4284 29316 4340 36206
rect 4508 35922 4564 36428
rect 4620 36372 4676 36382
rect 4732 36372 4788 39200
rect 4620 36370 4788 36372
rect 4620 36318 4622 36370
rect 4674 36318 4788 36370
rect 4620 36316 4788 36318
rect 4844 36482 4900 36494
rect 4844 36430 4846 36482
rect 4898 36430 4900 36482
rect 4620 36306 4676 36316
rect 4508 35870 4510 35922
rect 4562 35870 4564 35922
rect 4508 35858 4564 35870
rect 4620 35476 4676 35486
rect 4844 35476 4900 36430
rect 5404 35924 5460 39200
rect 6076 37044 6132 39200
rect 5740 36988 6132 37044
rect 5740 36484 5796 36988
rect 5874 36876 6138 36886
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 5874 36810 6138 36820
rect 6524 36484 6580 36494
rect 6748 36484 6804 39200
rect 5740 36482 5908 36484
rect 5740 36430 5742 36482
rect 5794 36430 5908 36482
rect 5740 36428 5908 36430
rect 5740 36418 5796 36428
rect 5628 35924 5684 35934
rect 5404 35922 5684 35924
rect 5404 35870 5406 35922
rect 5458 35870 5630 35922
rect 5682 35870 5684 35922
rect 5404 35868 5684 35870
rect 5404 35858 5460 35868
rect 5628 35858 5684 35868
rect 5852 35588 5908 36428
rect 6524 36482 7028 36484
rect 6524 36430 6526 36482
rect 6578 36430 7028 36482
rect 6524 36428 7028 36430
rect 6524 36418 6580 36428
rect 6076 36260 6132 36270
rect 6076 36258 6692 36260
rect 6076 36206 6078 36258
rect 6130 36206 6692 36258
rect 6076 36204 6692 36206
rect 6076 36194 6132 36204
rect 5964 35812 6020 35822
rect 5964 35810 6580 35812
rect 5964 35758 5966 35810
rect 6018 35758 6580 35810
rect 5964 35756 6580 35758
rect 5964 35746 6020 35756
rect 6412 35588 6468 35598
rect 5852 35586 6468 35588
rect 5852 35534 6414 35586
rect 6466 35534 6468 35586
rect 5852 35532 6468 35534
rect 6412 35522 6468 35532
rect 4620 35474 4900 35476
rect 4620 35422 4622 35474
rect 4674 35422 4900 35474
rect 4620 35420 4900 35422
rect 4620 35410 4676 35420
rect 5874 35308 6138 35318
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 5874 35242 6138 35252
rect 5874 33740 6138 33750
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 5874 33674 6138 33684
rect 5874 32172 6138 32182
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 5874 32106 6138 32116
rect 5874 30604 6138 30614
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 5874 30538 6138 30548
rect 4284 29250 4340 29260
rect 5874 29036 6138 29046
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 5874 28970 6138 28980
rect 5874 27468 6138 27478
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 5874 27402 6138 27412
rect 4172 27010 4228 27020
rect 5874 25900 6138 25910
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 5874 25834 6138 25844
rect 5068 25172 5124 25182
rect 5068 23268 5124 25116
rect 6524 25172 6580 35756
rect 6636 29540 6692 36204
rect 6636 29474 6692 29484
rect 6748 36258 6804 36270
rect 6748 36206 6750 36258
rect 6802 36206 6804 36258
rect 6748 29428 6804 36206
rect 6972 35922 7028 36428
rect 6972 35870 6974 35922
rect 7026 35870 7028 35922
rect 6972 35858 7028 35870
rect 7084 36370 7140 36382
rect 7084 36318 7086 36370
rect 7138 36318 7140 36370
rect 6748 29362 6804 29372
rect 6860 30884 6916 30894
rect 6524 25106 6580 25116
rect 6748 26964 6804 26974
rect 5874 24332 6138 24342
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 5874 24266 6138 24276
rect 5068 23202 5124 23212
rect 5874 22764 6138 22774
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 5874 22698 6138 22708
rect 4060 22530 4116 22540
rect 6748 22372 6804 26908
rect 6748 22306 6804 22316
rect 6860 21700 6916 30828
rect 7084 26516 7140 36318
rect 7420 36370 7476 39200
rect 7420 36318 7422 36370
rect 7474 36318 7476 36370
rect 7420 36306 7476 36318
rect 7868 36482 7924 36494
rect 7868 36430 7870 36482
rect 7922 36430 7924 36482
rect 7868 30212 7924 36430
rect 8092 36370 8148 39200
rect 8092 36318 8094 36370
rect 8146 36318 8148 36370
rect 8092 36306 8148 36318
rect 8428 36370 8484 36382
rect 8428 36318 8430 36370
rect 8482 36318 8484 36370
rect 7868 30146 7924 30156
rect 8428 27972 8484 36318
rect 8764 36370 8820 39200
rect 8764 36318 8766 36370
rect 8818 36318 8820 36370
rect 8764 36306 8820 36318
rect 9100 35924 9156 35934
rect 9436 35924 9492 39200
rect 9660 36484 9716 36494
rect 9660 36482 9828 36484
rect 9660 36430 9662 36482
rect 9714 36430 9828 36482
rect 9660 36428 9828 36430
rect 9660 36418 9716 36428
rect 9660 35924 9716 35934
rect 9100 35922 9716 35924
rect 9100 35870 9102 35922
rect 9154 35870 9662 35922
rect 9714 35870 9716 35922
rect 9100 35868 9716 35870
rect 9100 35858 9156 35868
rect 9660 35858 9716 35868
rect 9772 35588 9828 36428
rect 9884 36372 9940 36382
rect 10108 36372 10164 39200
rect 9884 36370 10164 36372
rect 9884 36318 9886 36370
rect 9938 36318 10164 36370
rect 9884 36316 10164 36318
rect 10332 36482 10388 36494
rect 10332 36430 10334 36482
rect 10386 36430 10388 36482
rect 9884 36306 9940 36316
rect 9996 35812 10052 35822
rect 9996 35718 10052 35756
rect 9772 35522 9828 35532
rect 10332 33796 10388 36430
rect 10556 36372 10612 36382
rect 10780 36372 10836 39200
rect 11004 36484 11060 36494
rect 11004 36482 11172 36484
rect 11004 36430 11006 36482
rect 11058 36430 11172 36482
rect 11004 36428 11172 36430
rect 11004 36418 11060 36428
rect 10556 36370 10836 36372
rect 10556 36318 10558 36370
rect 10610 36318 10836 36370
rect 10556 36316 10836 36318
rect 10556 36306 10612 36316
rect 10536 36092 10800 36102
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10536 36026 10800 36036
rect 10444 35588 10500 35598
rect 10444 35494 10500 35532
rect 10536 34524 10800 34534
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10536 34458 10800 34468
rect 10332 33730 10388 33740
rect 10536 32956 10800 32966
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10536 32890 10800 32900
rect 11116 32340 11172 36428
rect 11228 36372 11284 36382
rect 11452 36372 11508 39200
rect 11228 36370 11508 36372
rect 11228 36318 11230 36370
rect 11282 36318 11508 36370
rect 11228 36316 11508 36318
rect 11676 36482 11732 36494
rect 11676 36430 11678 36482
rect 11730 36430 11732 36482
rect 11228 36306 11284 36316
rect 11676 33684 11732 36430
rect 11900 36372 11956 36382
rect 12124 36372 12180 39200
rect 12796 37716 12852 39200
rect 12572 37660 12852 37716
rect 11900 36370 12180 36372
rect 11900 36318 11902 36370
rect 11954 36318 12180 36370
rect 11900 36316 12180 36318
rect 12236 36370 12292 36382
rect 12236 36318 12238 36370
rect 12290 36318 12292 36370
rect 11900 36306 11956 36316
rect 11676 33618 11732 33628
rect 11116 32284 11508 32340
rect 8428 27906 8484 27916
rect 9324 31556 9380 31566
rect 7084 26450 7140 26460
rect 6860 21634 6916 21644
rect 6972 25172 7028 25182
rect 6972 21476 7028 25116
rect 9212 22260 9268 22270
rect 9212 22166 9268 22204
rect 6972 21410 7028 21420
rect 5874 21196 6138 21206
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 5874 21130 6138 21140
rect 9324 21140 9380 31500
rect 10536 31388 10800 31398
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10536 31322 10800 31332
rect 10108 30100 10164 30110
rect 9436 27860 9492 27870
rect 9436 26962 9492 27804
rect 10108 27412 10164 30044
rect 10536 29820 10800 29830
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10536 29754 10800 29764
rect 11452 28530 11508 32284
rect 11452 28478 11454 28530
rect 11506 28478 11508 28530
rect 11452 28466 11508 28478
rect 11564 30212 11620 30222
rect 11564 28420 11620 30156
rect 12236 30100 12292 36318
rect 12572 36370 12628 37660
rect 12572 36318 12574 36370
rect 12626 36318 12628 36370
rect 12572 36306 12628 36318
rect 13356 36372 13412 36382
rect 13468 36372 13524 39200
rect 13356 36370 13524 36372
rect 13356 36318 13358 36370
rect 13410 36318 13524 36370
rect 13356 36316 13524 36318
rect 13692 36372 13748 36382
rect 14028 36372 14084 36382
rect 14140 36372 14196 39200
rect 14812 36484 14868 39200
rect 15484 37044 15540 39200
rect 15484 36988 15652 37044
rect 15198 36876 15462 36886
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15198 36810 15462 36820
rect 15484 36484 15540 36494
rect 15596 36484 15652 36988
rect 14812 36482 15316 36484
rect 14812 36430 14814 36482
rect 14866 36430 15316 36482
rect 14812 36428 15316 36430
rect 14812 36418 14868 36428
rect 13692 36370 13860 36372
rect 13692 36318 13694 36370
rect 13746 36318 13860 36370
rect 13692 36316 13860 36318
rect 13356 36306 13412 36316
rect 13692 36306 13748 36316
rect 12236 30034 12292 30044
rect 13692 33684 13748 33694
rect 13692 30098 13748 33628
rect 13692 30046 13694 30098
rect 13746 30046 13748 30098
rect 13692 30034 13748 30046
rect 13244 29426 13300 29438
rect 13244 29374 13246 29426
rect 13298 29374 13300 29426
rect 12684 28756 12740 28766
rect 11564 28354 11620 28364
rect 11788 28530 11844 28542
rect 11788 28478 11790 28530
rect 11842 28478 11844 28530
rect 10536 28252 10800 28262
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10536 28186 10800 28196
rect 10108 27346 10164 27356
rect 11228 27804 11508 27860
rect 10444 27300 10500 27310
rect 10444 27206 10500 27244
rect 10668 27300 10724 27310
rect 11228 27300 11284 27804
rect 10668 27298 11284 27300
rect 10668 27246 10670 27298
rect 10722 27246 11284 27298
rect 10668 27244 11284 27246
rect 10668 27234 10724 27244
rect 10220 27076 10276 27086
rect 10220 27074 10388 27076
rect 10220 27022 10222 27074
rect 10274 27022 10388 27074
rect 10220 27020 10388 27022
rect 10220 27010 10276 27020
rect 9436 26910 9438 26962
rect 9490 26910 9492 26962
rect 9436 26898 9492 26910
rect 9772 26964 9828 26974
rect 10108 26964 10164 26974
rect 9772 26962 10164 26964
rect 9772 26910 9774 26962
rect 9826 26910 10110 26962
rect 10162 26910 10164 26962
rect 9772 26908 10164 26910
rect 9772 26898 9828 26908
rect 10108 26898 10164 26908
rect 10220 26852 10276 26862
rect 10108 26516 10164 26526
rect 10220 26516 10276 26796
rect 10108 26514 10276 26516
rect 10108 26462 10110 26514
rect 10162 26462 10276 26514
rect 10108 26460 10276 26462
rect 10108 26450 10164 26460
rect 9660 26292 9716 26302
rect 9660 24722 9716 26236
rect 9660 24670 9662 24722
rect 9714 24670 9716 24722
rect 9660 24658 9716 24670
rect 9772 26290 9828 26302
rect 9772 26238 9774 26290
rect 9826 26238 9828 26290
rect 9772 25732 9828 26238
rect 9772 24500 9828 25676
rect 10332 24948 10388 27020
rect 10892 27074 10948 27086
rect 10892 27022 10894 27074
rect 10946 27022 10948 27074
rect 10892 26908 10948 27022
rect 11228 27074 11284 27244
rect 11228 27022 11230 27074
rect 11282 27022 11284 27074
rect 11228 27010 11284 27022
rect 11340 27634 11396 27646
rect 11340 27582 11342 27634
rect 11394 27582 11396 27634
rect 11340 26962 11396 27582
rect 11452 27636 11508 27804
rect 11676 27636 11732 27646
rect 11452 27634 11620 27636
rect 11452 27582 11454 27634
rect 11506 27582 11620 27634
rect 11452 27580 11620 27582
rect 11452 27570 11508 27580
rect 11340 26910 11342 26962
rect 11394 26910 11396 26962
rect 11340 26908 11396 26910
rect 10892 26852 11396 26908
rect 10892 26786 10948 26796
rect 10536 26684 10800 26694
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10536 26618 10800 26628
rect 10444 26402 10500 26414
rect 10444 26350 10446 26402
rect 10498 26350 10500 26402
rect 10444 26068 10500 26350
rect 10668 26292 10724 26302
rect 10668 26198 10724 26236
rect 11116 26290 11172 26852
rect 11564 26404 11620 27580
rect 11676 27542 11732 27580
rect 11788 27300 11844 28478
rect 12348 28532 12404 28542
rect 12348 28082 12404 28476
rect 12348 28030 12350 28082
rect 12402 28030 12404 28082
rect 12348 28018 12404 28030
rect 12572 27858 12628 27870
rect 12572 27806 12574 27858
rect 12626 27806 12628 27858
rect 12012 27748 12068 27758
rect 12572 27748 12628 27806
rect 12012 27746 12628 27748
rect 12012 27694 12014 27746
rect 12066 27694 12628 27746
rect 12012 27692 12628 27694
rect 12012 27682 12068 27692
rect 11676 27244 11844 27300
rect 11900 27634 11956 27646
rect 11900 27582 11902 27634
rect 11954 27582 11956 27634
rect 11676 26908 11732 27244
rect 11900 27076 11956 27582
rect 12348 27076 12404 27086
rect 12684 27076 12740 28700
rect 13132 28644 13188 28654
rect 13244 28644 13300 29374
rect 13188 28588 13300 28644
rect 13468 29202 13524 29214
rect 13468 29150 13470 29202
rect 13522 29150 13524 29202
rect 13132 27860 13188 28588
rect 11900 27020 12068 27076
rect 11676 26852 11956 26908
rect 11900 26850 11956 26852
rect 11900 26798 11902 26850
rect 11954 26798 11956 26850
rect 11900 26786 11956 26798
rect 11340 26348 11620 26404
rect 11676 26514 11732 26526
rect 11676 26462 11678 26514
rect 11730 26462 11732 26514
rect 11340 26292 11396 26348
rect 11116 26238 11118 26290
rect 11170 26238 11172 26290
rect 11116 26226 11172 26238
rect 11228 26290 11396 26292
rect 11228 26238 11342 26290
rect 11394 26238 11396 26290
rect 11228 26236 11396 26238
rect 11228 26068 11284 26236
rect 11340 26226 11396 26236
rect 11564 26180 11620 26190
rect 11564 26086 11620 26124
rect 10444 26012 11284 26068
rect 11564 25508 11620 25518
rect 11452 25284 11508 25294
rect 11452 25190 11508 25228
rect 10536 25116 10800 25126
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10536 25050 10800 25060
rect 10332 24892 10724 24948
rect 9884 24836 9940 24846
rect 10220 24836 10276 24846
rect 9884 24834 10164 24836
rect 9884 24782 9886 24834
rect 9938 24782 10164 24834
rect 9884 24780 10164 24782
rect 9884 24770 9940 24780
rect 9548 24444 9828 24500
rect 9436 23940 9492 23950
rect 9548 23940 9604 24444
rect 10108 24164 10164 24780
rect 10220 24742 10276 24780
rect 10220 24164 10276 24174
rect 10108 24162 10276 24164
rect 10108 24110 10222 24162
rect 10274 24110 10276 24162
rect 10108 24108 10276 24110
rect 9996 23940 10052 23950
rect 9436 23938 9604 23940
rect 9436 23886 9438 23938
rect 9490 23886 9604 23938
rect 9436 23884 9604 23886
rect 9660 23938 10052 23940
rect 9660 23886 9998 23938
rect 10050 23886 10052 23938
rect 9660 23884 10052 23886
rect 9436 23874 9492 23884
rect 9660 23826 9716 23884
rect 9660 23774 9662 23826
rect 9714 23774 9716 23826
rect 9660 23762 9716 23774
rect 9996 22594 10052 23884
rect 10108 23380 10164 23390
rect 10108 23286 10164 23324
rect 9996 22542 9998 22594
rect 10050 22542 10052 22594
rect 9548 22260 9604 22270
rect 9548 22258 9940 22260
rect 9548 22206 9550 22258
rect 9602 22206 9940 22258
rect 9548 22204 9940 22206
rect 9548 22194 9604 22204
rect 9884 21812 9940 22204
rect 9996 22036 10052 22542
rect 10108 22596 10164 22606
rect 10220 22596 10276 24108
rect 10332 23380 10388 24892
rect 10556 24722 10612 24734
rect 10556 24670 10558 24722
rect 10610 24670 10612 24722
rect 10444 23940 10500 23950
rect 10444 23846 10500 23884
rect 10556 23714 10612 24670
rect 10668 24162 10724 24892
rect 11452 24724 11508 24734
rect 10668 24110 10670 24162
rect 10722 24110 10724 24162
rect 10668 24098 10724 24110
rect 11340 24722 11508 24724
rect 11340 24670 11454 24722
rect 11506 24670 11508 24722
rect 11340 24668 11508 24670
rect 10556 23662 10558 23714
rect 10610 23662 10612 23714
rect 10556 23650 10612 23662
rect 10536 23548 10800 23558
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10536 23482 10800 23492
rect 11116 23380 11172 23390
rect 10332 23324 10612 23380
rect 10108 22594 10276 22596
rect 10108 22542 10110 22594
rect 10162 22542 10276 22594
rect 10108 22540 10276 22542
rect 10108 22530 10164 22540
rect 9996 21980 10164 22036
rect 9996 21812 10052 21822
rect 9884 21810 10052 21812
rect 9884 21758 9998 21810
rect 10050 21758 10052 21810
rect 9884 21756 10052 21758
rect 9996 21746 10052 21756
rect 9324 21074 9380 21084
rect 9996 21588 10052 21598
rect 10108 21588 10164 21980
rect 9996 21586 10164 21588
rect 9996 21534 9998 21586
rect 10050 21534 10164 21586
rect 9996 21532 10164 21534
rect 9996 21026 10052 21532
rect 9996 20974 9998 21026
rect 10050 20974 10052 21026
rect 9996 20962 10052 20974
rect 10108 21364 10164 21374
rect 10220 21364 10276 22540
rect 10444 23154 10500 23166
rect 10444 23102 10446 23154
rect 10498 23102 10500 23154
rect 10332 22370 10388 22382
rect 10332 22318 10334 22370
rect 10386 22318 10388 22370
rect 10332 22260 10388 22318
rect 10332 22194 10388 22204
rect 10444 22146 10500 23102
rect 10556 22596 10612 23324
rect 10556 22594 10948 22596
rect 10556 22542 10558 22594
rect 10610 22542 10948 22594
rect 10556 22540 10948 22542
rect 10556 22530 10612 22540
rect 10444 22094 10446 22146
rect 10498 22094 10500 22146
rect 10444 22082 10500 22094
rect 10536 21980 10800 21990
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10536 21914 10800 21924
rect 10892 21812 10948 22540
rect 10556 21756 10948 21812
rect 11116 21812 11172 23324
rect 11228 22148 11284 22158
rect 11228 22054 11284 22092
rect 11340 21924 11396 24668
rect 11452 24658 11508 24668
rect 11564 23938 11620 25452
rect 11676 25506 11732 26462
rect 11676 25454 11678 25506
rect 11730 25454 11732 25506
rect 11676 25442 11732 25454
rect 11788 26068 11844 26078
rect 12012 26068 12068 27020
rect 12348 27074 12740 27076
rect 12348 27022 12350 27074
rect 12402 27022 12740 27074
rect 12348 27020 12740 27022
rect 12908 27858 13188 27860
rect 12908 27806 13134 27858
rect 13186 27806 13188 27858
rect 12908 27804 13188 27806
rect 12348 27010 12404 27020
rect 12796 26962 12852 26974
rect 12796 26910 12798 26962
rect 12850 26910 12852 26962
rect 12796 26908 12852 26910
rect 11788 26066 12068 26068
rect 11788 26014 11790 26066
rect 11842 26014 12068 26066
rect 11788 26012 12068 26014
rect 12572 26852 12852 26908
rect 11676 24836 11732 24846
rect 11788 24836 11844 26012
rect 12460 25394 12516 25406
rect 12460 25342 12462 25394
rect 12514 25342 12516 25394
rect 12460 25172 12516 25342
rect 11676 24834 11844 24836
rect 11676 24782 11678 24834
rect 11730 24782 11844 24834
rect 11676 24780 11844 24782
rect 12012 24836 12068 24846
rect 12348 24836 12404 24846
rect 12460 24836 12516 25116
rect 12012 24834 12180 24836
rect 12012 24782 12014 24834
rect 12066 24782 12180 24834
rect 12012 24780 12180 24782
rect 11676 24724 11732 24780
rect 12012 24770 12068 24780
rect 11676 24658 11732 24668
rect 11564 23886 11566 23938
rect 11618 23886 11620 23938
rect 11564 23874 11620 23886
rect 11788 24052 11844 24062
rect 11788 23826 11844 23996
rect 12124 23940 12180 24780
rect 12348 24834 12516 24836
rect 12348 24782 12350 24834
rect 12402 24782 12516 24834
rect 12348 24780 12516 24782
rect 12348 24770 12404 24780
rect 12572 24724 12628 26852
rect 12684 26290 12740 26302
rect 12684 26238 12686 26290
rect 12738 26238 12740 26290
rect 12684 25508 12740 26238
rect 12684 25442 12740 25452
rect 12796 25396 12852 25406
rect 12908 25396 12964 27804
rect 13132 27794 13188 27804
rect 13468 28084 13524 29150
rect 13692 29204 13748 29214
rect 13692 29110 13748 29148
rect 13580 28644 13636 28654
rect 13580 28550 13636 28588
rect 13692 28642 13748 28654
rect 13692 28590 13694 28642
rect 13746 28590 13748 28642
rect 13692 28084 13748 28590
rect 13804 28644 13860 36316
rect 14028 36370 14196 36372
rect 14028 36318 14030 36370
rect 14082 36318 14196 36370
rect 14028 36316 14196 36318
rect 14364 36370 14420 36382
rect 14364 36318 14366 36370
rect 14418 36318 14420 36370
rect 14028 36306 14084 36316
rect 14140 33796 14196 33806
rect 14196 33740 14308 33796
rect 14140 33730 14196 33740
rect 14028 30098 14084 30110
rect 14028 30046 14030 30098
rect 14082 30046 14084 30098
rect 14028 29538 14084 30046
rect 14252 29652 14308 33740
rect 14364 30212 14420 36318
rect 15036 36260 15092 36270
rect 14364 30146 14420 30156
rect 14700 36258 15092 36260
rect 14700 36206 15038 36258
rect 15090 36206 15092 36258
rect 14700 36204 15092 36206
rect 14364 29652 14420 29662
rect 14252 29650 14420 29652
rect 14252 29598 14366 29650
rect 14418 29598 14420 29650
rect 14252 29596 14420 29598
rect 14364 29586 14420 29596
rect 14028 29486 14030 29538
rect 14082 29486 14084 29538
rect 14028 29474 14084 29486
rect 14588 29428 14644 29438
rect 14476 29426 14644 29428
rect 14476 29374 14590 29426
rect 14642 29374 14644 29426
rect 14476 29372 14644 29374
rect 13916 29204 13972 29214
rect 13916 29202 14084 29204
rect 13916 29150 13918 29202
rect 13970 29150 14084 29202
rect 13916 29148 14084 29150
rect 13916 29138 13972 29148
rect 13916 28756 13972 28766
rect 13916 28662 13972 28700
rect 14028 28644 14084 29148
rect 14252 28868 14308 28878
rect 14476 28868 14532 29372
rect 14588 29362 14644 29372
rect 14700 29204 14756 36204
rect 15036 36194 15092 36204
rect 15260 35922 15316 36428
rect 15484 36482 15988 36484
rect 15484 36430 15486 36482
rect 15538 36430 15988 36482
rect 15484 36428 15988 36430
rect 15484 36418 15540 36428
rect 15260 35870 15262 35922
rect 15314 35870 15316 35922
rect 15260 35858 15316 35870
rect 15708 36258 15764 36270
rect 15708 36206 15710 36258
rect 15762 36206 15764 36258
rect 15198 35308 15462 35318
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15198 35242 15462 35252
rect 15198 33740 15462 33750
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15198 33674 15462 33684
rect 15198 32172 15462 32182
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15198 32106 15462 32116
rect 15198 30604 15462 30614
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15198 30538 15462 30548
rect 15596 30212 15652 30222
rect 14812 30100 14868 30110
rect 14868 30044 14980 30100
rect 14812 30034 14868 30044
rect 14252 28866 14532 28868
rect 14252 28814 14254 28866
rect 14306 28814 14532 28866
rect 14252 28812 14532 28814
rect 14588 29148 14756 29204
rect 14252 28802 14308 28812
rect 14140 28644 14196 28654
rect 14028 28642 14196 28644
rect 14028 28590 14142 28642
rect 14194 28590 14196 28642
rect 14028 28588 14196 28590
rect 13804 28578 13860 28588
rect 14140 28084 14196 28588
rect 13468 28028 13748 28084
rect 13804 28028 14196 28084
rect 14252 28644 14308 28654
rect 13356 27636 13412 27646
rect 13468 27636 13524 28028
rect 13356 27634 13524 27636
rect 13356 27582 13358 27634
rect 13410 27582 13524 27634
rect 13356 27580 13524 27582
rect 13356 27570 13412 27580
rect 13020 26516 13076 26526
rect 13468 26516 13524 27580
rect 13580 27636 13636 27646
rect 13580 27542 13636 27580
rect 13804 27634 13860 28028
rect 13804 27582 13806 27634
rect 13858 27582 13860 27634
rect 13580 27412 13636 27422
rect 13580 26962 13636 27356
rect 13580 26910 13582 26962
rect 13634 26910 13636 26962
rect 13580 26898 13636 26910
rect 13020 26514 13524 26516
rect 13020 26462 13022 26514
rect 13074 26462 13524 26514
rect 13020 26460 13524 26462
rect 13020 26450 13076 26460
rect 13468 26292 13524 26460
rect 13804 26404 13860 27582
rect 13916 27634 13972 27646
rect 13916 27582 13918 27634
rect 13970 27582 13972 27634
rect 13916 27074 13972 27582
rect 13916 27022 13918 27074
rect 13970 27022 13972 27074
rect 13916 27010 13972 27022
rect 13692 26348 13860 26404
rect 13580 26292 13636 26302
rect 13468 26290 13636 26292
rect 13468 26238 13582 26290
rect 13634 26238 13636 26290
rect 13468 26236 13636 26238
rect 13580 26226 13636 26236
rect 13468 26066 13524 26078
rect 13468 26014 13470 26066
rect 13522 26014 13524 26066
rect 12852 25340 12964 25396
rect 13020 25620 13076 25630
rect 12796 25302 12852 25340
rect 13020 24946 13076 25564
rect 13356 25396 13412 25406
rect 13468 25396 13524 26014
rect 13412 25340 13524 25396
rect 13356 25330 13412 25340
rect 13692 25172 13748 26348
rect 14140 26292 14196 26302
rect 14140 26198 14196 26236
rect 13804 26180 13860 26190
rect 13804 26086 13860 26124
rect 14028 26066 14084 26078
rect 14028 26014 14030 26066
rect 14082 26014 14084 26066
rect 14028 25620 14084 26014
rect 14028 25554 14084 25564
rect 14252 25284 14308 28588
rect 14476 26516 14532 26526
rect 14476 26422 14532 26460
rect 14476 25620 14532 25630
rect 14364 25284 14420 25294
rect 14252 25228 14364 25284
rect 14364 25218 14420 25228
rect 13020 24894 13022 24946
rect 13074 24894 13076 24946
rect 13020 24882 13076 24894
rect 13244 25116 13748 25172
rect 12572 24658 12628 24668
rect 12348 24052 12404 24062
rect 12348 23958 12404 23996
rect 12572 23940 12628 23950
rect 11788 23774 11790 23826
rect 11842 23774 11844 23826
rect 11788 23548 11844 23774
rect 11900 23938 12180 23940
rect 11900 23886 12126 23938
rect 12178 23886 12180 23938
rect 11900 23884 12180 23886
rect 11900 23716 11956 23884
rect 12124 23874 12180 23884
rect 12460 23884 12572 23940
rect 11900 23660 12180 23716
rect 11788 23492 11956 23548
rect 11900 22372 11956 23492
rect 12012 22596 12068 22606
rect 12124 22596 12180 23660
rect 12236 23268 12292 23278
rect 12236 23174 12292 23212
rect 12012 22594 12292 22596
rect 12012 22542 12014 22594
rect 12066 22542 12292 22594
rect 12012 22540 12292 22542
rect 12012 22530 12068 22540
rect 12124 22372 12180 22382
rect 11900 22370 12180 22372
rect 11900 22318 12126 22370
rect 12178 22318 12180 22370
rect 11900 22316 12180 22318
rect 11564 22258 11620 22270
rect 11564 22206 11566 22258
rect 11618 22206 11620 22258
rect 11564 22148 11620 22206
rect 12012 22148 12068 22158
rect 11564 22146 12068 22148
rect 11564 22094 12014 22146
rect 12066 22094 12068 22146
rect 11564 22092 12068 22094
rect 12012 22082 12068 22092
rect 12124 22148 12180 22316
rect 12124 22082 12180 22092
rect 11340 21868 11732 21924
rect 11116 21756 11396 21812
rect 10556 21588 10612 21756
rect 11004 21700 11060 21710
rect 11004 21606 11060 21644
rect 11228 21588 11284 21598
rect 10444 21586 10612 21588
rect 10444 21534 10558 21586
rect 10610 21534 10612 21586
rect 10444 21532 10612 21534
rect 10108 21362 10276 21364
rect 10108 21310 10110 21362
rect 10162 21310 10276 21362
rect 10108 21308 10276 21310
rect 10332 21364 10388 21374
rect 10108 21026 10164 21308
rect 10332 21270 10388 21308
rect 10108 20974 10110 21026
rect 10162 20974 10164 21026
rect 10108 20962 10164 20974
rect 10332 20916 10388 20926
rect 10332 20822 10388 20860
rect 10444 20580 10500 21532
rect 10556 21522 10612 21532
rect 11116 21586 11284 21588
rect 11116 21534 11230 21586
rect 11282 21534 11284 21586
rect 11116 21532 11284 21534
rect 11116 21140 11172 21532
rect 11228 21522 11284 21532
rect 11340 21364 11396 21756
rect 10668 21084 11172 21140
rect 11228 21308 11396 21364
rect 10668 21026 10724 21084
rect 10668 20974 10670 21026
rect 10722 20974 10724 21026
rect 10668 20962 10724 20974
rect 10556 20804 10612 20814
rect 10556 20802 11060 20804
rect 10556 20750 10558 20802
rect 10610 20750 11060 20802
rect 10556 20748 11060 20750
rect 10556 20738 10612 20748
rect 10332 20524 10500 20580
rect 10332 20244 10388 20524
rect 10536 20412 10800 20422
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10536 20346 10800 20356
rect 10556 20244 10612 20254
rect 10332 20242 10612 20244
rect 10332 20190 10558 20242
rect 10610 20190 10612 20242
rect 10332 20188 10612 20190
rect 10556 20178 10612 20188
rect 9884 20130 9940 20142
rect 9884 20078 9886 20130
rect 9938 20078 9940 20130
rect 2940 19730 2996 19740
rect 9660 20018 9716 20030
rect 9660 19966 9662 20018
rect 9714 19966 9716 20018
rect 5874 19628 6138 19638
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 5874 19562 6138 19572
rect 9660 19572 9716 19966
rect 9884 20020 9940 20078
rect 10332 20020 10388 20030
rect 9884 20018 10388 20020
rect 9884 19966 10334 20018
rect 10386 19966 10388 20018
rect 9884 19964 10388 19966
rect 2492 19506 2548 19516
rect 9660 19506 9716 19516
rect 10332 19348 10388 19964
rect 10556 19348 10612 19358
rect 10892 19348 10948 20748
rect 11004 20690 11060 20748
rect 11004 20638 11006 20690
rect 11058 20638 11060 20690
rect 11004 20626 11060 20638
rect 11228 20188 11284 21308
rect 10332 19292 10556 19348
rect 10556 19234 10612 19292
rect 10556 19182 10558 19234
rect 10610 19182 10612 19234
rect 10556 19170 10612 19182
rect 10668 19292 10948 19348
rect 11004 20132 11284 20188
rect 11340 20690 11396 20702
rect 11340 20638 11342 20690
rect 11394 20638 11396 20690
rect 11340 20188 11396 20638
rect 11676 20188 11732 21868
rect 12236 21812 12292 22540
rect 12348 22370 12404 22382
rect 12348 22318 12350 22370
rect 12402 22318 12404 22370
rect 12348 22260 12404 22318
rect 12348 21924 12404 22204
rect 12460 22036 12516 23884
rect 12572 23846 12628 23884
rect 12796 23940 12852 23950
rect 12796 23846 12852 23884
rect 13244 23940 13300 25116
rect 13356 24724 13412 24734
rect 13692 24724 13748 24734
rect 13356 24722 13748 24724
rect 13356 24670 13358 24722
rect 13410 24670 13694 24722
rect 13746 24670 13748 24722
rect 13356 24668 13748 24670
rect 13356 24658 13412 24668
rect 13692 24658 13748 24668
rect 13804 24724 13860 24734
rect 14252 24724 14308 24734
rect 13804 24630 13860 24668
rect 13916 24668 14252 24724
rect 13244 23874 13300 23884
rect 13804 23940 13860 23950
rect 12684 23716 12740 23726
rect 12572 23714 12740 23716
rect 12572 23662 12686 23714
rect 12738 23662 12740 23714
rect 12572 23660 12740 23662
rect 12572 23266 12628 23660
rect 12684 23650 12740 23660
rect 12572 23214 12574 23266
rect 12626 23214 12628 23266
rect 12572 23202 12628 23214
rect 13692 23156 13748 23166
rect 13692 23062 13748 23100
rect 13468 22932 13524 22942
rect 13804 22932 13860 23884
rect 13916 23154 13972 24668
rect 14252 24630 14308 24668
rect 14364 24612 14420 24622
rect 14028 24500 14084 24510
rect 14028 24406 14084 24444
rect 14364 24498 14420 24556
rect 14364 24446 14366 24498
rect 14418 24446 14420 24498
rect 14364 24276 14420 24446
rect 14140 24220 14420 24276
rect 13916 23102 13918 23154
rect 13970 23102 13972 23154
rect 13916 23090 13972 23102
rect 14028 23378 14084 23390
rect 14028 23326 14030 23378
rect 14082 23326 14084 23378
rect 13468 22930 13636 22932
rect 13468 22878 13470 22930
rect 13522 22878 13636 22930
rect 13468 22876 13636 22878
rect 13804 22876 13972 22932
rect 13468 22866 13524 22876
rect 12572 22372 12628 22382
rect 12572 22370 12852 22372
rect 12572 22318 12574 22370
rect 12626 22318 12852 22370
rect 12572 22316 12852 22318
rect 12572 22306 12628 22316
rect 12460 21970 12516 21980
rect 12572 22148 12628 22158
rect 12348 21858 12404 21868
rect 12012 21756 12292 21812
rect 12012 21588 12068 21756
rect 12348 21588 12404 21598
rect 12572 21588 12628 22092
rect 12012 21532 12180 21588
rect 12124 21476 12180 21532
rect 12348 21586 12628 21588
rect 12348 21534 12350 21586
rect 12402 21534 12628 21586
rect 12348 21532 12628 21534
rect 12796 21586 12852 22316
rect 13468 22148 13524 22158
rect 13244 21812 13300 21822
rect 13468 21812 13524 22092
rect 13244 21718 13300 21756
rect 13356 21756 13524 21812
rect 12796 21534 12798 21586
rect 12850 21534 12852 21586
rect 12236 21476 12292 21486
rect 12124 21474 12292 21476
rect 12124 21422 12238 21474
rect 12290 21422 12292 21474
rect 12124 21420 12292 21422
rect 12236 21026 12292 21420
rect 12236 20974 12238 21026
rect 12290 20974 12292 21026
rect 12236 20962 12292 20974
rect 12348 21026 12404 21532
rect 12572 21364 12628 21374
rect 12572 21270 12628 21308
rect 12348 20974 12350 21026
rect 12402 20974 12404 21026
rect 12348 20962 12404 20974
rect 12796 21026 12852 21534
rect 12908 21588 12964 21598
rect 12908 21494 12964 21532
rect 12796 20974 12798 21026
rect 12850 20974 12852 21026
rect 12572 20916 12628 20926
rect 12572 20822 12628 20860
rect 12796 20356 12852 20974
rect 13244 21364 13300 21374
rect 13356 21364 13412 21756
rect 13468 21588 13524 21598
rect 13468 21494 13524 21532
rect 13356 21308 13524 21364
rect 12236 20300 12852 20356
rect 12236 20242 12292 20300
rect 12236 20190 12238 20242
rect 12290 20190 12292 20242
rect 11340 20132 11508 20188
rect 1708 19010 1764 19022
rect 1708 18958 1710 19010
rect 1762 18958 1764 19010
rect 1708 18900 1764 18958
rect 2044 19012 2100 19022
rect 2044 18918 2100 18956
rect 2492 19010 2548 19022
rect 10668 19012 10724 19292
rect 11004 19236 11060 20132
rect 11228 20018 11284 20030
rect 11228 19966 11230 20018
rect 11282 19966 11284 20018
rect 11228 19572 11284 19966
rect 11228 19506 11284 19516
rect 11452 19348 11508 20132
rect 11564 20132 12068 20188
rect 12236 20178 12292 20190
rect 11564 20130 11620 20132
rect 11564 20078 11566 20130
rect 11618 20078 11620 20130
rect 11564 20066 11620 20078
rect 12012 20020 12068 20132
rect 12012 19926 12068 19964
rect 12572 20130 12628 20142
rect 12572 20078 12574 20130
rect 12626 20078 12628 20130
rect 12572 19796 12628 20078
rect 12572 19730 12628 19740
rect 12684 20020 12740 20030
rect 10780 19180 11396 19236
rect 10780 19122 10836 19180
rect 10780 19070 10782 19122
rect 10834 19070 10836 19122
rect 10780 19058 10836 19070
rect 2492 18958 2494 19010
rect 2546 18958 2548 19010
rect 1708 18834 1764 18844
rect 2492 18900 2548 18958
rect 2492 18834 2548 18844
rect 10332 18956 10724 19012
rect 11116 19012 11172 19022
rect 11116 19010 11284 19012
rect 11116 18958 11118 19010
rect 11170 18958 11284 19010
rect 11116 18956 11284 18958
rect 1708 18562 1764 18574
rect 1708 18510 1710 18562
rect 1762 18510 1764 18562
rect 1708 18228 1764 18510
rect 2044 18452 2100 18462
rect 10332 18452 10388 18956
rect 11116 18946 11172 18956
rect 10536 18844 10800 18854
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10536 18778 10800 18788
rect 10892 18562 10948 18574
rect 10892 18510 10894 18562
rect 10946 18510 10948 18562
rect 10444 18452 10500 18462
rect 10332 18450 10724 18452
rect 10332 18398 10446 18450
rect 10498 18398 10724 18450
rect 10332 18396 10724 18398
rect 2044 18358 2100 18396
rect 10444 18386 10500 18396
rect 1708 18162 1764 18172
rect 8764 18228 8820 18238
rect 5874 18060 6138 18070
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 5874 17994 6138 18004
rect 2716 17780 2772 17790
rect 2716 17666 2772 17724
rect 2716 17614 2718 17666
rect 2770 17614 2772 17666
rect 2716 17602 2772 17614
rect 8764 17666 8820 18172
rect 8764 17614 8766 17666
rect 8818 17614 8820 17666
rect 8764 17602 8820 17614
rect 9884 18226 9940 18238
rect 9884 18174 9886 18226
rect 9938 18174 9940 18226
rect 9884 17668 9940 18174
rect 9996 18226 10052 18238
rect 10220 18228 10276 18238
rect 9996 18174 9998 18226
rect 10050 18174 10052 18226
rect 9996 17892 10052 18174
rect 10108 18226 10276 18228
rect 10108 18174 10222 18226
rect 10274 18174 10276 18226
rect 10108 18172 10276 18174
rect 10108 18116 10164 18172
rect 10220 18162 10276 18172
rect 10556 18228 10612 18238
rect 10556 18134 10612 18172
rect 10108 18050 10164 18060
rect 10332 18116 10388 18126
rect 10220 17892 10276 17902
rect 9996 17890 10276 17892
rect 9996 17838 10222 17890
rect 10274 17838 10276 17890
rect 9996 17836 10276 17838
rect 10108 17668 10164 17678
rect 9884 17666 10164 17668
rect 9884 17614 10110 17666
rect 10162 17614 10164 17666
rect 9884 17612 10164 17614
rect 1708 17556 1764 17566
rect 1708 17462 1764 17500
rect 2044 17556 2100 17566
rect 2044 17462 2100 17500
rect 8428 17556 8484 17566
rect 8428 17462 8484 17500
rect 2380 17442 2436 17454
rect 2380 17390 2382 17442
rect 2434 17390 2436 17442
rect 1708 16994 1764 17006
rect 1708 16942 1710 16994
rect 1762 16942 1764 16994
rect 1708 16212 1764 16942
rect 2044 16996 2100 17006
rect 2044 16902 2100 16940
rect 2380 16884 2436 17390
rect 2380 16818 2436 16828
rect 2156 16772 2212 16782
rect 1708 16146 1764 16156
rect 2044 16660 2100 16670
rect 2044 16098 2100 16604
rect 2044 16046 2046 16098
rect 2098 16046 2100 16098
rect 2044 16034 2100 16046
rect 1708 15876 1764 15886
rect 1708 15782 1764 15820
rect 1708 15426 1764 15438
rect 1708 15374 1710 15426
rect 1762 15374 1764 15426
rect 1708 14868 1764 15374
rect 2044 15428 2100 15438
rect 2156 15428 2212 16716
rect 10108 16658 10164 17612
rect 10220 16884 10276 17836
rect 10332 16996 10388 18060
rect 10444 17892 10500 17902
rect 10444 17798 10500 17836
rect 10668 17890 10724 18396
rect 10892 18116 10948 18510
rect 11116 18452 11172 18462
rect 10892 18050 10948 18060
rect 11004 18450 11172 18452
rect 11004 18398 11118 18450
rect 11170 18398 11172 18450
rect 11004 18396 11172 18398
rect 10668 17838 10670 17890
rect 10722 17838 10724 17890
rect 10668 17556 10724 17838
rect 10780 17892 10836 17902
rect 11004 17892 11060 18396
rect 11116 18386 11172 18396
rect 10780 17890 11060 17892
rect 10780 17838 10782 17890
rect 10834 17838 11060 17890
rect 10780 17836 11060 17838
rect 10780 17826 10836 17836
rect 11228 17668 11284 18956
rect 11340 17892 11396 19180
rect 11452 19122 11508 19292
rect 12684 19234 12740 19964
rect 12684 19182 12686 19234
rect 12738 19182 12740 19234
rect 12684 19170 12740 19182
rect 11452 19070 11454 19122
rect 11506 19070 11508 19122
rect 11452 19058 11508 19070
rect 11564 18562 11620 18574
rect 11564 18510 11566 18562
rect 11618 18510 11620 18562
rect 11340 17836 11508 17892
rect 10668 17490 10724 17500
rect 10892 17612 11284 17668
rect 11340 17666 11396 17678
rect 11340 17614 11342 17666
rect 11394 17614 11396 17666
rect 10536 17276 10800 17286
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10536 17210 10800 17220
rect 10780 17108 10836 17118
rect 10332 16940 10612 16996
rect 10220 16882 10388 16884
rect 10220 16830 10222 16882
rect 10274 16830 10388 16882
rect 10220 16828 10388 16830
rect 10220 16818 10276 16828
rect 10108 16606 10110 16658
rect 10162 16606 10164 16658
rect 5874 16492 6138 16502
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 5874 16426 6138 16436
rect 8876 16324 8932 16334
rect 8540 16100 8596 16110
rect 8876 16100 8932 16268
rect 9772 16212 9828 16222
rect 8540 16098 8932 16100
rect 8540 16046 8542 16098
rect 8594 16046 8878 16098
rect 8930 16046 8932 16098
rect 8540 16044 8932 16046
rect 2044 15426 2212 15428
rect 2044 15374 2046 15426
rect 2098 15374 2212 15426
rect 2044 15372 2212 15374
rect 2268 15876 2324 15886
rect 2044 15362 2100 15372
rect 1708 14802 1764 14812
rect 2044 14418 2100 14430
rect 2044 14366 2046 14418
rect 2098 14366 2100 14418
rect 1708 14308 1764 14318
rect 1708 14214 1764 14252
rect 2044 14084 2100 14366
rect 2044 14018 2100 14028
rect 1708 13858 1764 13870
rect 1708 13806 1710 13858
rect 1762 13806 1764 13858
rect 1708 13524 1764 13806
rect 2044 13860 2100 13870
rect 2044 13766 2100 13804
rect 1708 13458 1764 13468
rect 2044 12964 2100 12974
rect 2044 12870 2100 12908
rect 1708 12852 1764 12862
rect 1708 12758 1764 12796
rect 1708 12290 1764 12302
rect 1708 12238 1710 12290
rect 1762 12238 1764 12290
rect 1708 11508 1764 12238
rect 2044 12292 2100 12302
rect 2268 12292 2324 15820
rect 8204 15540 8260 15550
rect 6300 15316 6356 15326
rect 5874 14924 6138 14934
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 5874 14858 6138 14868
rect 5874 13356 6138 13366
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 5874 13290 6138 13300
rect 2716 13188 2772 13198
rect 2716 12962 2772 13132
rect 2716 12910 2718 12962
rect 2770 12910 2772 12962
rect 2716 12898 2772 12910
rect 2044 12290 2324 12292
rect 2044 12238 2046 12290
rect 2098 12238 2324 12290
rect 2044 12236 2324 12238
rect 2380 12738 2436 12750
rect 2380 12686 2382 12738
rect 2434 12686 2436 12738
rect 2044 12226 2100 12236
rect 2380 12180 2436 12686
rect 2380 12114 2436 12124
rect 5874 11788 6138 11798
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 5874 11722 6138 11732
rect 1708 11442 1764 11452
rect 2044 11508 2100 11518
rect 2044 11394 2100 11452
rect 2044 11342 2046 11394
rect 2098 11342 2100 11394
rect 2044 11330 2100 11342
rect 1708 11172 1764 11182
rect 1708 11078 1764 11116
rect 1708 10722 1764 10734
rect 1708 10670 1710 10722
rect 1762 10670 1764 10722
rect 1708 10164 1764 10670
rect 2044 10724 2100 10734
rect 2044 10630 2100 10668
rect 5874 10220 6138 10230
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 5874 10154 6138 10164
rect 1708 10098 1764 10108
rect 2044 9828 2100 9838
rect 2044 9734 2100 9772
rect 1708 9604 1764 9614
rect 1708 9510 1764 9548
rect 1708 9154 1764 9166
rect 1708 9102 1710 9154
rect 1762 9102 1764 9154
rect 1708 8820 1764 9102
rect 2044 9156 2100 9166
rect 2044 9062 2100 9100
rect 1708 8754 1764 8764
rect 5874 8652 6138 8662
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 5874 8586 6138 8596
rect 2604 8372 2660 8382
rect 2604 8258 2660 8316
rect 3164 8372 3220 8382
rect 3164 8278 3220 8316
rect 2604 8206 2606 8258
rect 2658 8206 2660 8258
rect 2604 8194 2660 8206
rect 1708 8148 1764 8158
rect 1708 8054 1764 8092
rect 2044 8146 2100 8158
rect 2044 8094 2046 8146
rect 2098 8094 2100 8146
rect 2044 7364 2100 8094
rect 2380 8034 2436 8046
rect 2380 7982 2382 8034
rect 2434 7982 2436 8034
rect 2380 7700 2436 7982
rect 2380 7634 2436 7644
rect 2380 7364 2436 7374
rect 2044 7308 2380 7364
rect 2380 7270 2436 7308
rect 5874 7084 6138 7094
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 5874 7018 6138 7028
rect 5874 5516 6138 5526
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 5874 5450 6138 5460
rect 6300 5348 6356 15260
rect 7644 14756 7700 14766
rect 5964 5292 6356 5348
rect 6412 14644 6468 14654
rect 5964 4562 6020 5292
rect 6412 4564 6468 14588
rect 5964 4510 5966 4562
rect 6018 4510 6020 4562
rect 5964 4498 6020 4510
rect 6300 4562 6468 4564
rect 6300 4510 6414 4562
rect 6466 4510 6468 4562
rect 6300 4508 6468 4510
rect 5628 4338 5684 4350
rect 5628 4286 5630 4338
rect 5682 4286 5684 4338
rect 5404 4228 5460 4238
rect 5628 4228 5684 4286
rect 5404 4226 5684 4228
rect 5404 4174 5406 4226
rect 5458 4174 5684 4226
rect 5404 4172 5684 4174
rect 5404 800 5460 4172
rect 5874 3948 6138 3958
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 5874 3882 6138 3892
rect 6300 3780 6356 4508
rect 6412 4498 6468 4508
rect 6748 13748 6804 13758
rect 5852 3724 6356 3780
rect 5852 3554 5908 3724
rect 5852 3502 5854 3554
rect 5906 3502 5908 3554
rect 5852 3490 5908 3502
rect 6412 3442 6468 3454
rect 6412 3390 6414 3442
rect 6466 3390 6468 3442
rect 6412 3388 6468 3390
rect 6748 3442 6804 13692
rect 7644 4564 7700 14700
rect 7196 4562 7700 4564
rect 7196 4510 7646 4562
rect 7698 4510 7700 4562
rect 7196 4508 7700 4510
rect 6748 3390 6750 3442
rect 6802 3390 6804 3442
rect 6076 3330 6132 3342
rect 6412 3332 6692 3388
rect 6748 3378 6804 3390
rect 6972 4226 7028 4238
rect 6972 4174 6974 4226
rect 7026 4174 7028 4226
rect 6076 3278 6078 3330
rect 6130 3278 6132 3330
rect 6076 800 6132 3278
rect 6636 3220 6692 3332
rect 6972 3220 7028 4174
rect 7196 3554 7252 4508
rect 7644 4498 7700 4508
rect 8092 4228 8148 4238
rect 7196 3502 7198 3554
rect 7250 3502 7252 3554
rect 7196 3490 7252 3502
rect 7868 4226 8148 4228
rect 7868 4174 8094 4226
rect 8146 4174 8148 4226
rect 7868 4172 8148 4174
rect 7868 3554 7924 4172
rect 8092 4162 8148 4172
rect 7868 3502 7870 3554
rect 7922 3502 7924 3554
rect 6636 3164 7028 3220
rect 7420 3330 7476 3342
rect 7420 3278 7422 3330
rect 7474 3278 7476 3330
rect 6748 800 6804 3164
rect 7420 800 7476 3278
rect 7868 2548 7924 3502
rect 8092 3444 8148 3454
rect 8204 3444 8260 15484
rect 8540 14644 8596 16044
rect 8876 16034 8932 16044
rect 9548 16098 9604 16110
rect 9548 16046 9550 16098
rect 9602 16046 9604 16098
rect 9100 15988 9156 15998
rect 9100 15894 9156 15932
rect 9548 15428 9604 16046
rect 9772 15986 9828 16156
rect 9772 15934 9774 15986
rect 9826 15934 9828 15986
rect 9772 15922 9828 15934
rect 10108 16098 10164 16606
rect 10332 16322 10388 16828
rect 10444 16772 10500 16782
rect 10444 16678 10500 16716
rect 10556 16436 10612 16940
rect 10780 16994 10836 17052
rect 10780 16942 10782 16994
rect 10834 16942 10836 16994
rect 10780 16930 10836 16942
rect 10332 16270 10334 16322
rect 10386 16270 10388 16322
rect 10332 16212 10388 16270
rect 10332 16146 10388 16156
rect 10444 16380 10612 16436
rect 10668 16658 10724 16670
rect 10668 16606 10670 16658
rect 10722 16606 10724 16658
rect 10668 16436 10724 16606
rect 10108 16046 10110 16098
rect 10162 16046 10164 16098
rect 10108 15988 10164 16046
rect 10108 15922 10164 15932
rect 10444 15876 10500 16380
rect 10668 16370 10724 16380
rect 10780 16324 10836 16334
rect 10892 16324 10948 17612
rect 11116 17442 11172 17454
rect 11116 17390 11118 17442
rect 11170 17390 11172 17442
rect 11116 16660 11172 17390
rect 11228 17108 11284 17118
rect 11340 17108 11396 17614
rect 11284 17052 11396 17108
rect 11228 17042 11284 17052
rect 11116 16594 11172 16604
rect 10780 16322 11172 16324
rect 10780 16270 10782 16322
rect 10834 16270 11172 16322
rect 10780 16268 11172 16270
rect 10780 16258 10836 16268
rect 10556 16212 10612 16222
rect 10556 16118 10612 16156
rect 10444 15810 10500 15820
rect 10892 15986 10948 15998
rect 10892 15934 10894 15986
rect 10946 15934 10948 15986
rect 10536 15708 10800 15718
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10536 15642 10800 15652
rect 9548 15362 9604 15372
rect 9996 15428 10052 15438
rect 10332 15428 10388 15438
rect 9996 15334 10052 15372
rect 10108 15426 10388 15428
rect 10108 15374 10334 15426
rect 10386 15374 10388 15426
rect 10108 15372 10388 15374
rect 8540 14642 8932 14644
rect 8540 14590 8542 14642
rect 8594 14590 8932 14642
rect 8540 14588 8932 14590
rect 8540 14578 8596 14588
rect 8876 14530 8932 14588
rect 8876 14478 8878 14530
rect 8930 14478 8932 14530
rect 8876 14466 8932 14478
rect 9212 14532 9268 14542
rect 9212 14418 9268 14476
rect 9212 14366 9214 14418
rect 9266 14366 9268 14418
rect 9212 14354 9268 14366
rect 9884 14420 9940 14430
rect 9884 14326 9940 14364
rect 9548 14306 9604 14318
rect 9548 14254 9550 14306
rect 9602 14254 9604 14306
rect 9548 12964 9604 14254
rect 9548 12898 9604 12908
rect 9996 13636 10052 13646
rect 9884 12404 9940 12414
rect 8764 11172 8820 11182
rect 8652 4228 8708 4238
rect 8092 3442 8260 3444
rect 8092 3390 8094 3442
rect 8146 3390 8260 3442
rect 8092 3388 8260 3390
rect 8540 4226 8708 4228
rect 8540 4174 8654 4226
rect 8706 4174 8708 4226
rect 8540 4172 8708 4174
rect 8540 3554 8596 4172
rect 8652 4162 8708 4172
rect 8540 3502 8542 3554
rect 8594 3502 8596 3554
rect 8092 3378 8148 3388
rect 8540 2548 8596 3502
rect 8764 3442 8820 11116
rect 9100 4340 9156 4350
rect 9660 4340 9716 4350
rect 9100 4338 9716 4340
rect 9100 4286 9102 4338
rect 9154 4286 9662 4338
rect 9714 4286 9716 4338
rect 9100 4284 9716 4286
rect 9100 4274 9156 4284
rect 8764 3390 8766 3442
rect 8818 3390 8820 3442
rect 8764 3378 8820 3390
rect 7868 2492 8148 2548
rect 8540 2492 8820 2548
rect 8092 800 8148 2492
rect 8764 800 8820 2492
rect 9436 800 9492 4284
rect 9660 4274 9716 4284
rect 9548 3444 9604 3482
rect 9548 3378 9604 3388
rect 9884 3442 9940 12348
rect 9996 4562 10052 13580
rect 10108 9828 10164 15372
rect 10332 15362 10388 15372
rect 10668 15428 10724 15438
rect 10892 15428 10948 15934
rect 10668 15426 10948 15428
rect 10668 15374 10670 15426
rect 10722 15374 10948 15426
rect 10668 15372 10948 15374
rect 11004 15426 11060 15438
rect 11004 15374 11006 15426
rect 11058 15374 11060 15426
rect 10668 15362 10724 15372
rect 11004 14980 11060 15374
rect 10444 14924 11060 14980
rect 10444 14868 10500 14924
rect 10444 14754 10500 14812
rect 10444 14702 10446 14754
rect 10498 14702 10500 14754
rect 10444 14690 10500 14702
rect 10892 14756 10948 14766
rect 11116 14756 11172 16268
rect 11452 16212 11508 17836
rect 10892 14754 11172 14756
rect 10892 14702 10894 14754
rect 10946 14702 11172 14754
rect 10892 14700 11172 14702
rect 11228 16156 11508 16212
rect 10220 14532 10276 14542
rect 10220 13748 10276 14476
rect 10668 14532 10724 14542
rect 10668 14438 10724 14476
rect 10332 14420 10388 14430
rect 10332 14306 10388 14364
rect 10332 14254 10334 14306
rect 10386 14254 10388 14306
rect 10332 14242 10388 14254
rect 10536 14140 10800 14150
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10536 14074 10800 14084
rect 10556 13972 10612 13982
rect 10332 13748 10388 13758
rect 10556 13748 10612 13916
rect 10220 13746 10388 13748
rect 10220 13694 10334 13746
rect 10386 13694 10388 13746
rect 10220 13692 10388 13694
rect 10220 13186 10276 13692
rect 10332 13682 10388 13692
rect 10444 13746 10612 13748
rect 10444 13694 10558 13746
rect 10610 13694 10612 13746
rect 10444 13692 10612 13694
rect 10220 13134 10222 13186
rect 10274 13134 10276 13186
rect 10220 12178 10276 13134
rect 10220 12126 10222 12178
rect 10274 12126 10276 12178
rect 10220 12114 10276 12126
rect 10332 13188 10388 13198
rect 10444 13188 10500 13692
rect 10556 13682 10612 13692
rect 10780 13522 10836 13534
rect 10780 13470 10782 13522
rect 10834 13470 10836 13522
rect 10780 13412 10836 13470
rect 10780 13346 10836 13356
rect 10332 13186 10500 13188
rect 10332 13134 10334 13186
rect 10386 13134 10500 13186
rect 10332 13132 10500 13134
rect 10780 13188 10836 13198
rect 10892 13188 10948 14700
rect 11228 13860 11284 16156
rect 11452 15988 11508 15998
rect 11452 15894 11508 15932
rect 11340 15764 11396 15774
rect 11340 15428 11396 15708
rect 11340 15334 11396 15372
rect 11004 13804 11284 13860
rect 11452 13860 11508 13870
rect 11004 13746 11060 13804
rect 11452 13766 11508 13804
rect 11004 13694 11006 13746
rect 11058 13694 11060 13746
rect 11004 13300 11060 13694
rect 11116 13524 11172 13534
rect 11116 13430 11172 13468
rect 11004 13244 11172 13300
rect 10780 13186 11060 13188
rect 10780 13134 10782 13186
rect 10834 13134 11060 13186
rect 10780 13132 11060 13134
rect 10332 12178 10388 13132
rect 10780 13122 10836 13132
rect 10556 12964 10612 12974
rect 10556 12870 10612 12908
rect 10892 12850 10948 12862
rect 10892 12798 10894 12850
rect 10946 12798 10948 12850
rect 10536 12572 10800 12582
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10536 12506 10800 12516
rect 10668 12402 10724 12414
rect 10668 12350 10670 12402
rect 10722 12350 10724 12402
rect 10556 12292 10612 12302
rect 10668 12292 10724 12350
rect 10612 12236 10724 12292
rect 10556 12226 10612 12236
rect 10892 12180 10948 12798
rect 10332 12126 10334 12178
rect 10386 12126 10388 12178
rect 10332 12114 10388 12126
rect 10668 12124 10948 12180
rect 10556 12068 10612 12078
rect 10556 11974 10612 12012
rect 10332 11508 10388 11518
rect 10108 9762 10164 9772
rect 10220 11452 10332 11508
rect 9996 4510 9998 4562
rect 10050 4510 10052 4562
rect 9996 4498 10052 4510
rect 10220 3554 10276 11452
rect 10332 11442 10388 11452
rect 10668 11394 10724 12124
rect 11004 12068 11060 13132
rect 11116 13186 11172 13244
rect 11116 13134 11118 13186
rect 11170 13134 11172 13186
rect 11116 13122 11172 13134
rect 11452 13186 11508 13198
rect 11452 13134 11454 13186
rect 11506 13134 11508 13186
rect 11452 13074 11508 13134
rect 11452 13022 11454 13074
rect 11506 13022 11508 13074
rect 11452 13010 11508 13022
rect 11564 12852 11620 18510
rect 11900 18450 11956 18462
rect 11900 18398 11902 18450
rect 11954 18398 11956 18450
rect 11900 18004 11956 18398
rect 12236 18450 12292 18462
rect 12236 18398 12238 18450
rect 12290 18398 12292 18450
rect 12124 18004 12180 18014
rect 11900 17948 12124 18004
rect 12124 17938 12180 17948
rect 12236 17890 12292 18398
rect 12796 18452 12852 20300
rect 12908 20690 12964 20702
rect 12908 20638 12910 20690
rect 12962 20638 12964 20690
rect 12908 20130 12964 20638
rect 13244 20468 13300 21308
rect 13244 20402 13300 20412
rect 13468 20802 13524 21308
rect 13468 20750 13470 20802
rect 13522 20750 13524 20802
rect 12908 20078 12910 20130
rect 12962 20078 12964 20130
rect 12908 20066 12964 20078
rect 13244 20020 13300 20030
rect 13244 19926 13300 19964
rect 12908 19010 12964 19022
rect 12908 18958 12910 19010
rect 12962 18958 12964 19010
rect 12908 18676 12964 18958
rect 13468 18788 13524 20750
rect 13580 20132 13636 22876
rect 13692 21588 13748 21598
rect 13692 20356 13748 21532
rect 13804 20692 13860 20702
rect 13804 20598 13860 20636
rect 13692 20290 13748 20300
rect 13916 20188 13972 22876
rect 14028 22596 14084 23326
rect 14140 23154 14196 24220
rect 14476 24162 14532 25564
rect 14476 24110 14478 24162
rect 14530 24110 14532 24162
rect 14476 24098 14532 24110
rect 14588 23940 14644 29148
rect 14700 28420 14756 28430
rect 14700 27970 14756 28364
rect 14700 27918 14702 27970
rect 14754 27918 14756 27970
rect 14700 27906 14756 27918
rect 14812 28084 14868 28094
rect 14812 27858 14868 28028
rect 14812 27806 14814 27858
rect 14866 27806 14868 27858
rect 14812 27794 14868 27806
rect 14924 27636 14980 30044
rect 15372 29316 15428 29326
rect 15372 29222 15428 29260
rect 14812 27580 14980 27636
rect 15036 29204 15092 29214
rect 15036 27634 15092 29148
rect 15198 29036 15462 29046
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15198 28970 15462 28980
rect 15484 28868 15540 28878
rect 15596 28868 15652 30156
rect 15708 29092 15764 36206
rect 15932 35922 15988 36428
rect 16044 36372 16100 36382
rect 16156 36372 16212 39200
rect 16828 36932 16884 39200
rect 16380 36876 16884 36932
rect 16156 36316 16324 36372
rect 16044 36278 16100 36316
rect 15932 35870 15934 35922
rect 15986 35870 15988 35922
rect 15932 35858 15988 35870
rect 16268 35924 16324 36316
rect 16380 36370 16436 36876
rect 16380 36318 16382 36370
rect 16434 36318 16436 36370
rect 16380 36306 16436 36318
rect 17276 36482 17332 36494
rect 17276 36430 17278 36482
rect 17330 36430 17332 36482
rect 16380 35924 16436 35934
rect 16268 35922 16436 35924
rect 16268 35870 16382 35922
rect 16434 35870 16436 35922
rect 16268 35868 16436 35870
rect 16380 35858 16436 35868
rect 16604 35700 16660 35710
rect 16380 35698 16660 35700
rect 16380 35646 16606 35698
rect 16658 35646 16660 35698
rect 16380 35644 16660 35646
rect 15820 29428 15876 29438
rect 15820 29334 15876 29372
rect 16268 29316 16324 29326
rect 16268 29222 16324 29260
rect 16156 29204 16212 29214
rect 16156 29110 16212 29148
rect 15708 29036 16100 29092
rect 16044 28980 16100 29036
rect 16044 28924 16324 28980
rect 15484 28866 15652 28868
rect 15484 28814 15486 28866
rect 15538 28814 15652 28866
rect 15484 28812 15652 28814
rect 15820 28868 15876 28878
rect 15484 28802 15540 28812
rect 15820 28774 15876 28812
rect 15596 28644 15652 28654
rect 15596 28642 15764 28644
rect 15596 28590 15598 28642
rect 15650 28590 15764 28642
rect 15596 28588 15764 28590
rect 15596 28578 15652 28588
rect 15708 28084 15764 28588
rect 15596 27972 15652 27982
rect 15596 27878 15652 27916
rect 15036 27582 15038 27634
rect 15090 27582 15092 27634
rect 14700 26292 14756 26302
rect 14700 26198 14756 26236
rect 14700 25844 14756 25854
rect 14700 24724 14756 25788
rect 14812 24946 14868 27580
rect 15036 27300 15092 27582
rect 15260 27858 15316 27870
rect 15260 27806 15262 27858
rect 15314 27806 15316 27858
rect 15260 27636 15316 27806
rect 15708 27858 15764 28028
rect 15708 27806 15710 27858
rect 15762 27806 15764 27858
rect 15708 27794 15764 27806
rect 16044 28642 16100 28654
rect 16044 28590 16046 28642
rect 16098 28590 16100 28642
rect 16044 27858 16100 28590
rect 16044 27806 16046 27858
rect 16098 27806 16100 27858
rect 15932 27636 15988 27646
rect 15260 27580 15652 27636
rect 15198 27468 15462 27478
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15198 27402 15462 27412
rect 15596 27412 15652 27580
rect 15932 27542 15988 27580
rect 16044 27412 16100 27806
rect 15596 27356 16100 27412
rect 16156 28084 16212 28094
rect 15596 27300 15652 27356
rect 15036 27234 15092 27244
rect 15148 27244 15652 27300
rect 14924 27074 14980 27086
rect 14924 27022 14926 27074
rect 14978 27022 14980 27074
rect 14924 26908 14980 27022
rect 15148 26962 15204 27244
rect 15932 27186 15988 27356
rect 15932 27134 15934 27186
rect 15986 27134 15988 27186
rect 15932 27122 15988 27134
rect 15372 27076 15428 27086
rect 15372 26982 15428 27020
rect 15708 27074 15764 27086
rect 16156 27076 16212 28028
rect 15708 27022 15710 27074
rect 15762 27022 15764 27074
rect 15148 26910 15150 26962
rect 15202 26910 15204 26962
rect 14924 26852 15092 26908
rect 15148 26898 15204 26910
rect 15036 25844 15092 26852
rect 15708 26516 15764 27022
rect 16044 27074 16212 27076
rect 16044 27022 16158 27074
rect 16210 27022 16212 27074
rect 16044 27020 16212 27022
rect 15596 26404 15652 26414
rect 15596 26310 15652 26348
rect 15708 26180 15764 26460
rect 15932 26516 15988 26526
rect 16044 26516 16100 27020
rect 16156 27010 16212 27020
rect 15932 26514 16100 26516
rect 15932 26462 15934 26514
rect 15986 26462 16100 26514
rect 15932 26460 16100 26462
rect 16156 26852 16212 26862
rect 15932 26450 15988 26460
rect 15708 26114 15764 26124
rect 15820 26068 15876 26078
rect 15198 25900 15462 25910
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15198 25834 15462 25844
rect 15036 25732 15092 25788
rect 15260 25732 15316 25742
rect 15036 25730 15316 25732
rect 15036 25678 15262 25730
rect 15314 25678 15316 25730
rect 15036 25676 15316 25678
rect 15260 25666 15316 25676
rect 14812 24894 14814 24946
rect 14866 24894 14868 24946
rect 14812 24882 14868 24894
rect 14924 25620 14980 25630
rect 14700 24668 14868 24724
rect 14700 24500 14756 24510
rect 14700 24162 14756 24444
rect 14700 24110 14702 24162
rect 14754 24110 14756 24162
rect 14700 24098 14756 24110
rect 14812 24162 14868 24668
rect 14812 24110 14814 24162
rect 14866 24110 14868 24162
rect 14812 23940 14868 24110
rect 14588 23874 14644 23884
rect 14700 23884 14868 23940
rect 14364 23828 14420 23838
rect 14364 23734 14420 23772
rect 14140 23102 14142 23154
rect 14194 23102 14196 23154
rect 14140 23090 14196 23102
rect 14700 23042 14756 23884
rect 14812 23156 14868 23166
rect 14812 23062 14868 23100
rect 14924 23156 14980 25564
rect 15148 25508 15204 25546
rect 15148 25442 15204 25452
rect 15148 25284 15204 25294
rect 15260 25284 15316 25294
rect 15204 25282 15316 25284
rect 15204 25230 15262 25282
rect 15314 25230 15316 25282
rect 15204 25228 15316 25230
rect 15148 25218 15204 25228
rect 15260 25218 15316 25228
rect 15820 25284 15876 26012
rect 16156 25618 16212 26796
rect 16268 26628 16324 28924
rect 16268 26562 16324 26572
rect 16268 26290 16324 26302
rect 16268 26238 16270 26290
rect 16322 26238 16324 26290
rect 16268 26068 16324 26238
rect 16268 26002 16324 26012
rect 16380 25620 16436 35644
rect 16604 35634 16660 35644
rect 16940 29540 16996 29550
rect 16716 29428 16772 29438
rect 16716 29334 16772 29372
rect 16492 29204 16548 29214
rect 16492 28754 16548 29148
rect 16604 29202 16660 29214
rect 16604 29150 16606 29202
rect 16658 29150 16660 29202
rect 16604 28868 16660 29150
rect 16604 28802 16660 28812
rect 16940 28756 16996 29484
rect 16492 28702 16494 28754
rect 16546 28702 16548 28754
rect 16492 28690 16548 28702
rect 16828 28754 16996 28756
rect 16828 28702 16942 28754
rect 16994 28702 16996 28754
rect 16828 28700 16996 28702
rect 16828 27748 16884 28700
rect 16940 28690 16996 28700
rect 17276 28644 17332 36430
rect 17500 36370 17556 39200
rect 17500 36318 17502 36370
rect 17554 36318 17556 36370
rect 17500 36306 17556 36318
rect 17948 36482 18004 36494
rect 17948 36430 17950 36482
rect 18002 36430 18004 36482
rect 17388 35812 17444 35822
rect 17444 35756 17556 35812
rect 17388 35746 17444 35756
rect 17388 29986 17444 29998
rect 17388 29934 17390 29986
rect 17442 29934 17444 29986
rect 17388 29428 17444 29934
rect 17388 29362 17444 29372
rect 17388 28756 17444 28766
rect 17500 28756 17556 35756
rect 17388 28754 17556 28756
rect 17388 28702 17390 28754
rect 17442 28702 17556 28754
rect 17388 28700 17556 28702
rect 17388 28690 17444 28700
rect 17276 28578 17332 28588
rect 17500 27972 17556 28700
rect 17500 27906 17556 27916
rect 17724 35588 17780 35598
rect 16828 27682 16884 27692
rect 16940 27746 16996 27758
rect 16940 27694 16942 27746
rect 16994 27694 16996 27746
rect 16940 27076 16996 27694
rect 17500 27748 17556 27758
rect 17500 27654 17556 27692
rect 17388 27636 17444 27646
rect 17724 27636 17780 35532
rect 17948 31892 18004 36430
rect 18172 36370 18228 39200
rect 18172 36318 18174 36370
rect 18226 36318 18228 36370
rect 18172 36306 18228 36318
rect 18508 36370 18564 36382
rect 18508 36318 18510 36370
rect 18562 36318 18564 36370
rect 17948 31826 18004 31836
rect 18396 29988 18452 29998
rect 17836 29426 17892 29438
rect 17836 29374 17838 29426
rect 17890 29374 17892 29426
rect 17836 28642 17892 29374
rect 17948 29428 18004 29438
rect 17948 29334 18004 29372
rect 18060 29426 18116 29438
rect 18060 29374 18062 29426
rect 18114 29374 18116 29426
rect 17836 28590 17838 28642
rect 17890 28590 17892 28642
rect 17836 27748 17892 28590
rect 17948 29204 18004 29214
rect 17948 28642 18004 29148
rect 17948 28590 17950 28642
rect 18002 28590 18004 28642
rect 17948 28578 18004 28590
rect 18060 28644 18116 29374
rect 18284 29426 18340 29438
rect 18284 29374 18286 29426
rect 18338 29374 18340 29426
rect 18284 28644 18340 29374
rect 18396 29204 18452 29932
rect 18508 29428 18564 36318
rect 18508 29362 18564 29372
rect 18620 36372 18676 36382
rect 18620 29204 18676 36316
rect 18844 36370 18900 39200
rect 19292 36484 19348 36494
rect 19292 36482 19460 36484
rect 19292 36430 19294 36482
rect 19346 36430 19460 36482
rect 19292 36428 19460 36430
rect 19292 36418 19348 36428
rect 18844 36318 18846 36370
rect 18898 36318 18900 36370
rect 18844 36306 18900 36318
rect 18732 31892 18788 31902
rect 18732 30098 18788 31836
rect 18956 30212 19012 30222
rect 18732 30046 18734 30098
rect 18786 30046 18788 30098
rect 18732 30034 18788 30046
rect 18844 30210 19012 30212
rect 18844 30158 18958 30210
rect 19010 30158 19012 30210
rect 18844 30156 19012 30158
rect 18732 29652 18788 29662
rect 18844 29652 18900 30156
rect 18956 30146 19012 30156
rect 18732 29650 18900 29652
rect 18732 29598 18734 29650
rect 18786 29598 18900 29650
rect 18732 29596 18900 29598
rect 19292 29988 19348 29998
rect 18732 29586 18788 29596
rect 19292 29538 19348 29932
rect 19292 29486 19294 29538
rect 19346 29486 19348 29538
rect 19292 29474 19348 29486
rect 19404 29316 19460 36428
rect 19516 36370 19572 39200
rect 19852 36372 19908 36382
rect 19516 36318 19518 36370
rect 19570 36318 19572 36370
rect 19516 36306 19572 36318
rect 19740 36370 19908 36372
rect 19740 36318 19854 36370
rect 19906 36318 19908 36370
rect 19740 36316 19908 36318
rect 19628 29988 19684 29998
rect 19516 29986 19684 29988
rect 19516 29934 19630 29986
rect 19682 29934 19684 29986
rect 19516 29932 19684 29934
rect 19516 29540 19572 29932
rect 19628 29922 19684 29932
rect 19628 29652 19684 29662
rect 19628 29558 19684 29596
rect 19516 29474 19572 29484
rect 19404 29260 19684 29316
rect 18396 29138 18452 29148
rect 18508 29148 18676 29204
rect 18396 28644 18452 28654
rect 18060 28642 18228 28644
rect 18060 28590 18062 28642
rect 18114 28590 18228 28642
rect 18060 28588 18228 28590
rect 18284 28642 18452 28644
rect 18284 28590 18398 28642
rect 18450 28590 18452 28642
rect 18284 28588 18452 28590
rect 18060 28578 18116 28588
rect 18172 28084 18228 28588
rect 18396 28196 18452 28588
rect 18508 28308 18564 29148
rect 18732 28868 18788 28878
rect 18732 28866 19236 28868
rect 18732 28814 18734 28866
rect 18786 28814 19236 28866
rect 18732 28812 19236 28814
rect 18732 28802 18788 28812
rect 19180 28642 19236 28812
rect 19180 28590 19182 28642
rect 19234 28590 19236 28642
rect 19180 28578 19236 28590
rect 18956 28420 19012 28430
rect 18956 28326 19012 28364
rect 18508 28252 18788 28308
rect 18396 28140 18676 28196
rect 18172 28028 18452 28084
rect 17948 27972 18004 27982
rect 18004 27916 18340 27972
rect 17948 27906 18004 27916
rect 18284 27858 18340 27916
rect 18284 27806 18286 27858
rect 18338 27806 18340 27858
rect 18060 27748 18116 27758
rect 17836 27746 18116 27748
rect 17836 27694 18062 27746
rect 18114 27694 18116 27746
rect 17836 27692 18116 27694
rect 17724 27580 18004 27636
rect 17388 27542 17444 27580
rect 17948 27300 18004 27580
rect 18060 27524 18116 27692
rect 18060 27458 18116 27468
rect 18172 27748 18228 27758
rect 17948 27244 18116 27300
rect 17388 27076 17444 27086
rect 16940 27074 17444 27076
rect 16940 27022 17390 27074
rect 17442 27022 17444 27074
rect 16940 27020 17444 27022
rect 17388 26964 17444 27020
rect 17836 27076 17892 27086
rect 17388 26898 17444 26908
rect 17612 26964 17668 27002
rect 17612 26898 17668 26908
rect 16604 26516 16660 26526
rect 16604 26422 16660 26460
rect 17836 26514 17892 27020
rect 17948 27074 18004 27086
rect 17948 27022 17950 27074
rect 18002 27022 18004 27074
rect 17948 26852 18004 27022
rect 17948 26786 18004 26796
rect 17836 26462 17838 26514
rect 17890 26462 17892 26514
rect 17836 26450 17892 26462
rect 17948 26628 18004 26638
rect 17164 26404 17220 26414
rect 17052 26348 17164 26404
rect 16716 26178 16772 26190
rect 16716 26126 16718 26178
rect 16770 26126 16772 26178
rect 16156 25566 16158 25618
rect 16210 25566 16212 25618
rect 16156 25554 16212 25566
rect 16268 25564 16436 25620
rect 16604 25732 16660 25742
rect 15820 25190 15876 25228
rect 15932 25060 15988 25070
rect 15148 24724 15204 24734
rect 15484 24724 15540 24734
rect 15148 24722 15540 24724
rect 15148 24670 15150 24722
rect 15202 24670 15486 24722
rect 15538 24670 15540 24722
rect 15148 24668 15540 24670
rect 15148 24658 15204 24668
rect 15484 24658 15540 24668
rect 15596 24498 15652 24510
rect 15596 24446 15598 24498
rect 15650 24446 15652 24498
rect 15198 24332 15462 24342
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15198 24266 15462 24276
rect 15372 23828 15428 23838
rect 15596 23828 15652 24446
rect 15820 24500 15876 24510
rect 15932 24500 15988 25004
rect 16268 24948 16324 25564
rect 16604 25508 16660 25676
rect 16380 25394 16436 25406
rect 16380 25342 16382 25394
rect 16434 25342 16436 25394
rect 16380 25284 16436 25342
rect 16380 25218 16436 25228
rect 16492 25394 16548 25406
rect 16492 25342 16494 25394
rect 16546 25342 16548 25394
rect 16492 25060 16548 25342
rect 16492 24994 16548 25004
rect 16268 24882 16324 24892
rect 15820 24498 15988 24500
rect 15820 24446 15822 24498
rect 15874 24446 15988 24498
rect 15820 24444 15988 24446
rect 15820 24434 15876 24444
rect 15372 23826 15652 23828
rect 15372 23774 15374 23826
rect 15426 23774 15652 23826
rect 15372 23772 15652 23774
rect 15372 23762 15428 23772
rect 15596 23268 15652 23772
rect 15596 23202 15652 23212
rect 15036 23156 15092 23166
rect 14924 23154 15092 23156
rect 14924 23102 15038 23154
rect 15090 23102 15092 23154
rect 14924 23100 15092 23102
rect 14700 22990 14702 23042
rect 14754 22990 14756 23042
rect 14588 22930 14644 22942
rect 14588 22878 14590 22930
rect 14642 22878 14644 22930
rect 14588 22596 14644 22878
rect 14028 22540 14420 22596
rect 14140 22372 14196 22382
rect 14140 22258 14196 22316
rect 14364 22370 14420 22540
rect 14588 22530 14644 22540
rect 14364 22318 14366 22370
rect 14418 22318 14420 22370
rect 14364 22306 14420 22318
rect 14476 22484 14532 22494
rect 14140 22206 14142 22258
rect 14194 22206 14196 22258
rect 14140 22194 14196 22206
rect 14476 21364 14532 22428
rect 14700 22260 14756 22990
rect 14700 22194 14756 22204
rect 14812 22260 14868 22270
rect 14924 22260 14980 23100
rect 15036 23090 15092 23100
rect 15198 22764 15462 22774
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15198 22698 15462 22708
rect 14812 22258 14980 22260
rect 14812 22206 14814 22258
rect 14866 22206 14980 22258
rect 14812 22204 14980 22206
rect 15036 22370 15092 22382
rect 15036 22318 15038 22370
rect 15090 22318 15092 22370
rect 14812 22194 14868 22204
rect 15036 21588 15092 22318
rect 15484 22260 15540 22270
rect 15932 22260 15988 24444
rect 16044 24836 16100 24846
rect 16044 24722 16100 24780
rect 16044 24670 16046 24722
rect 16098 24670 16100 24722
rect 16044 24276 16100 24670
rect 16604 24612 16660 25452
rect 16156 24556 16660 24612
rect 16716 25284 16772 26126
rect 16940 26068 16996 26078
rect 16716 24612 16772 25228
rect 16828 25506 16884 25518
rect 16828 25454 16830 25506
rect 16882 25454 16884 25506
rect 16828 24836 16884 25454
rect 16828 24770 16884 24780
rect 16940 25508 16996 26012
rect 16828 24612 16884 24622
rect 16716 24610 16884 24612
rect 16716 24558 16830 24610
rect 16882 24558 16884 24610
rect 16716 24556 16884 24558
rect 16156 24498 16212 24556
rect 16828 24546 16884 24556
rect 16156 24446 16158 24498
rect 16210 24446 16212 24498
rect 16156 24434 16212 24446
rect 16044 24220 16324 24276
rect 16268 23826 16324 24220
rect 16268 23774 16270 23826
rect 16322 23774 16324 23826
rect 16268 23762 16324 23774
rect 16380 23996 16660 24052
rect 16380 23156 16436 23996
rect 16604 23938 16660 23996
rect 16604 23886 16606 23938
rect 16658 23886 16660 23938
rect 16604 23874 16660 23886
rect 16492 23828 16548 23838
rect 16492 23378 16548 23772
rect 16492 23326 16494 23378
rect 16546 23326 16548 23378
rect 16492 23314 16548 23326
rect 16716 23156 16772 23166
rect 16380 23044 16436 23100
rect 16604 23154 16772 23156
rect 16604 23102 16718 23154
rect 16770 23102 16772 23154
rect 16604 23100 16772 23102
rect 16380 22988 16548 23044
rect 16268 22260 16324 22270
rect 15932 22258 16324 22260
rect 15932 22206 16270 22258
rect 16322 22206 16324 22258
rect 15932 22204 16324 22206
rect 15484 22166 15540 22204
rect 16268 22194 16324 22204
rect 15820 22148 15876 22158
rect 15820 22054 15876 22092
rect 14476 21298 14532 21308
rect 14700 21532 15036 21588
rect 14364 20916 14420 20926
rect 14364 20822 14420 20860
rect 14140 20802 14196 20814
rect 14140 20750 14142 20802
rect 14194 20750 14196 20802
rect 14140 20692 14196 20750
rect 14140 20626 14196 20636
rect 14588 20802 14644 20814
rect 14588 20750 14590 20802
rect 14642 20750 14644 20802
rect 14588 20692 14644 20750
rect 14588 20626 14644 20636
rect 14252 20580 14308 20590
rect 14252 20486 14308 20524
rect 14700 20188 14756 21532
rect 15036 21522 15092 21532
rect 15260 22036 15316 22046
rect 15260 21586 15316 21980
rect 15708 21924 15764 21934
rect 15764 21868 15876 21924
rect 15708 21858 15764 21868
rect 15260 21534 15262 21586
rect 15314 21534 15316 21586
rect 15260 21522 15316 21534
rect 15484 21588 15540 21598
rect 15484 21586 15652 21588
rect 15484 21534 15486 21586
rect 15538 21534 15652 21586
rect 15484 21532 15652 21534
rect 15484 21522 15540 21532
rect 14924 21364 14980 21402
rect 14924 21298 14980 21308
rect 15036 21362 15092 21374
rect 15036 21310 15038 21362
rect 15090 21310 15092 21362
rect 14924 21140 14980 21150
rect 14924 20802 14980 21084
rect 14924 20750 14926 20802
rect 14978 20750 14980 20802
rect 14924 20738 14980 20750
rect 15036 20692 15092 21310
rect 15198 21196 15462 21206
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15198 21130 15462 21140
rect 15596 20914 15652 21532
rect 15596 20862 15598 20914
rect 15650 20862 15652 20914
rect 15596 20804 15652 20862
rect 15148 20692 15204 20702
rect 15036 20636 15148 20692
rect 14924 20356 14980 20366
rect 14924 20188 14980 20300
rect 13916 20132 14196 20188
rect 14700 20132 14868 20188
rect 14924 20132 15092 20188
rect 13580 20130 13860 20132
rect 13580 20078 13582 20130
rect 13634 20078 13860 20130
rect 13580 20076 13860 20078
rect 13580 20066 13636 20076
rect 13468 18722 13524 18732
rect 12908 18620 13188 18676
rect 12908 18452 12964 18462
rect 12796 18450 12964 18452
rect 12796 18398 12910 18450
rect 12962 18398 12964 18450
rect 12796 18396 12964 18398
rect 12908 18386 12964 18396
rect 13020 18452 13076 18462
rect 13020 18358 13076 18396
rect 12460 18228 12516 18238
rect 12236 17838 12238 17890
rect 12290 17838 12292 17890
rect 11676 17556 11732 17566
rect 11676 16772 11732 17500
rect 11676 16706 11732 16716
rect 12236 16882 12292 17838
rect 12348 18226 12516 18228
rect 12348 18174 12462 18226
rect 12514 18174 12516 18226
rect 12348 18172 12516 18174
rect 12348 17666 12404 18172
rect 12460 18162 12516 18172
rect 12684 18226 12740 18238
rect 12684 18174 12686 18226
rect 12738 18174 12740 18226
rect 12684 17892 12740 18174
rect 12684 17826 12740 17836
rect 12908 18004 12964 18014
rect 12908 17890 12964 17948
rect 12908 17838 12910 17890
rect 12962 17838 12964 17890
rect 12908 17826 12964 17838
rect 12348 17614 12350 17666
rect 12402 17614 12404 17666
rect 12348 17108 12404 17614
rect 12572 17666 12628 17678
rect 12572 17614 12574 17666
rect 12626 17614 12628 17666
rect 12572 17556 12628 17614
rect 12572 17490 12628 17500
rect 12796 17668 12852 17678
rect 13132 17668 13188 18620
rect 13356 18562 13412 18574
rect 13356 18510 13358 18562
rect 13410 18510 13412 18562
rect 13356 18340 13412 18510
rect 13692 18452 13748 18462
rect 13692 18358 13748 18396
rect 13356 18274 13412 18284
rect 12796 17666 13188 17668
rect 12796 17614 12798 17666
rect 12850 17614 13188 17666
rect 12796 17612 13188 17614
rect 12348 17052 12628 17108
rect 12236 16830 12238 16882
rect 12290 16830 12292 16882
rect 12236 16324 12292 16830
rect 12460 16660 12516 16670
rect 12572 16660 12628 17052
rect 11788 16322 12292 16324
rect 11788 16270 12238 16322
rect 12290 16270 12292 16322
rect 11788 16268 12292 16270
rect 11788 15986 11844 16268
rect 12236 16258 12292 16268
rect 12348 16658 12628 16660
rect 12348 16606 12462 16658
rect 12514 16606 12628 16658
rect 12348 16604 12628 16606
rect 12684 16658 12740 16670
rect 12684 16606 12686 16658
rect 12738 16606 12740 16658
rect 12348 16098 12404 16604
rect 12460 16594 12516 16604
rect 12684 16548 12740 16606
rect 12684 16482 12740 16492
rect 12796 16660 12852 17612
rect 13356 16994 13412 17006
rect 13356 16942 13358 16994
rect 13410 16942 13412 16994
rect 13020 16884 13076 16894
rect 13020 16790 13076 16828
rect 12908 16660 12964 16670
rect 12796 16658 12964 16660
rect 12796 16606 12910 16658
rect 12962 16606 12964 16658
rect 12796 16604 12964 16606
rect 12572 16212 12628 16222
rect 12572 16118 12628 16156
rect 12348 16046 12350 16098
rect 12402 16046 12404 16098
rect 11788 15934 11790 15986
rect 11842 15934 11844 15986
rect 11788 15922 11844 15934
rect 12012 15988 12068 15998
rect 11676 15764 11732 15774
rect 11676 14642 11732 15708
rect 11676 14590 11678 14642
rect 11730 14590 11732 14642
rect 11676 14578 11732 14590
rect 12012 15202 12068 15932
rect 12348 15988 12404 16046
rect 12796 16100 12852 16604
rect 12908 16594 12964 16604
rect 12796 16006 12852 16044
rect 12348 15922 12404 15932
rect 12908 15988 12964 15998
rect 12908 15986 13076 15988
rect 12908 15934 12910 15986
rect 12962 15934 13076 15986
rect 12908 15932 13076 15934
rect 12908 15922 12964 15932
rect 12460 15876 12516 15886
rect 12460 15540 12516 15820
rect 12012 15150 12014 15202
rect 12066 15150 12068 15202
rect 11900 14420 11956 14430
rect 11788 14364 11900 14420
rect 11676 13746 11732 13758
rect 11676 13694 11678 13746
rect 11730 13694 11732 13746
rect 11676 13524 11732 13694
rect 11676 13458 11732 13468
rect 10780 12012 11060 12068
rect 11228 12796 11620 12852
rect 10780 11954 10836 12012
rect 10780 11902 10782 11954
rect 10834 11902 10836 11954
rect 10780 11890 10836 11902
rect 11004 11732 11060 11742
rect 10668 11342 10670 11394
rect 10722 11342 10724 11394
rect 10668 11330 10724 11342
rect 10892 11676 11004 11732
rect 10332 11170 10388 11182
rect 10332 11118 10334 11170
rect 10386 11118 10388 11170
rect 10332 9156 10388 11118
rect 10536 11004 10800 11014
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10536 10938 10800 10948
rect 10536 9436 10800 9446
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10536 9370 10800 9380
rect 10332 9090 10388 9100
rect 10536 7868 10800 7878
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10536 7802 10800 7812
rect 10536 6300 10800 6310
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10536 6234 10800 6244
rect 10536 4732 10800 4742
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10536 4666 10800 4676
rect 10220 3502 10222 3554
rect 10274 3502 10276 3554
rect 10220 3490 10276 3502
rect 10444 4226 10500 4238
rect 10444 4174 10446 4226
rect 10498 4174 10500 4226
rect 9884 3390 9886 3442
rect 9938 3390 9940 3442
rect 9884 3378 9940 3390
rect 10108 3444 10164 3454
rect 10108 3332 10164 3388
rect 10444 3332 10500 4174
rect 10892 3554 10948 11676
rect 11004 11666 11060 11676
rect 11004 11170 11060 11182
rect 11004 11118 11006 11170
rect 11058 11118 11060 11170
rect 11004 10724 11060 11118
rect 11004 10658 11060 10668
rect 11228 8372 11284 12796
rect 11340 12292 11396 12302
rect 11676 12292 11732 12302
rect 11340 11394 11396 12236
rect 11340 11342 11342 11394
rect 11394 11342 11396 11394
rect 11340 11330 11396 11342
rect 11564 12236 11676 12292
rect 11228 8306 11284 8316
rect 10892 3502 10894 3554
rect 10946 3502 10948 3554
rect 10892 3490 10948 3502
rect 11564 3554 11620 12236
rect 11676 12226 11732 12236
rect 11788 12178 11844 14364
rect 11900 14326 11956 14364
rect 12012 14196 12068 15150
rect 12236 15538 12516 15540
rect 12236 15486 12462 15538
rect 12514 15486 12516 15538
rect 12236 15484 12516 15486
rect 12236 14530 12292 15484
rect 12460 15474 12516 15484
rect 12796 15428 12852 15438
rect 12236 14478 12238 14530
rect 12290 14478 12292 14530
rect 12236 14466 12292 14478
rect 12684 15426 12852 15428
rect 12684 15374 12798 15426
rect 12850 15374 12852 15426
rect 12684 15372 12852 15374
rect 12572 14308 12628 14318
rect 12572 14214 12628 14252
rect 12460 14196 12516 14206
rect 12012 14140 12460 14196
rect 12460 13746 12516 14140
rect 12684 14084 12740 15372
rect 12796 15362 12852 15372
rect 13020 15314 13076 15932
rect 13020 15262 13022 15314
rect 13074 15262 13076 15314
rect 13020 15250 13076 15262
rect 12796 14530 12852 14542
rect 12796 14478 12798 14530
rect 12850 14478 12852 14530
rect 12796 14308 12852 14478
rect 12796 14242 12852 14252
rect 12908 14420 12964 14430
rect 12460 13694 12462 13746
rect 12514 13694 12516 13746
rect 12460 13682 12516 13694
rect 12572 14028 12740 14084
rect 12572 12964 12628 14028
rect 12796 13972 12852 13982
rect 12460 12908 12628 12964
rect 12684 13916 12796 13972
rect 12684 13858 12740 13916
rect 12796 13906 12852 13916
rect 12684 13806 12686 13858
rect 12738 13806 12740 13858
rect 11788 12126 11790 12178
rect 11842 12126 11844 12178
rect 11788 12114 11844 12126
rect 12236 12404 12292 12414
rect 12236 12178 12292 12348
rect 12236 12126 12238 12178
rect 12290 12126 12292 12178
rect 12236 12114 12292 12126
rect 12012 12068 12068 12078
rect 12012 11974 12068 12012
rect 11676 11956 11732 11966
rect 11676 11862 11732 11900
rect 12348 11954 12404 11966
rect 12348 11902 12350 11954
rect 12402 11902 12404 11954
rect 12348 11396 12404 11902
rect 12460 11732 12516 12908
rect 12572 12738 12628 12750
rect 12572 12686 12574 12738
rect 12626 12686 12628 12738
rect 12572 11844 12628 12686
rect 12684 12178 12740 13806
rect 12796 12962 12852 12974
rect 12796 12910 12798 12962
rect 12850 12910 12852 12962
rect 12796 12740 12852 12910
rect 12796 12674 12852 12684
rect 12684 12126 12686 12178
rect 12738 12126 12740 12178
rect 12684 11956 12740 12126
rect 12908 12178 12964 14364
rect 13244 14196 13300 14206
rect 13244 13970 13300 14140
rect 13244 13918 13246 13970
rect 13298 13918 13300 13970
rect 13244 13906 13300 13918
rect 12908 12126 12910 12178
rect 12962 12126 12964 12178
rect 12908 12114 12964 12126
rect 13132 13412 13188 13422
rect 13356 13412 13412 16942
rect 13580 16884 13636 16894
rect 13580 16790 13636 16828
rect 13804 16212 13860 20076
rect 14140 20130 14196 20132
rect 14140 20078 14142 20130
rect 14194 20078 14196 20130
rect 14140 20066 14196 20078
rect 14476 20018 14532 20030
rect 14476 19966 14478 20018
rect 14530 19966 14532 20018
rect 14476 19460 14532 19966
rect 14476 19394 14532 19404
rect 14700 19572 14756 19582
rect 14700 19122 14756 19516
rect 14700 19070 14702 19122
rect 14754 19070 14756 19122
rect 14364 19012 14420 19022
rect 14364 18918 14420 18956
rect 14252 18788 14308 18798
rect 14308 18732 14532 18788
rect 14252 18722 14308 18732
rect 14252 18340 14308 18350
rect 14252 18246 14308 18284
rect 13804 16156 13972 16212
rect 13468 15988 13524 15998
rect 13468 15894 13524 15932
rect 13804 15988 13860 15998
rect 13804 15894 13860 15932
rect 13916 15148 13972 16156
rect 14140 16100 14196 16110
rect 14028 15988 14084 15998
rect 14028 15538 14084 15932
rect 14028 15486 14030 15538
rect 14082 15486 14084 15538
rect 14028 15474 14084 15486
rect 13916 15092 14084 15148
rect 13132 12852 13188 13356
rect 13132 12178 13188 12796
rect 13132 12126 13134 12178
rect 13186 12126 13188 12178
rect 13132 12114 13188 12126
rect 13244 13356 13412 13412
rect 13468 14530 13524 14542
rect 13468 14478 13470 14530
rect 13522 14478 13524 14530
rect 13468 13972 13524 14478
rect 13692 14530 13748 14542
rect 13692 14478 13694 14530
rect 13746 14478 13748 14530
rect 13692 14420 13748 14478
rect 13916 14532 13972 14542
rect 13916 14438 13972 14476
rect 13580 14308 13636 14318
rect 13580 14214 13636 14252
rect 12684 11890 12740 11900
rect 12572 11778 12628 11788
rect 12460 11666 12516 11676
rect 12348 11330 12404 11340
rect 11564 3502 11566 3554
rect 11618 3502 11620 3554
rect 11564 3490 11620 3502
rect 12348 8484 12404 8494
rect 12348 3554 12404 8428
rect 13244 7364 13300 13356
rect 13356 13188 13412 13198
rect 13356 12404 13412 13132
rect 13468 12962 13524 13916
rect 13692 13186 13748 14364
rect 13692 13134 13694 13186
rect 13746 13134 13748 13186
rect 13692 13122 13748 13134
rect 14028 13188 14084 15092
rect 14140 14754 14196 16044
rect 14140 14702 14142 14754
rect 14194 14702 14196 14754
rect 14140 14690 14196 14702
rect 14252 15202 14308 15214
rect 14252 15150 14254 15202
rect 14306 15150 14308 15202
rect 14252 14308 14308 15150
rect 14364 14420 14420 18732
rect 14476 18450 14532 18732
rect 14700 18676 14756 19070
rect 14812 19124 14868 20132
rect 15036 20130 15092 20132
rect 15036 20078 15038 20130
rect 15090 20078 15092 20130
rect 15036 20066 15092 20078
rect 15148 20018 15204 20636
rect 15148 19966 15150 20018
rect 15202 19966 15204 20018
rect 15148 19954 15204 19966
rect 15372 20580 15428 20590
rect 15372 20018 15428 20524
rect 15372 19966 15374 20018
rect 15426 19966 15428 20018
rect 15372 19954 15428 19966
rect 15596 20018 15652 20748
rect 15708 20802 15764 20814
rect 15708 20750 15710 20802
rect 15762 20750 15764 20802
rect 15708 20692 15764 20750
rect 15820 20802 15876 21868
rect 15932 21476 15988 21486
rect 16380 21476 16436 21486
rect 15932 21474 16436 21476
rect 15932 21422 15934 21474
rect 15986 21422 16382 21474
rect 16434 21422 16436 21474
rect 15932 21420 16436 21422
rect 15932 21410 15988 21420
rect 16380 21364 16436 21420
rect 16380 21298 16436 21308
rect 15820 20750 15822 20802
rect 15874 20750 15876 20802
rect 15820 20738 15876 20750
rect 15708 20626 15764 20636
rect 15596 19966 15598 20018
rect 15650 19966 15652 20018
rect 15596 19954 15652 19966
rect 16268 20468 16324 20478
rect 15198 19628 15462 19638
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15198 19562 15462 19572
rect 15596 19460 15652 19470
rect 15036 19124 15092 19134
rect 14812 19122 15092 19124
rect 14812 19070 15038 19122
rect 15090 19070 15092 19122
rect 14812 19068 15092 19070
rect 14700 18610 14756 18620
rect 14476 18398 14478 18450
rect 14530 18398 14532 18450
rect 14476 18386 14532 18398
rect 14812 18562 14868 18574
rect 14812 18510 14814 18562
rect 14866 18510 14868 18562
rect 14700 17892 14756 17902
rect 14812 17892 14868 18510
rect 14700 17890 14812 17892
rect 14700 17838 14702 17890
rect 14754 17838 14812 17890
rect 14700 17836 14812 17838
rect 14588 17108 14644 17118
rect 14476 15874 14532 15886
rect 14476 15822 14478 15874
rect 14530 15822 14532 15874
rect 14476 15540 14532 15822
rect 14588 15540 14644 17052
rect 14700 16882 14756 17836
rect 14812 17826 14868 17836
rect 14812 17668 14868 17678
rect 14812 17574 14868 17612
rect 14700 16830 14702 16882
rect 14754 16830 14756 16882
rect 14700 16818 14756 16830
rect 14812 16658 14868 16670
rect 14812 16606 14814 16658
rect 14866 16606 14868 16658
rect 14812 16548 14868 16606
rect 14812 16482 14868 16492
rect 14924 16098 14980 19068
rect 15036 19058 15092 19068
rect 15596 19122 15652 19404
rect 15596 19070 15598 19122
rect 15650 19070 15652 19122
rect 15596 19058 15652 19070
rect 15932 19124 15988 19134
rect 15932 19030 15988 19068
rect 16268 19122 16324 20412
rect 16380 20020 16436 20030
rect 16380 19926 16436 19964
rect 16268 19070 16270 19122
rect 16322 19070 16324 19122
rect 16268 19058 16324 19070
rect 15372 19012 15428 19022
rect 15372 18450 15428 18956
rect 15372 18398 15374 18450
rect 15426 18398 15428 18450
rect 15372 18340 15428 18398
rect 15372 18274 15428 18284
rect 16156 18338 16212 18350
rect 16156 18286 16158 18338
rect 16210 18286 16212 18338
rect 15260 18228 15316 18238
rect 16044 18228 16100 18238
rect 15036 18226 15316 18228
rect 15036 18174 15262 18226
rect 15314 18174 15316 18226
rect 15036 18172 15316 18174
rect 15036 17892 15092 18172
rect 15260 18162 15316 18172
rect 15708 18226 16100 18228
rect 15708 18174 16046 18226
rect 16098 18174 16100 18226
rect 15708 18172 16100 18174
rect 15198 18060 15462 18070
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15198 17994 15462 18004
rect 15484 17892 15540 17902
rect 15036 17836 15204 17892
rect 15148 17780 15204 17836
rect 15148 17714 15204 17724
rect 14924 16046 14926 16098
rect 14978 16046 14980 16098
rect 14588 15484 14756 15540
rect 14476 15474 14532 15484
rect 14588 15316 14644 15326
rect 14476 15314 14644 15316
rect 14476 15262 14590 15314
rect 14642 15262 14644 15314
rect 14476 15260 14644 15262
rect 14476 15202 14532 15260
rect 14588 15250 14644 15260
rect 14476 15150 14478 15202
rect 14530 15150 14532 15202
rect 14476 15138 14532 15150
rect 14588 14420 14644 14430
rect 14364 14364 14588 14420
rect 14140 13188 14196 13198
rect 14084 13186 14196 13188
rect 14084 13134 14142 13186
rect 14194 13134 14196 13186
rect 14084 13132 14196 13134
rect 14028 13094 14084 13132
rect 14140 13122 14196 13132
rect 13468 12910 13470 12962
rect 13522 12910 13524 12962
rect 13468 12898 13524 12910
rect 13916 12964 13972 12974
rect 13916 12870 13972 12908
rect 13580 12740 13636 12750
rect 13580 12646 13636 12684
rect 14252 12516 14308 14252
rect 14588 13858 14644 14364
rect 14588 13806 14590 13858
rect 14642 13806 14644 13858
rect 14588 13794 14644 13806
rect 14364 13636 14420 13646
rect 14364 13542 14420 13580
rect 14700 12964 14756 15484
rect 14924 15426 14980 16046
rect 15036 17666 15092 17678
rect 15036 17614 15038 17666
rect 15090 17614 15092 17666
rect 15036 16884 15092 17614
rect 15484 17666 15540 17836
rect 15484 17614 15486 17666
rect 15538 17614 15540 17666
rect 15148 17554 15204 17566
rect 15148 17502 15150 17554
rect 15202 17502 15204 17554
rect 15148 16996 15204 17502
rect 15148 16930 15204 16940
rect 15036 15988 15092 16828
rect 15484 16882 15540 17614
rect 15708 17890 15764 18172
rect 16044 18162 16100 18172
rect 16156 18228 16212 18286
rect 15708 17838 15710 17890
rect 15762 17838 15764 17890
rect 15708 17556 15764 17838
rect 16156 17780 16212 18172
rect 16156 17714 16212 17724
rect 15708 17490 15764 17500
rect 15932 17666 15988 17678
rect 15932 17614 15934 17666
rect 15986 17614 15988 17666
rect 15596 17444 15652 17454
rect 15596 17350 15652 17388
rect 15484 16830 15486 16882
rect 15538 16830 15540 16882
rect 15484 16818 15540 16830
rect 15932 16884 15988 17614
rect 16492 17444 16548 22988
rect 16604 22370 16660 23100
rect 16716 23090 16772 23100
rect 16604 22318 16606 22370
rect 16658 22318 16660 22370
rect 16604 20916 16660 22318
rect 16716 21924 16772 21934
rect 16716 21810 16772 21868
rect 16716 21758 16718 21810
rect 16770 21758 16772 21810
rect 16716 21746 16772 21758
rect 16828 21474 16884 21486
rect 16828 21422 16830 21474
rect 16882 21422 16884 21474
rect 16828 21364 16884 21422
rect 16828 21298 16884 21308
rect 16604 20860 16772 20916
rect 16604 20692 16660 20702
rect 16604 20598 16660 20636
rect 16604 19124 16660 19134
rect 16604 18564 16660 19068
rect 16604 17666 16660 18508
rect 16604 17614 16606 17666
rect 16658 17614 16660 17666
rect 16604 17602 16660 17614
rect 16492 17388 16660 17444
rect 16492 16996 16548 17006
rect 15932 16790 15988 16828
rect 16156 16940 16492 16996
rect 15148 16772 15204 16782
rect 15148 16678 15204 16716
rect 15708 16658 15764 16670
rect 15708 16606 15710 16658
rect 15762 16606 15764 16658
rect 15198 16492 15462 16502
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15198 16426 15462 16436
rect 15484 16324 15540 16334
rect 15708 16324 15764 16606
rect 15484 16322 15764 16324
rect 15484 16270 15486 16322
rect 15538 16270 15764 16322
rect 15484 16268 15764 16270
rect 16044 16658 16100 16670
rect 16044 16606 16046 16658
rect 16098 16606 16100 16658
rect 15484 16212 15540 16268
rect 15484 16146 15540 16156
rect 15148 15988 15204 15998
rect 15036 15986 15204 15988
rect 15036 15934 15150 15986
rect 15202 15934 15204 15986
rect 15036 15932 15204 15934
rect 15148 15922 15204 15932
rect 15596 15986 15652 15998
rect 15932 15988 15988 15998
rect 15596 15934 15598 15986
rect 15650 15934 15652 15986
rect 15596 15540 15652 15934
rect 15820 15986 15988 15988
rect 15820 15934 15934 15986
rect 15986 15934 15988 15986
rect 15820 15932 15988 15934
rect 15820 15764 15876 15932
rect 15932 15922 15988 15932
rect 16044 15764 16100 16606
rect 15820 15698 15876 15708
rect 15932 15708 16100 15764
rect 15596 15474 15652 15484
rect 14924 15374 14926 15426
rect 14978 15374 14980 15426
rect 14924 15362 14980 15374
rect 15260 15426 15316 15438
rect 15260 15374 15262 15426
rect 15314 15374 15316 15426
rect 15260 15092 15316 15374
rect 15036 15036 15316 15092
rect 15036 14756 15092 15036
rect 15198 14924 15462 14934
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15198 14858 15462 14868
rect 15036 14700 15204 14756
rect 14812 14530 14868 14542
rect 14812 14478 14814 14530
rect 14866 14478 14868 14530
rect 14812 13860 14868 14478
rect 14924 14532 14980 14542
rect 14924 14438 14980 14476
rect 15148 14530 15204 14700
rect 15148 14478 15150 14530
rect 15202 14478 15204 14530
rect 14924 13860 14980 13870
rect 14812 13858 14980 13860
rect 14812 13806 14926 13858
rect 14978 13806 14980 13858
rect 14812 13804 14980 13806
rect 14812 13188 14868 13804
rect 14924 13794 14980 13804
rect 15148 13636 15204 14478
rect 15596 14532 15652 14542
rect 15596 14438 15652 14476
rect 14812 13122 14868 13132
rect 14924 13580 15204 13636
rect 15260 14418 15316 14430
rect 15260 14366 15262 14418
rect 15314 14366 15316 14418
rect 14588 12908 14756 12964
rect 14924 12964 14980 13580
rect 15260 13524 15316 14366
rect 15708 14418 15764 14430
rect 15708 14366 15710 14418
rect 15762 14366 15764 14418
rect 15708 14308 15764 14366
rect 15708 14242 15764 14252
rect 15708 13636 15764 13646
rect 15708 13542 15764 13580
rect 14588 12740 14644 12908
rect 14924 12870 14980 12908
rect 15036 13468 15316 13524
rect 15596 13522 15652 13534
rect 15596 13470 15598 13522
rect 15650 13470 15652 13522
rect 14252 12450 14308 12460
rect 14476 12684 14644 12740
rect 14812 12850 14868 12862
rect 14812 12798 14814 12850
rect 14866 12798 14868 12850
rect 13356 12178 13412 12348
rect 13804 12292 13860 12302
rect 13804 12198 13860 12236
rect 13356 12126 13358 12178
rect 13410 12126 13412 12178
rect 13356 12114 13412 12126
rect 13468 12180 13524 12190
rect 13468 12086 13524 12124
rect 14028 12180 14084 12190
rect 14028 12086 14084 12124
rect 13804 11956 13860 11966
rect 13692 11396 13748 11406
rect 13692 11302 13748 11340
rect 13468 11170 13524 11182
rect 13468 11118 13470 11170
rect 13522 11118 13524 11170
rect 13468 8484 13524 11118
rect 13468 8418 13524 8428
rect 13244 7298 13300 7308
rect 12348 3502 12350 3554
rect 12402 3502 12404 3554
rect 12348 3490 12404 3502
rect 13692 3556 13748 3566
rect 13804 3556 13860 11900
rect 13692 3554 13860 3556
rect 13692 3502 13694 3554
rect 13746 3502 13860 3554
rect 13692 3500 13860 3502
rect 14476 3556 14532 12684
rect 14812 12292 14868 12798
rect 13692 3490 13748 3500
rect 14476 3490 14532 3500
rect 14588 12236 14868 12292
rect 13356 3444 13412 3454
rect 13356 3442 13524 3444
rect 13356 3390 13358 3442
rect 13410 3390 13524 3442
rect 13356 3388 13524 3390
rect 13356 3378 13412 3388
rect 10108 3276 10500 3332
rect 10556 3332 10612 3342
rect 11228 3332 11284 3342
rect 11900 3332 11956 3342
rect 12572 3332 12628 3342
rect 10556 3330 10948 3332
rect 10556 3278 10558 3330
rect 10610 3278 10948 3330
rect 10556 3276 10948 3278
rect 10108 800 10164 3276
rect 10556 3266 10612 3276
rect 10536 3164 10800 3174
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10536 3098 10800 3108
rect 10892 1652 10948 3276
rect 11228 3330 11508 3332
rect 11228 3278 11230 3330
rect 11282 3278 11508 3330
rect 11228 3276 11508 3278
rect 11228 3266 11284 3276
rect 10780 1596 10948 1652
rect 10780 800 10836 1596
rect 11452 800 11508 3276
rect 11900 3330 12180 3332
rect 11900 3278 11902 3330
rect 11954 3278 12180 3330
rect 11900 3276 12180 3278
rect 11900 3266 11956 3276
rect 12124 800 12180 3276
rect 12572 3330 12852 3332
rect 12572 3278 12574 3330
rect 12626 3278 12852 3330
rect 12572 3276 12852 3278
rect 12572 3266 12628 3276
rect 12796 800 12852 3276
rect 13468 800 13524 3388
rect 14364 3442 14420 3454
rect 14364 3390 14366 3442
rect 14418 3390 14420 3442
rect 14364 3388 14420 3390
rect 14588 3388 14644 12236
rect 15036 12180 15092 13468
rect 15198 13356 15462 13366
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15198 13290 15462 13300
rect 15260 13188 15316 13198
rect 15316 13132 15540 13188
rect 15260 13094 15316 13132
rect 15148 12962 15204 12974
rect 15148 12910 15150 12962
rect 15202 12910 15204 12962
rect 15148 12852 15204 12910
rect 15148 12786 15204 12796
rect 15372 12964 15428 12974
rect 15372 12292 15428 12908
rect 14812 12124 15092 12180
rect 15148 12236 15428 12292
rect 14812 3556 14868 12124
rect 14924 11954 14980 11966
rect 14924 11902 14926 11954
rect 14978 11902 14980 11954
rect 14924 11508 14980 11902
rect 15036 11956 15092 11966
rect 15148 11956 15204 12236
rect 15484 12178 15540 13132
rect 15596 13076 15652 13470
rect 15932 13412 15988 15708
rect 16044 15540 16100 15550
rect 16156 15540 16212 16940
rect 16492 16902 16548 16940
rect 16604 16772 16660 17388
rect 16492 16716 16660 16772
rect 16380 16660 16436 16670
rect 16380 16566 16436 16604
rect 16268 15876 16324 15886
rect 16268 15782 16324 15820
rect 16492 15764 16548 16716
rect 16716 16100 16772 20860
rect 16828 20804 16884 20814
rect 16940 20804 16996 25452
rect 17052 24164 17108 26348
rect 17164 26338 17220 26348
rect 17500 26404 17556 26414
rect 17500 26310 17556 26348
rect 17948 25620 18004 26572
rect 18060 26516 18116 27244
rect 18172 27074 18228 27692
rect 18172 27022 18174 27074
rect 18226 27022 18228 27074
rect 18172 27010 18228 27022
rect 18172 26516 18228 26526
rect 18060 26514 18228 26516
rect 18060 26462 18174 26514
rect 18226 26462 18228 26514
rect 18060 26460 18228 26462
rect 18172 26450 18228 26460
rect 17388 25508 17444 25518
rect 17388 25414 17444 25452
rect 17948 25506 18004 25564
rect 17948 25454 17950 25506
rect 18002 25454 18004 25506
rect 17948 25442 18004 25454
rect 17612 25396 17668 25406
rect 17164 25282 17220 25294
rect 17164 25230 17166 25282
rect 17218 25230 17220 25282
rect 17164 24724 17220 25230
rect 17388 24948 17444 24958
rect 17612 24948 17668 25340
rect 17724 25394 17780 25406
rect 17724 25342 17726 25394
rect 17778 25342 17780 25394
rect 17724 25172 17780 25342
rect 17724 25106 17780 25116
rect 17948 25172 18004 25182
rect 17612 24892 17780 24948
rect 17388 24854 17444 24892
rect 17164 24658 17220 24668
rect 17612 24724 17668 24734
rect 17612 24630 17668 24668
rect 17612 24388 17668 24398
rect 17052 24108 17556 24164
rect 17276 23940 17332 23950
rect 16828 20802 16996 20804
rect 16828 20750 16830 20802
rect 16882 20750 16996 20802
rect 16828 20748 16996 20750
rect 17052 23938 17332 23940
rect 17052 23886 17278 23938
rect 17330 23886 17332 23938
rect 17052 23884 17332 23886
rect 16828 20468 16884 20748
rect 16828 20402 16884 20412
rect 17052 20244 17108 23884
rect 17276 23874 17332 23884
rect 17388 23940 17444 23950
rect 17388 23826 17444 23884
rect 17388 23774 17390 23826
rect 17442 23774 17444 23826
rect 17388 23762 17444 23774
rect 17388 23156 17444 23166
rect 17388 23062 17444 23100
rect 17276 22148 17332 22158
rect 17164 22092 17276 22148
rect 17164 20356 17220 22092
rect 17276 22054 17332 22092
rect 17388 21588 17444 21598
rect 17388 21494 17444 21532
rect 17388 21028 17444 21038
rect 17388 20914 17444 20972
rect 17388 20862 17390 20914
rect 17442 20862 17444 20914
rect 17388 20692 17444 20862
rect 17388 20626 17444 20636
rect 17276 20580 17332 20590
rect 17276 20486 17332 20524
rect 17164 20300 17332 20356
rect 17052 20188 17220 20244
rect 16940 20132 16996 20142
rect 16828 20020 16884 20030
rect 16828 19926 16884 19964
rect 16940 19796 16996 20076
rect 16828 19740 16996 19796
rect 16828 18674 16884 19740
rect 17164 19348 17220 20188
rect 17276 19908 17332 20300
rect 17500 20132 17556 24108
rect 17612 20468 17668 24332
rect 17724 23828 17780 24892
rect 17724 23734 17780 23772
rect 17836 23940 17892 23950
rect 17948 23940 18004 25116
rect 18284 24724 18340 27806
rect 18396 27970 18452 28028
rect 18396 27918 18398 27970
rect 18450 27918 18452 27970
rect 18396 26964 18452 27918
rect 18620 27860 18676 28140
rect 18508 27858 18676 27860
rect 18508 27806 18622 27858
rect 18674 27806 18676 27858
rect 18508 27804 18676 27806
rect 18508 27076 18564 27804
rect 18620 27794 18676 27804
rect 18508 26982 18564 27020
rect 18396 26898 18452 26908
rect 18396 26290 18452 26302
rect 18396 26238 18398 26290
rect 18450 26238 18452 26290
rect 18396 25730 18452 26238
rect 18396 25678 18398 25730
rect 18450 25678 18452 25730
rect 18396 25666 18452 25678
rect 17836 23938 18004 23940
rect 17836 23886 17838 23938
rect 17890 23886 18004 23938
rect 17836 23884 18004 23886
rect 18060 24668 18340 24724
rect 17724 23380 17780 23390
rect 17836 23380 17892 23884
rect 17724 23378 17892 23380
rect 17724 23326 17726 23378
rect 17778 23326 17892 23378
rect 17724 23324 17892 23326
rect 17948 23492 18004 23502
rect 17724 23314 17780 23324
rect 17836 22594 17892 22606
rect 17836 22542 17838 22594
rect 17890 22542 17892 22594
rect 17836 22482 17892 22542
rect 17836 22430 17838 22482
rect 17890 22430 17892 22482
rect 17836 22418 17892 22430
rect 17724 21812 17780 21822
rect 17724 21718 17780 21756
rect 17948 21588 18004 23436
rect 18060 23268 18116 24668
rect 18396 24612 18452 24622
rect 18284 24500 18340 24510
rect 18284 24406 18340 24444
rect 18396 24276 18452 24556
rect 18172 24220 18452 24276
rect 18172 23940 18228 24220
rect 18732 24164 18788 28252
rect 19068 27860 19124 27870
rect 19516 27860 19572 27870
rect 19068 27858 19572 27860
rect 19068 27806 19070 27858
rect 19122 27806 19518 27858
rect 19570 27806 19572 27858
rect 19068 27804 19572 27806
rect 19068 27794 19124 27804
rect 19516 27794 19572 27804
rect 18956 26964 19012 26974
rect 19404 26964 19460 26974
rect 18956 26962 19460 26964
rect 18956 26910 18958 26962
rect 19010 26910 19406 26962
rect 19458 26910 19460 26962
rect 18956 26908 19460 26910
rect 18956 26898 19012 26908
rect 19404 26898 19460 26908
rect 19180 26404 19236 26414
rect 19180 26310 19236 26348
rect 18844 26290 18900 26302
rect 18844 26238 18846 26290
rect 18898 26238 18900 26290
rect 18844 25620 18900 26238
rect 19516 26178 19572 26190
rect 19516 26126 19518 26178
rect 19570 26126 19572 26178
rect 19516 26068 19572 26126
rect 19516 26002 19572 26012
rect 18956 25732 19012 25742
rect 18956 25638 19012 25676
rect 18844 25526 18900 25564
rect 19628 25508 19684 29260
rect 19740 28084 19796 36316
rect 19852 36306 19908 36316
rect 20188 36370 20244 39200
rect 20188 36318 20190 36370
rect 20242 36318 20244 36370
rect 20188 36306 20244 36318
rect 20748 36372 20804 36382
rect 20860 36372 20916 39200
rect 21084 36372 21140 36382
rect 20860 36370 21140 36372
rect 20860 36318 21086 36370
rect 21138 36318 21140 36370
rect 20860 36316 21140 36318
rect 19860 36092 20124 36102
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 19860 36026 20124 36036
rect 19860 34524 20124 34534
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 19860 34458 20124 34468
rect 19860 32956 20124 32966
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 19860 32890 20124 32900
rect 19860 31388 20124 31398
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 19860 31322 20124 31332
rect 19860 29820 20124 29830
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 19860 29754 20124 29764
rect 19964 29540 20020 29550
rect 19964 29446 20020 29484
rect 20300 29538 20356 29550
rect 20300 29486 20302 29538
rect 20354 29486 20356 29538
rect 20300 29316 20356 29486
rect 20300 29250 20356 29260
rect 19852 28644 19908 28654
rect 19852 28642 20244 28644
rect 19852 28590 19854 28642
rect 19906 28590 20244 28642
rect 19852 28588 20244 28590
rect 19852 28578 19908 28588
rect 19860 28252 20124 28262
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 19860 28186 20124 28196
rect 19852 28084 19908 28094
rect 19740 28082 19908 28084
rect 19740 28030 19854 28082
rect 19906 28030 19908 28082
rect 19740 28028 19908 28030
rect 19852 28018 19908 28028
rect 20188 27970 20244 28588
rect 20188 27918 20190 27970
rect 20242 27918 20244 27970
rect 20188 27748 20244 27918
rect 20524 27972 20580 27982
rect 20524 27878 20580 27916
rect 19740 27300 19796 27310
rect 19740 26962 19796 27244
rect 20188 27186 20244 27692
rect 20188 27134 20190 27186
rect 20242 27134 20244 27186
rect 20188 27122 20244 27134
rect 19740 26910 19742 26962
rect 19794 26910 19796 26962
rect 19740 26898 19796 26910
rect 20412 26852 20468 26862
rect 19860 26684 20124 26694
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 19860 26618 20124 26628
rect 20076 26404 20132 26414
rect 19740 26292 19796 26302
rect 19740 26198 19796 26236
rect 19852 26290 19908 26302
rect 19852 26238 19854 26290
rect 19906 26238 19908 26290
rect 19852 25844 19908 26238
rect 19852 25778 19908 25788
rect 20076 26290 20132 26348
rect 20076 26238 20078 26290
rect 20130 26238 20132 26290
rect 19292 25452 19684 25508
rect 20076 25508 20132 26238
rect 18956 24724 19012 24734
rect 18956 24630 19012 24668
rect 18844 24498 18900 24510
rect 18844 24446 18846 24498
rect 18898 24446 18900 24498
rect 18844 24276 18900 24446
rect 19180 24500 19236 24510
rect 19180 24406 19236 24444
rect 18844 24220 19012 24276
rect 18732 24108 18900 24164
rect 18172 23874 18228 23884
rect 18284 23940 18340 23950
rect 18732 23940 18788 23950
rect 18284 23938 18788 23940
rect 18284 23886 18286 23938
rect 18338 23886 18734 23938
rect 18786 23886 18788 23938
rect 18284 23884 18788 23886
rect 18284 23874 18340 23884
rect 18732 23874 18788 23884
rect 18508 23716 18564 23726
rect 18844 23716 18900 24108
rect 18508 23714 18900 23716
rect 18508 23662 18510 23714
rect 18562 23662 18900 23714
rect 18508 23660 18900 23662
rect 18956 23716 19012 24220
rect 19180 23828 19236 23838
rect 19292 23828 19348 25452
rect 20076 25442 20132 25452
rect 20300 26068 20356 26078
rect 20188 25396 20244 25406
rect 19180 23826 19348 23828
rect 19180 23774 19182 23826
rect 19234 23774 19348 23826
rect 19180 23772 19348 23774
rect 19404 25282 19460 25294
rect 19404 25230 19406 25282
rect 19458 25230 19460 25282
rect 19404 24610 19460 25230
rect 20076 25284 20132 25322
rect 20188 25284 20244 25340
rect 20132 25228 20244 25284
rect 20076 25218 20132 25228
rect 19860 25116 20124 25126
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 19860 25050 20124 25060
rect 19404 24558 19406 24610
rect 19458 24558 19460 24610
rect 19180 23762 19236 23772
rect 18508 23650 18564 23660
rect 18172 23268 18228 23278
rect 18060 23212 18172 23268
rect 18060 22930 18116 22942
rect 18060 22878 18062 22930
rect 18114 22878 18116 22930
rect 18060 22036 18116 22878
rect 18172 22594 18228 23212
rect 18172 22542 18174 22594
rect 18226 22542 18228 22594
rect 18172 22530 18228 22542
rect 18284 23156 18340 23166
rect 18284 22482 18340 23100
rect 18844 23156 18900 23166
rect 18956 23156 19012 23660
rect 18844 23154 19012 23156
rect 18844 23102 18846 23154
rect 18898 23102 19012 23154
rect 18844 23100 19012 23102
rect 19292 23604 19348 23614
rect 18844 23090 18900 23100
rect 18620 23044 18676 23054
rect 18620 22594 18676 22988
rect 19180 23044 19236 23054
rect 19180 22950 19236 22988
rect 18956 22932 19012 22942
rect 18956 22838 19012 22876
rect 18620 22542 18622 22594
rect 18674 22542 18676 22594
rect 18620 22530 18676 22542
rect 18284 22430 18286 22482
rect 18338 22430 18340 22482
rect 18284 22418 18340 22430
rect 18732 22258 18788 22270
rect 18732 22206 18734 22258
rect 18786 22206 18788 22258
rect 18732 22148 18788 22206
rect 18732 22082 18788 22092
rect 18060 21970 18116 21980
rect 19292 21810 19348 23548
rect 19404 23156 19460 24558
rect 20188 24722 20244 24734
rect 20188 24670 20190 24722
rect 20242 24670 20244 24722
rect 20188 24612 20244 24670
rect 20188 24546 20244 24556
rect 19516 24498 19572 24510
rect 19516 24446 19518 24498
rect 19570 24446 19572 24498
rect 19516 23938 19572 24446
rect 19516 23886 19518 23938
rect 19570 23886 19572 23938
rect 19516 23874 19572 23886
rect 20300 23716 20356 26012
rect 20412 24612 20468 26796
rect 20524 26066 20580 26078
rect 20524 26014 20526 26066
rect 20578 26014 20580 26066
rect 20524 25506 20580 26014
rect 20524 25454 20526 25506
rect 20578 25454 20580 25506
rect 20524 25442 20580 25454
rect 20748 25394 20804 36316
rect 21084 36306 21140 36316
rect 21420 36370 21476 36382
rect 21420 36318 21422 36370
rect 21474 36318 21476 36370
rect 20972 29314 21028 29326
rect 20972 29262 20974 29314
rect 21026 29262 21028 29314
rect 20972 27972 21028 29262
rect 21196 29204 21252 29214
rect 21196 29110 21252 29148
rect 20972 27906 21028 27916
rect 21308 26292 21364 26302
rect 21308 26198 21364 26236
rect 20748 25342 20750 25394
rect 20802 25342 20804 25394
rect 20748 25330 20804 25342
rect 21196 26180 21252 26190
rect 20524 24836 20580 24846
rect 20972 24836 21028 24846
rect 20524 24834 21028 24836
rect 20524 24782 20526 24834
rect 20578 24782 20974 24834
rect 21026 24782 21028 24834
rect 20524 24780 21028 24782
rect 20524 24770 20580 24780
rect 20860 24612 20916 24622
rect 20412 24610 20916 24612
rect 20412 24558 20862 24610
rect 20914 24558 20916 24610
rect 20412 24556 20916 24558
rect 20188 23660 20356 23716
rect 19860 23548 20124 23558
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 19860 23482 20124 23492
rect 19404 23062 19460 23100
rect 19628 23380 19684 23390
rect 19516 22930 19572 22942
rect 19516 22878 19518 22930
rect 19570 22878 19572 22930
rect 19404 22372 19460 22382
rect 19516 22372 19572 22878
rect 19404 22370 19572 22372
rect 19404 22318 19406 22370
rect 19458 22318 19572 22370
rect 19404 22316 19572 22318
rect 19404 22306 19460 22316
rect 19628 22258 19684 23324
rect 19964 23268 20020 23278
rect 19964 23174 20020 23212
rect 19628 22206 19630 22258
rect 19682 22206 19684 22258
rect 19628 22194 19684 22206
rect 20076 22148 20132 22186
rect 20076 22082 20132 22092
rect 19860 21980 20124 21990
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 19860 21914 20124 21924
rect 19292 21758 19294 21810
rect 19346 21758 19348 21810
rect 19292 21746 19348 21758
rect 18508 21698 18564 21710
rect 18508 21646 18510 21698
rect 18562 21646 18564 21698
rect 18060 21588 18116 21598
rect 17948 21586 18116 21588
rect 17948 21534 18062 21586
rect 18114 21534 18116 21586
rect 17948 21532 18116 21534
rect 17724 20916 17780 20926
rect 17724 20822 17780 20860
rect 17836 20692 17892 20702
rect 17836 20690 18004 20692
rect 17836 20638 17838 20690
rect 17890 20638 18004 20690
rect 17836 20636 18004 20638
rect 17836 20626 17892 20636
rect 17612 20412 17780 20468
rect 17500 20038 17556 20076
rect 17612 20244 17668 20254
rect 17276 19852 17556 19908
rect 16940 19292 17220 19348
rect 16940 19122 16996 19292
rect 16940 19070 16942 19122
rect 16994 19070 16996 19122
rect 16940 19058 16996 19070
rect 16828 18622 16830 18674
rect 16882 18622 16884 18674
rect 16828 16884 16884 18622
rect 17052 17556 17108 19292
rect 17276 19122 17332 19134
rect 17276 19070 17278 19122
rect 17330 19070 17332 19122
rect 17276 18564 17332 19070
rect 17276 18498 17332 18508
rect 17052 17490 17108 17500
rect 16940 17442 16996 17454
rect 16940 17390 16942 17442
rect 16994 17390 16996 17442
rect 16940 16996 16996 17390
rect 17388 17442 17444 17454
rect 17388 17390 17390 17442
rect 17442 17390 17444 17442
rect 17388 17108 17444 17390
rect 17500 17332 17556 19852
rect 17612 18450 17668 20188
rect 17724 19236 17780 20412
rect 17836 20132 17892 20142
rect 17836 20038 17892 20076
rect 17948 20020 18004 20636
rect 17948 19954 18004 19964
rect 17836 19236 17892 19246
rect 17724 19234 17892 19236
rect 17724 19182 17838 19234
rect 17890 19182 17892 19234
rect 17724 19180 17892 19182
rect 17836 19124 17892 19180
rect 17836 19058 17892 19068
rect 18060 18674 18116 21532
rect 18284 21586 18340 21598
rect 18284 21534 18286 21586
rect 18338 21534 18340 21586
rect 18284 21364 18340 21534
rect 18284 21298 18340 21308
rect 18508 20916 18564 21646
rect 18844 21588 18900 21598
rect 18844 21586 19012 21588
rect 18844 21534 18846 21586
rect 18898 21534 19012 21586
rect 18844 21532 19012 21534
rect 18844 21522 18900 21532
rect 18508 20860 18788 20916
rect 18396 20802 18452 20814
rect 18396 20750 18398 20802
rect 18450 20750 18452 20802
rect 18396 19908 18452 20750
rect 18732 20804 18788 20860
rect 18956 20804 19012 21532
rect 19516 21586 19572 21598
rect 19964 21588 20020 21598
rect 19516 21534 19518 21586
rect 19570 21534 19572 21586
rect 19068 21476 19124 21486
rect 19516 21476 19572 21534
rect 19068 21474 19572 21476
rect 19068 21422 19070 21474
rect 19122 21422 19572 21474
rect 19068 21420 19572 21422
rect 19628 21586 20020 21588
rect 19628 21534 19966 21586
rect 20018 21534 20020 21586
rect 19628 21532 20020 21534
rect 19068 21410 19124 21420
rect 19628 21140 19684 21532
rect 19964 21522 20020 21532
rect 19404 21084 19684 21140
rect 19404 21026 19460 21084
rect 19404 20974 19406 21026
rect 19458 20974 19460 21026
rect 19404 20962 19460 20974
rect 19068 20804 19124 20814
rect 18732 20802 18900 20804
rect 18732 20750 18734 20802
rect 18786 20750 18900 20802
rect 18732 20748 18900 20750
rect 18956 20802 19124 20804
rect 18956 20750 19070 20802
rect 19122 20750 19124 20802
rect 18956 20748 19124 20750
rect 18732 20738 18788 20748
rect 18508 20692 18564 20702
rect 18508 20244 18564 20636
rect 18508 20178 18564 20188
rect 18844 20130 18900 20748
rect 18844 20078 18846 20130
rect 18898 20078 18900 20130
rect 18732 20020 18788 20030
rect 18732 19926 18788 19964
rect 18508 19908 18564 19918
rect 18396 19906 18564 19908
rect 18396 19854 18510 19906
rect 18562 19854 18564 19906
rect 18396 19852 18564 19854
rect 18172 19236 18228 19246
rect 18172 19122 18228 19180
rect 18172 19070 18174 19122
rect 18226 19070 18228 19122
rect 18172 19058 18228 19070
rect 18508 19234 18564 19852
rect 18508 19182 18510 19234
rect 18562 19182 18564 19234
rect 18060 18622 18062 18674
rect 18114 18622 18116 18674
rect 18060 18610 18116 18622
rect 17612 18398 17614 18450
rect 17666 18398 17668 18450
rect 17612 18386 17668 18398
rect 18396 18452 18452 18462
rect 18396 18358 18452 18396
rect 18508 18228 18564 19182
rect 18844 19236 18900 20078
rect 18844 19142 18900 19180
rect 19068 20132 19124 20748
rect 19852 20692 19908 20702
rect 19516 20690 19908 20692
rect 19516 20638 19854 20690
rect 19906 20638 19908 20690
rect 19516 20636 19908 20638
rect 19516 20242 19572 20636
rect 19852 20626 19908 20636
rect 20188 20690 20244 23660
rect 20860 23604 20916 24556
rect 20972 24612 21028 24780
rect 20972 24546 21028 24556
rect 21196 24834 21252 26124
rect 21420 26068 21476 36318
rect 21532 36372 21588 39200
rect 21756 36372 21812 36382
rect 21532 36370 21812 36372
rect 21532 36318 21758 36370
rect 21810 36318 21812 36370
rect 21532 36316 21812 36318
rect 21756 36306 21812 36316
rect 22092 36372 22148 36382
rect 22204 36372 22260 39200
rect 22652 36482 22708 36494
rect 22652 36430 22654 36482
rect 22706 36430 22708 36482
rect 22428 36372 22484 36382
rect 22204 36370 22484 36372
rect 22204 36318 22430 36370
rect 22482 36318 22484 36370
rect 22204 36316 22484 36318
rect 22092 36278 22148 36316
rect 22428 36306 22484 36316
rect 22428 35476 22484 35486
rect 21756 33124 21812 33134
rect 21532 30210 21588 30222
rect 21532 30158 21534 30210
rect 21586 30158 21588 30210
rect 21532 29650 21588 30158
rect 21756 30098 21812 33068
rect 22092 30100 22148 30110
rect 21756 30046 21758 30098
rect 21810 30046 21812 30098
rect 21756 30034 21812 30046
rect 21868 30098 22148 30100
rect 21868 30046 22094 30098
rect 22146 30046 22148 30098
rect 21868 30044 22148 30046
rect 21532 29598 21534 29650
rect 21586 29598 21588 29650
rect 21532 29586 21588 29598
rect 21868 29650 21924 30044
rect 22092 30034 22148 30044
rect 22428 30098 22484 35420
rect 22652 33124 22708 36430
rect 22876 36372 22932 39200
rect 23548 37828 23604 39200
rect 23548 37772 24164 37828
rect 23324 36484 23380 36494
rect 23212 36482 23380 36484
rect 23212 36430 23326 36482
rect 23378 36430 23380 36482
rect 23212 36428 23380 36430
rect 24108 36484 24164 37772
rect 24220 36708 24276 39200
rect 24892 36932 24948 39200
rect 25564 37828 25620 39200
rect 25564 37772 26180 37828
rect 24522 36876 24786 36886
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24892 36866 24948 36876
rect 25900 36932 25956 36942
rect 24522 36810 24786 36820
rect 24220 36642 24276 36652
rect 25228 36708 25284 36718
rect 24108 36428 24612 36484
rect 23100 36372 23156 36382
rect 22876 36370 23156 36372
rect 22876 36318 23102 36370
rect 23154 36318 23156 36370
rect 22876 36316 23156 36318
rect 23100 36306 23156 36316
rect 22652 33058 22708 33068
rect 22428 30046 22430 30098
rect 22482 30046 22484 30098
rect 22428 30034 22484 30046
rect 21868 29598 21870 29650
rect 21922 29598 21924 29650
rect 21868 29586 21924 29598
rect 21980 29652 22036 29662
rect 21980 29428 22036 29596
rect 22428 29428 22484 29438
rect 21980 29372 22428 29428
rect 21868 29316 21924 29326
rect 21756 28642 21812 28654
rect 21756 28590 21758 28642
rect 21810 28590 21812 28642
rect 21756 27860 21812 28590
rect 21868 28642 21924 29260
rect 21868 28590 21870 28642
rect 21922 28590 21924 28642
rect 21868 28578 21924 28590
rect 21980 28308 22036 29372
rect 22428 29334 22484 29372
rect 22764 29316 22820 29326
rect 22764 29222 22820 29260
rect 22204 29204 22260 29214
rect 22204 29110 22260 29148
rect 22988 29204 23044 29214
rect 22988 29110 23044 29148
rect 22428 28642 22484 28654
rect 22428 28590 22430 28642
rect 22482 28590 22484 28642
rect 22092 28532 22148 28542
rect 22092 28530 22260 28532
rect 22092 28478 22094 28530
rect 22146 28478 22260 28530
rect 22092 28476 22260 28478
rect 22092 28466 22148 28476
rect 21980 28252 22148 28308
rect 21980 27972 22036 27982
rect 21868 27860 21924 27870
rect 21756 27858 21924 27860
rect 21756 27806 21870 27858
rect 21922 27806 21924 27858
rect 21756 27804 21924 27806
rect 21756 27188 21812 27804
rect 21868 27794 21924 27804
rect 21756 27186 21924 27188
rect 21756 27134 21758 27186
rect 21810 27134 21924 27186
rect 21756 27132 21924 27134
rect 21756 26908 21812 27132
rect 21532 26852 21812 26908
rect 21532 26514 21588 26852
rect 21532 26462 21534 26514
rect 21586 26462 21588 26514
rect 21532 26450 21588 26462
rect 21868 26290 21924 27132
rect 21980 27074 22036 27916
rect 22092 27970 22148 28252
rect 22092 27918 22094 27970
rect 22146 27918 22148 27970
rect 22092 27906 22148 27918
rect 22204 27970 22260 28476
rect 22204 27918 22206 27970
rect 22258 27918 22260 27970
rect 21980 27022 21982 27074
rect 22034 27022 22036 27074
rect 21980 27010 22036 27022
rect 22204 26962 22260 27918
rect 22428 27860 22484 28590
rect 22652 28420 22708 28430
rect 22652 28418 22820 28420
rect 22652 28366 22654 28418
rect 22706 28366 22820 28418
rect 22652 28364 22820 28366
rect 22652 28354 22708 28364
rect 22316 27858 22484 27860
rect 22316 27806 22430 27858
rect 22482 27806 22484 27858
rect 22316 27804 22484 27806
rect 22316 27076 22372 27804
rect 22428 27794 22484 27804
rect 22652 27860 22708 27870
rect 22316 27010 22372 27020
rect 22204 26910 22206 26962
rect 22258 26910 22260 26962
rect 22204 26908 22260 26910
rect 22652 26964 22708 27804
rect 22764 27636 22820 28364
rect 23212 28084 23268 36428
rect 23324 36418 23380 36428
rect 23548 36372 23604 36382
rect 23436 33908 23492 33918
rect 23324 30098 23380 30110
rect 23324 30046 23326 30098
rect 23378 30046 23380 30098
rect 23324 29650 23380 30046
rect 23324 29598 23326 29650
rect 23378 29598 23380 29650
rect 23324 29586 23380 29598
rect 23212 28018 23268 28028
rect 23324 28532 23380 28542
rect 22876 27860 22932 27870
rect 23212 27860 23268 27870
rect 22876 27858 23268 27860
rect 22876 27806 22878 27858
rect 22930 27806 23214 27858
rect 23266 27806 23268 27858
rect 22876 27804 23268 27806
rect 22876 27794 22932 27804
rect 23212 27794 23268 27804
rect 22764 27580 23044 27636
rect 22988 27074 23044 27580
rect 22988 27022 22990 27074
rect 23042 27022 23044 27074
rect 22988 27010 23044 27022
rect 22764 26964 22820 26974
rect 22652 26962 22820 26964
rect 22652 26910 22766 26962
rect 22818 26910 22820 26962
rect 22652 26908 22820 26910
rect 22204 26852 22372 26908
rect 22764 26898 22820 26908
rect 23324 26962 23380 28476
rect 23324 26910 23326 26962
rect 23378 26910 23380 26962
rect 23324 26898 23380 26910
rect 21868 26238 21870 26290
rect 21922 26238 21924 26290
rect 21868 26226 21924 26238
rect 21980 26404 22036 26414
rect 21420 26002 21476 26012
rect 21420 25844 21476 25854
rect 21308 25396 21364 25406
rect 21308 25302 21364 25340
rect 21196 24782 21198 24834
rect 21250 24782 21252 24834
rect 21196 24500 21252 24782
rect 21420 24724 21476 25788
rect 21644 25396 21700 25406
rect 21980 25396 22036 26348
rect 21644 25394 22036 25396
rect 21644 25342 21646 25394
rect 21698 25342 22036 25394
rect 21644 25340 22036 25342
rect 22204 26290 22260 26302
rect 22204 26238 22206 26290
rect 22258 26238 22260 26290
rect 21644 25330 21700 25340
rect 21196 24434 21252 24444
rect 21308 24722 21476 24724
rect 21308 24670 21422 24722
rect 21474 24670 21476 24722
rect 21308 24668 21476 24670
rect 20524 23548 20916 23604
rect 21196 23940 21252 23950
rect 20300 23268 20356 23278
rect 20300 23174 20356 23212
rect 20412 22258 20468 22270
rect 20412 22206 20414 22258
rect 20466 22206 20468 22258
rect 20412 22148 20468 22206
rect 20412 22082 20468 22092
rect 20300 21700 20356 21710
rect 20300 21606 20356 21644
rect 20188 20638 20190 20690
rect 20242 20638 20244 20690
rect 20188 20626 20244 20638
rect 20524 20692 20580 23548
rect 20636 23266 20692 23278
rect 20636 23214 20638 23266
rect 20690 23214 20692 23266
rect 20636 22260 20692 23214
rect 20636 22194 20692 22204
rect 20748 22146 20804 22158
rect 20748 22094 20750 22146
rect 20802 22094 20804 22146
rect 20748 22036 20804 22094
rect 21196 22036 21252 23884
rect 21308 23826 21364 24668
rect 21420 24658 21476 24668
rect 21868 24724 21924 24734
rect 22092 24724 22148 24734
rect 21868 24722 22148 24724
rect 21868 24670 21870 24722
rect 21922 24670 22094 24722
rect 22146 24670 22148 24722
rect 21868 24668 22148 24670
rect 21868 24658 21924 24668
rect 22092 24658 22148 24668
rect 21980 24500 22036 24510
rect 21308 23774 21310 23826
rect 21362 23774 21364 23826
rect 21308 23762 21364 23774
rect 21644 23828 21700 23838
rect 21644 23734 21700 23772
rect 21980 23826 22036 24444
rect 22204 24052 22260 26238
rect 22316 24052 22372 26852
rect 23436 26514 23492 33852
rect 23548 28082 23604 36316
rect 24556 36370 24612 36428
rect 24556 36318 24558 36370
rect 24610 36318 24612 36370
rect 24556 36306 24612 36318
rect 24892 36370 24948 36382
rect 24892 36318 24894 36370
rect 24946 36318 24948 36370
rect 23996 35588 24052 35598
rect 23660 33124 23716 33134
rect 23660 30098 23716 33068
rect 23660 30046 23662 30098
rect 23714 30046 23716 30098
rect 23660 30034 23716 30046
rect 23548 28030 23550 28082
rect 23602 28030 23604 28082
rect 23548 28018 23604 28030
rect 23660 29314 23716 29326
rect 23660 29262 23662 29314
rect 23714 29262 23716 29314
rect 23436 26462 23438 26514
rect 23490 26462 23492 26514
rect 23436 26450 23492 26462
rect 23660 26404 23716 29262
rect 23884 29204 23940 29214
rect 23772 29148 23884 29204
rect 23772 28530 23828 29148
rect 23884 29110 23940 29148
rect 23772 28478 23774 28530
rect 23826 28478 23828 28530
rect 23772 28466 23828 28478
rect 23996 28084 24052 35532
rect 24522 35308 24786 35318
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24522 35242 24786 35252
rect 24892 33908 24948 36318
rect 25228 36370 25284 36652
rect 25228 36318 25230 36370
rect 25282 36318 25284 36370
rect 25228 36306 25284 36318
rect 25452 36482 25508 36494
rect 25452 36430 25454 36482
rect 25506 36430 25508 36482
rect 24892 33842 24948 33852
rect 25004 35924 25060 35934
rect 24522 33740 24786 33750
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24522 33674 24786 33684
rect 24522 32172 24786 32182
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24522 32106 24786 32116
rect 24522 30604 24786 30614
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24522 30538 24786 30548
rect 24332 30436 24388 30446
rect 24108 30212 24164 30222
rect 24108 30210 24276 30212
rect 24108 30158 24110 30210
rect 24162 30158 24276 30210
rect 24108 30156 24276 30158
rect 24108 30146 24164 30156
rect 24220 29650 24276 30156
rect 24332 30098 24388 30380
rect 24332 30046 24334 30098
rect 24386 30046 24388 30098
rect 24332 30034 24388 30046
rect 24220 29598 24222 29650
rect 24274 29598 24276 29650
rect 24220 29586 24276 29598
rect 24522 29036 24786 29046
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24522 28970 24786 28980
rect 25004 28868 25060 35868
rect 25452 33124 25508 36430
rect 25900 36370 25956 36876
rect 26124 36708 26180 37772
rect 26236 36932 26292 39200
rect 26908 37492 26964 39200
rect 27580 37828 27636 39200
rect 27580 37772 28196 37828
rect 26908 37436 27188 37492
rect 26236 36866 26292 36876
rect 26124 36652 26628 36708
rect 25900 36318 25902 36370
rect 25954 36318 25956 36370
rect 25900 36306 25956 36318
rect 26236 36372 26292 36382
rect 26236 36278 26292 36316
rect 26572 36370 26628 36652
rect 26796 36484 26852 36494
rect 26572 36318 26574 36370
rect 26626 36318 26628 36370
rect 26572 36306 26628 36318
rect 26684 36482 26852 36484
rect 26684 36430 26798 36482
rect 26850 36430 26852 36482
rect 26684 36428 26852 36430
rect 26684 33908 26740 36428
rect 26796 36418 26852 36428
rect 26236 33852 26740 33908
rect 26796 36260 26852 36270
rect 25452 33058 25508 33068
rect 25788 33572 25844 33582
rect 25564 30212 25620 30222
rect 25564 30210 25732 30212
rect 25564 30158 25566 30210
rect 25618 30158 25732 30210
rect 25564 30156 25732 30158
rect 25564 30146 25620 30156
rect 25676 29652 25732 30156
rect 25788 30098 25844 33516
rect 25788 30046 25790 30098
rect 25842 30046 25844 30098
rect 25788 30034 25844 30046
rect 26124 30098 26180 30110
rect 26124 30046 26126 30098
rect 26178 30046 26180 30098
rect 26124 29988 26180 30046
rect 25900 29932 26180 29988
rect 25788 29652 25844 29662
rect 25676 29650 25844 29652
rect 25676 29598 25790 29650
rect 25842 29598 25844 29650
rect 25676 29596 25844 29598
rect 25788 29586 25844 29596
rect 25228 29314 25284 29326
rect 25900 29316 25956 29932
rect 25228 29262 25230 29314
rect 25282 29262 25284 29314
rect 25228 29092 25284 29262
rect 25564 29260 25956 29316
rect 26124 29764 26180 29774
rect 25452 29204 25508 29214
rect 24780 28812 25060 28868
rect 25116 29036 25284 29092
rect 25340 29148 25452 29204
rect 24108 28532 24164 28542
rect 24780 28532 24836 28812
rect 25004 28644 25060 28654
rect 24108 28530 24388 28532
rect 24108 28478 24110 28530
rect 24162 28478 24388 28530
rect 24108 28476 24388 28478
rect 24108 28466 24164 28476
rect 24220 28084 24276 28094
rect 23996 28082 24276 28084
rect 23996 28030 24222 28082
rect 24274 28030 24276 28082
rect 23996 28028 24276 28030
rect 24220 28018 24276 28028
rect 23884 27860 23940 27870
rect 23884 27766 23940 27804
rect 24108 27860 24164 27870
rect 23660 26338 23716 26348
rect 24108 27076 24164 27804
rect 24108 26402 24164 27020
rect 24108 26350 24110 26402
rect 24162 26350 24164 26402
rect 22428 26290 22484 26302
rect 22428 26238 22430 26290
rect 22482 26238 22484 26290
rect 22428 25172 22484 26238
rect 22876 26292 22932 26302
rect 23100 26292 23156 26302
rect 22876 26290 23156 26292
rect 22876 26238 22878 26290
rect 22930 26238 23102 26290
rect 23154 26238 23156 26290
rect 22876 26236 23156 26238
rect 22876 26226 22932 26236
rect 23100 26226 23156 26236
rect 23772 26292 23828 26302
rect 23828 26236 23940 26292
rect 23772 26198 23828 26236
rect 22764 25732 22820 25742
rect 22764 25638 22820 25676
rect 23324 25732 23380 25742
rect 23324 25638 23380 25676
rect 22428 25106 22484 25116
rect 22876 25506 22932 25518
rect 22876 25454 22878 25506
rect 22930 25454 22932 25506
rect 22876 25172 22932 25454
rect 23100 25508 23156 25518
rect 23100 25506 23268 25508
rect 23100 25454 23102 25506
rect 23154 25454 23268 25506
rect 23100 25452 23268 25454
rect 23100 25442 23156 25452
rect 22428 24948 22484 24958
rect 22428 24854 22484 24892
rect 22876 24612 22932 25116
rect 22876 24556 23156 24612
rect 22876 24388 22932 24398
rect 22316 23996 22596 24052
rect 22204 23986 22260 23996
rect 21980 23774 21982 23826
rect 22034 23774 22036 23826
rect 21980 23762 22036 23774
rect 22316 23826 22372 23838
rect 22316 23774 22318 23826
rect 22370 23774 22372 23826
rect 22316 23604 22372 23774
rect 22316 23538 22372 23548
rect 22540 23492 22596 23996
rect 22652 23716 22708 23726
rect 22652 23622 22708 23660
rect 22540 23436 22708 23492
rect 21308 23042 21364 23054
rect 21308 22990 21310 23042
rect 21362 22990 21364 23042
rect 21308 22484 21364 22990
rect 22652 22596 22708 23436
rect 21868 22540 22708 22596
rect 21308 22428 21588 22484
rect 21532 22372 21588 22428
rect 21644 22372 21700 22382
rect 21532 22370 21700 22372
rect 21532 22318 21646 22370
rect 21698 22318 21700 22370
rect 21532 22316 21700 22318
rect 20748 21980 21252 22036
rect 20972 21586 21028 21598
rect 20972 21534 20974 21586
rect 21026 21534 21028 21586
rect 20972 21364 21028 21534
rect 20748 20916 20804 20926
rect 20972 20916 21028 21308
rect 20748 20914 21028 20916
rect 20748 20862 20750 20914
rect 20802 20862 21028 20914
rect 20748 20860 21028 20862
rect 20748 20850 20804 20860
rect 20524 20636 21028 20692
rect 19860 20412 20124 20422
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 19860 20346 20124 20356
rect 19516 20190 19518 20242
rect 19570 20190 19572 20242
rect 19516 20178 19572 20190
rect 19852 20244 19908 20254
rect 19852 20150 19908 20188
rect 19068 20018 19124 20076
rect 19068 19966 19070 20018
rect 19122 19966 19124 20018
rect 19068 19234 19124 19966
rect 20860 20018 20916 20030
rect 20860 19966 20862 20018
rect 20914 19966 20916 20018
rect 19068 19182 19070 19234
rect 19122 19182 19124 19234
rect 19068 19170 19124 19182
rect 19292 19908 19348 19918
rect 18732 19122 18788 19134
rect 18732 19070 18734 19122
rect 18786 19070 18788 19122
rect 18732 18788 18788 19070
rect 19180 19124 19236 19134
rect 18732 18732 18900 18788
rect 18732 18562 18788 18574
rect 18732 18510 18734 18562
rect 18786 18510 18788 18562
rect 18732 18228 18788 18510
rect 18844 18340 18900 18732
rect 18844 18274 18900 18284
rect 18956 18452 19012 18462
rect 18172 18172 18788 18228
rect 18172 17666 18228 18172
rect 18172 17614 18174 17666
rect 18226 17614 18228 17666
rect 18172 17602 18228 17614
rect 18284 17780 18340 17790
rect 18284 17666 18340 17724
rect 18620 17668 18676 17678
rect 18284 17614 18286 17666
rect 18338 17614 18340 17666
rect 18284 17602 18340 17614
rect 18508 17666 18676 17668
rect 18508 17614 18622 17666
rect 18674 17614 18676 17666
rect 18508 17612 18676 17614
rect 17724 17556 17780 17566
rect 17724 17554 18116 17556
rect 17724 17502 17726 17554
rect 17778 17502 18116 17554
rect 17724 17500 18116 17502
rect 17724 17490 17780 17500
rect 18060 17444 18116 17500
rect 18396 17554 18452 17566
rect 18396 17502 18398 17554
rect 18450 17502 18452 17554
rect 18396 17444 18452 17502
rect 18060 17388 18340 17444
rect 17500 17276 17780 17332
rect 17388 17042 17444 17052
rect 17612 17108 17668 17118
rect 16940 16940 17332 16996
rect 17276 16884 17332 16940
rect 17612 16994 17668 17052
rect 17612 16942 17614 16994
rect 17666 16942 17668 16994
rect 17388 16884 17444 16894
rect 16828 16828 17220 16884
rect 17276 16882 17556 16884
rect 17276 16830 17390 16882
rect 17442 16830 17556 16882
rect 17276 16828 17556 16830
rect 16492 15698 16548 15708
rect 16604 16098 16772 16100
rect 16604 16046 16718 16098
rect 16770 16046 16772 16098
rect 16604 16044 16772 16046
rect 16044 15538 16212 15540
rect 16044 15486 16046 15538
rect 16098 15486 16212 15538
rect 16044 15484 16212 15486
rect 16044 15316 16100 15484
rect 16044 15250 16100 15260
rect 16604 15148 16660 16044
rect 16716 16034 16772 16044
rect 17052 16436 17108 16446
rect 16940 15988 16996 15998
rect 16940 15894 16996 15932
rect 16492 15092 16660 15148
rect 16716 15764 16772 15774
rect 17052 15764 17108 16380
rect 16044 14306 16100 14318
rect 16044 14254 16046 14306
rect 16098 14254 16100 14306
rect 16044 14196 16100 14254
rect 16044 14130 16100 14140
rect 16380 14306 16436 14318
rect 16380 14254 16382 14306
rect 16434 14254 16436 14306
rect 16380 13972 16436 14254
rect 16380 13906 16436 13916
rect 16156 13748 16212 13758
rect 16156 13654 16212 13692
rect 15932 13346 15988 13356
rect 16156 13188 16212 13198
rect 16156 13094 16212 13132
rect 15596 13010 15652 13020
rect 16044 13076 16100 13086
rect 16044 12982 16100 13020
rect 15820 12964 15876 12974
rect 15820 12870 15876 12908
rect 16492 12964 16548 15092
rect 16716 14420 16772 15708
rect 16940 15708 17108 15764
rect 16828 15540 16884 15550
rect 16828 15446 16884 15484
rect 16604 14418 16772 14420
rect 16604 14366 16718 14418
rect 16770 14366 16772 14418
rect 16604 14364 16772 14366
rect 16604 13746 16660 14364
rect 16716 14354 16772 14364
rect 16940 14084 16996 15708
rect 16940 14018 16996 14028
rect 17052 14418 17108 14430
rect 17052 14366 17054 14418
rect 17106 14366 17108 14418
rect 17052 13972 17108 14366
rect 17164 14196 17220 16828
rect 17388 16818 17444 16828
rect 17276 16660 17332 16670
rect 17276 14644 17332 16604
rect 17388 16436 17444 16446
rect 17388 16210 17444 16380
rect 17388 16158 17390 16210
rect 17442 16158 17444 16210
rect 17388 16146 17444 16158
rect 17500 16212 17556 16828
rect 17612 16548 17668 16942
rect 17724 16660 17780 17276
rect 18172 17220 18228 17230
rect 17836 17164 18172 17220
rect 17836 16994 17892 17164
rect 17836 16942 17838 16994
rect 17890 16942 17892 16994
rect 17836 16930 17892 16942
rect 17724 16594 17780 16604
rect 17612 16482 17668 16492
rect 17724 16212 17780 16222
rect 18060 16212 18116 17164
rect 18172 17154 18228 17164
rect 18284 17108 18340 17388
rect 18396 17378 18452 17388
rect 18396 17108 18452 17118
rect 18284 17106 18452 17108
rect 18284 17054 18398 17106
rect 18450 17054 18452 17106
rect 18284 17052 18452 17054
rect 18396 17042 18452 17052
rect 18172 16884 18228 16894
rect 18508 16884 18564 17612
rect 18620 17602 18676 17612
rect 18956 16996 19012 18396
rect 18956 16930 19012 16940
rect 19068 17442 19124 17454
rect 19068 17390 19070 17442
rect 19122 17390 19124 17442
rect 19068 16994 19124 17390
rect 19068 16942 19070 16994
rect 19122 16942 19124 16994
rect 19068 16930 19124 16942
rect 18172 16882 18564 16884
rect 18172 16830 18174 16882
rect 18226 16830 18564 16882
rect 18172 16828 18564 16830
rect 18172 16818 18228 16828
rect 17500 16210 17780 16212
rect 17500 16158 17726 16210
rect 17778 16158 17780 16210
rect 17500 16156 17780 16158
rect 17500 15314 17556 16156
rect 17724 16146 17780 16156
rect 17836 16156 18116 16212
rect 17836 15988 17892 16156
rect 18060 16098 18116 16156
rect 18284 16100 18340 16828
rect 19180 16772 19236 19068
rect 19292 17556 19348 19852
rect 20524 19908 20580 19918
rect 20524 19814 20580 19852
rect 19516 19124 19572 19134
rect 19740 19124 19796 19134
rect 19516 19122 19796 19124
rect 19516 19070 19518 19122
rect 19570 19070 19742 19122
rect 19794 19070 19796 19122
rect 19516 19068 19796 19070
rect 19516 19058 19572 19068
rect 19740 19058 19796 19068
rect 20524 19124 20580 19134
rect 20076 19012 20132 19050
rect 20524 19030 20580 19068
rect 20076 18946 20132 18956
rect 20748 19012 20804 19022
rect 19860 18844 20124 18854
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 19860 18778 20124 18788
rect 20188 18676 20244 18686
rect 20188 18582 20244 18620
rect 19964 18564 20020 18574
rect 19404 18452 19460 18462
rect 19852 18452 19908 18462
rect 19404 17780 19460 18396
rect 19628 18450 19908 18452
rect 19628 18398 19854 18450
rect 19906 18398 19908 18450
rect 19628 18396 19908 18398
rect 19516 18340 19572 18350
rect 19516 18246 19572 18284
rect 19404 17686 19460 17724
rect 19292 17500 19572 17556
rect 19404 16996 19460 17006
rect 18060 16046 18062 16098
rect 18114 16046 18116 16098
rect 18060 16034 18116 16046
rect 18172 16098 18340 16100
rect 18172 16046 18286 16098
rect 18338 16046 18340 16098
rect 18172 16044 18340 16046
rect 17500 15262 17502 15314
rect 17554 15262 17556 15314
rect 17500 15148 17556 15262
rect 17276 14578 17332 14588
rect 17388 15092 17556 15148
rect 17612 15428 17668 15438
rect 17164 14130 17220 14140
rect 17052 13906 17108 13916
rect 17276 14084 17332 14094
rect 16828 13860 16884 13870
rect 16828 13858 16996 13860
rect 16828 13806 16830 13858
rect 16882 13806 16996 13858
rect 16828 13804 16996 13806
rect 16828 13794 16884 13804
rect 16604 13694 16606 13746
rect 16658 13694 16660 13746
rect 16604 13682 16660 13694
rect 16492 12898 16548 12908
rect 15484 12126 15486 12178
rect 15538 12126 15540 12178
rect 15484 12114 15540 12126
rect 15708 12850 15764 12862
rect 15708 12798 15710 12850
rect 15762 12798 15764 12850
rect 15260 12068 15316 12078
rect 15260 11974 15316 12012
rect 15036 11954 15204 11956
rect 15036 11902 15038 11954
rect 15090 11902 15204 11954
rect 15036 11900 15204 11902
rect 15708 11956 15764 12798
rect 16268 12852 16324 12862
rect 16268 12402 16324 12796
rect 16828 12852 16884 12862
rect 16828 12758 16884 12796
rect 16268 12350 16270 12402
rect 16322 12350 16324 12402
rect 16268 12338 16324 12350
rect 15820 12068 15876 12078
rect 15820 11974 15876 12012
rect 15932 12068 15988 12078
rect 16380 12068 16436 12078
rect 15932 12066 16212 12068
rect 15932 12014 15934 12066
rect 15986 12014 16212 12066
rect 15932 12012 16212 12014
rect 15932 12002 15988 12012
rect 15036 11890 15092 11900
rect 15708 11890 15764 11900
rect 15198 11788 15462 11798
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15198 11722 15462 11732
rect 14924 11442 14980 11452
rect 16044 11508 16100 11518
rect 16044 11394 16100 11452
rect 16044 11342 16046 11394
rect 16098 11342 16100 11394
rect 16044 11330 16100 11342
rect 16156 11282 16212 12012
rect 16156 11230 16158 11282
rect 16210 11230 16212 11282
rect 15036 11172 15092 11182
rect 15036 11078 15092 11116
rect 15484 11172 15540 11182
rect 15484 10836 15540 11116
rect 15484 10770 15540 10780
rect 16156 10836 16212 11230
rect 16156 10770 16212 10780
rect 16268 12066 16436 12068
rect 16268 12014 16382 12066
rect 16434 12014 16436 12066
rect 16268 12012 16436 12014
rect 16268 11060 16324 12012
rect 16380 12002 16436 12012
rect 16716 11396 16772 11406
rect 16940 11396 16996 13804
rect 17052 12964 17108 12974
rect 17052 12740 17108 12908
rect 17052 12674 17108 12684
rect 16772 11340 16996 11396
rect 17276 11508 17332 14028
rect 17388 13076 17444 15092
rect 17500 14308 17556 14318
rect 17612 14308 17668 15372
rect 17836 15426 17892 15932
rect 17948 15986 18004 15998
rect 17948 15934 17950 15986
rect 18002 15934 18004 15986
rect 17948 15540 18004 15934
rect 17948 15474 18004 15484
rect 18172 15876 18228 16044
rect 18284 16034 18340 16044
rect 18620 16716 19236 16772
rect 19292 16994 19460 16996
rect 19292 16942 19406 16994
rect 19458 16942 19460 16994
rect 19292 16940 19460 16942
rect 18620 16212 18676 16716
rect 18620 15876 18676 16156
rect 18732 16100 18788 16110
rect 19180 16100 19236 16110
rect 18732 16098 19236 16100
rect 18732 16046 18734 16098
rect 18786 16046 19182 16098
rect 19234 16046 19236 16098
rect 18732 16044 19236 16046
rect 18732 16034 18788 16044
rect 19180 16034 19236 16044
rect 18620 15820 18788 15876
rect 17836 15374 17838 15426
rect 17890 15374 17892 15426
rect 17836 15362 17892 15374
rect 18172 15314 18228 15820
rect 18620 15426 18676 15438
rect 18620 15374 18622 15426
rect 18674 15374 18676 15426
rect 18172 15262 18174 15314
rect 18226 15262 18228 15314
rect 18172 15250 18228 15262
rect 18396 15316 18452 15326
rect 18396 15222 18452 15260
rect 17836 14644 17892 14654
rect 17724 14420 17780 14430
rect 17724 14326 17780 14364
rect 17556 14252 17668 14308
rect 17500 14214 17556 14252
rect 17500 14084 17556 14094
rect 17556 14028 17668 14084
rect 17500 14018 17556 14028
rect 17612 13746 17668 14028
rect 17612 13694 17614 13746
rect 17666 13694 17668 13746
rect 17612 13682 17668 13694
rect 17724 13860 17780 13870
rect 17836 13860 17892 14588
rect 17948 14532 18004 14542
rect 17948 14418 18004 14476
rect 18508 14532 18564 14542
rect 18508 14438 18564 14476
rect 17948 14366 17950 14418
rect 18002 14366 18004 14418
rect 17948 14354 18004 14366
rect 18060 14420 18116 14430
rect 18060 14326 18116 14364
rect 18620 13860 18676 15374
rect 18732 14418 18788 15820
rect 18956 15874 19012 15886
rect 18956 15822 18958 15874
rect 19010 15822 19012 15874
rect 18844 15316 18900 15326
rect 18844 15222 18900 15260
rect 18956 15204 19012 15822
rect 19292 15540 19348 16940
rect 19404 16930 19460 16940
rect 19516 16324 19572 17500
rect 18956 15138 19012 15148
rect 19068 15484 19348 15540
rect 19404 15540 19460 15550
rect 19516 15540 19572 16268
rect 19628 16100 19684 18396
rect 19852 18386 19908 18396
rect 19740 17556 19796 17566
rect 19964 17556 20020 18508
rect 19740 17554 20020 17556
rect 19740 17502 19742 17554
rect 19794 17502 20020 17554
rect 19740 17500 20020 17502
rect 20076 17556 20132 17566
rect 20076 17554 20244 17556
rect 20076 17502 20078 17554
rect 20130 17502 20244 17554
rect 20076 17500 20244 17502
rect 19740 17490 19796 17500
rect 20076 17490 20132 17500
rect 19860 17276 20124 17286
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 19860 17210 20124 17220
rect 19964 16996 20020 17006
rect 19964 16902 20020 16940
rect 20188 16882 20244 17500
rect 20188 16830 20190 16882
rect 20242 16830 20244 16882
rect 19740 16100 19796 16110
rect 19628 16098 19796 16100
rect 19628 16046 19742 16098
rect 19794 16046 19796 16098
rect 19628 16044 19796 16046
rect 19404 15538 19572 15540
rect 19404 15486 19406 15538
rect 19458 15486 19572 15538
rect 19404 15484 19572 15486
rect 18732 14366 18734 14418
rect 18786 14366 18788 14418
rect 18732 14354 18788 14366
rect 18844 14756 18900 14766
rect 18844 13970 18900 14700
rect 19068 14084 19124 15484
rect 19404 15474 19460 15484
rect 19180 15316 19236 15326
rect 19180 14530 19236 15260
rect 19180 14478 19182 14530
rect 19234 14478 19236 14530
rect 19180 14308 19236 14478
rect 19628 15314 19684 15326
rect 19628 15262 19630 15314
rect 19682 15262 19684 15314
rect 19628 14530 19684 15262
rect 19628 14478 19630 14530
rect 19682 14478 19684 14530
rect 19628 14420 19684 14478
rect 19628 14354 19684 14364
rect 19180 14242 19236 14252
rect 19628 14196 19684 14206
rect 19068 14028 19348 14084
rect 18844 13918 18846 13970
rect 18898 13918 18900 13970
rect 18844 13906 18900 13918
rect 17724 13858 17892 13860
rect 17724 13806 17726 13858
rect 17778 13806 17892 13858
rect 17724 13804 17892 13806
rect 18508 13804 18676 13860
rect 17724 13748 17780 13804
rect 17724 13682 17780 13692
rect 17948 13746 18004 13758
rect 18172 13748 18228 13758
rect 17948 13694 17950 13746
rect 18002 13694 18004 13746
rect 17500 13636 17556 13646
rect 17500 13300 17556 13580
rect 17500 13244 17780 13300
rect 17500 13076 17556 13086
rect 17388 13074 17556 13076
rect 17388 13022 17502 13074
rect 17554 13022 17556 13074
rect 17388 13020 17556 13022
rect 17500 13010 17556 13020
rect 17724 12964 17780 13244
rect 17500 12852 17556 12862
rect 17556 12796 17668 12852
rect 17500 12786 17556 12796
rect 17500 12404 17556 12414
rect 17500 12310 17556 12348
rect 17276 11394 17332 11452
rect 17276 11342 17278 11394
rect 17330 11342 17332 11394
rect 16716 11302 16772 11340
rect 17276 11330 17332 11342
rect 16380 11284 16436 11294
rect 16380 11190 16436 11228
rect 17388 11282 17444 11294
rect 17388 11230 17390 11282
rect 17442 11230 17444 11282
rect 16940 11172 16996 11182
rect 16940 11078 16996 11116
rect 16268 10612 16324 11004
rect 17276 11060 17332 11070
rect 17388 11060 17444 11230
rect 17612 11284 17668 12796
rect 17724 12404 17780 12908
rect 17948 12852 18004 13694
rect 17948 12758 18004 12796
rect 18060 13746 18228 13748
rect 18060 13694 18174 13746
rect 18226 13694 18228 13746
rect 18060 13692 18228 13694
rect 18060 12962 18116 13692
rect 18172 13682 18228 13692
rect 18508 13188 18564 13804
rect 19068 13746 19124 13758
rect 19068 13694 19070 13746
rect 19122 13694 19124 13746
rect 18620 13636 18676 13646
rect 19068 13636 19124 13694
rect 18620 13634 19124 13636
rect 18620 13582 18622 13634
rect 18674 13582 19124 13634
rect 18620 13580 19124 13582
rect 18620 13570 18676 13580
rect 18060 12910 18062 12962
rect 18114 12910 18116 12962
rect 17724 12338 17780 12348
rect 17724 11396 17780 11406
rect 18060 11396 18116 12910
rect 18396 13132 18564 13188
rect 18396 12740 18452 13132
rect 18508 12964 18564 12974
rect 19068 12964 19124 12974
rect 18508 12962 19124 12964
rect 18508 12910 18510 12962
rect 18562 12910 19070 12962
rect 19122 12910 19124 12962
rect 18508 12908 19124 12910
rect 18508 12898 18564 12908
rect 19068 12898 19124 12908
rect 18396 12684 18564 12740
rect 17780 11340 18116 11396
rect 17724 11302 17780 11340
rect 17612 11190 17668 11228
rect 18396 11284 18452 11294
rect 18396 11190 18452 11228
rect 17332 11004 17444 11060
rect 18172 11170 18228 11182
rect 18172 11118 18174 11170
rect 18226 11118 18228 11170
rect 17276 10994 17332 11004
rect 16044 10556 16324 10612
rect 16716 10724 16772 10734
rect 18060 10724 18116 10734
rect 15198 10220 15462 10230
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15198 10154 15462 10164
rect 15198 8652 15462 8662
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15198 8586 15462 8596
rect 15198 7084 15462 7094
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15198 7018 15462 7028
rect 15198 5516 15462 5526
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15198 5450 15462 5460
rect 15932 4228 15988 4238
rect 15596 4226 15988 4228
rect 15596 4174 15934 4226
rect 15986 4174 15988 4226
rect 15596 4172 15988 4174
rect 15198 3948 15462 3958
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15198 3882 15462 3892
rect 15596 3668 15652 4172
rect 15932 4162 15988 4172
rect 16044 4004 16100 10556
rect 16380 4452 16436 4462
rect 15484 3612 15652 3668
rect 15932 3948 16100 4004
rect 16156 4450 16436 4452
rect 16156 4398 16382 4450
rect 16434 4398 16436 4450
rect 16156 4396 16436 4398
rect 14924 3556 14980 3566
rect 14812 3554 14980 3556
rect 14812 3502 14926 3554
rect 14978 3502 14980 3554
rect 14812 3500 14980 3502
rect 14924 3490 14980 3500
rect 15484 3554 15540 3612
rect 15484 3502 15486 3554
rect 15538 3502 15540 3554
rect 14028 3332 14084 3342
rect 14364 3332 14644 3388
rect 14700 3332 14756 3342
rect 14028 3330 14196 3332
rect 14028 3278 14030 3330
rect 14082 3278 14196 3330
rect 14028 3276 14196 3278
rect 14028 3266 14084 3276
rect 14140 800 14196 3276
rect 14700 3330 14868 3332
rect 14700 3278 14702 3330
rect 14754 3278 14868 3330
rect 14700 3276 14868 3278
rect 14700 3266 14756 3276
rect 14812 800 14868 3276
rect 15484 800 15540 3502
rect 15708 3444 15764 3454
rect 15932 3444 15988 3948
rect 16044 3556 16100 3566
rect 16044 3462 16100 3500
rect 15708 3442 15988 3444
rect 15708 3390 15710 3442
rect 15762 3390 15988 3442
rect 15708 3388 15988 3390
rect 15708 3378 15764 3388
rect 16156 800 16212 4396
rect 16380 4386 16436 4396
rect 16716 4450 16772 10668
rect 16716 4398 16718 4450
rect 16770 4398 16772 4450
rect 16716 4386 16772 4398
rect 17276 10722 18116 10724
rect 17276 10670 18062 10722
rect 18114 10670 18116 10722
rect 17276 10668 18116 10670
rect 17276 3554 17332 10668
rect 18060 10658 18116 10668
rect 18172 10612 18228 11118
rect 18284 10612 18340 10622
rect 18172 10610 18340 10612
rect 18172 10558 18286 10610
rect 18338 10558 18340 10610
rect 18172 10556 18340 10558
rect 18284 10546 18340 10556
rect 18508 5012 18564 12684
rect 18844 12738 18900 12750
rect 18844 12686 18846 12738
rect 18898 12686 18900 12738
rect 18732 11172 18788 11182
rect 18620 11170 18788 11172
rect 18620 11118 18734 11170
rect 18786 11118 18788 11170
rect 18620 11116 18788 11118
rect 18620 9156 18676 11116
rect 18732 11106 18788 11116
rect 18732 10724 18788 10734
rect 18732 10630 18788 10668
rect 18732 9156 18788 9166
rect 18620 9100 18732 9156
rect 18732 9090 18788 9100
rect 18844 8036 18900 12686
rect 19068 11282 19124 11294
rect 19068 11230 19070 11282
rect 19122 11230 19124 11282
rect 18956 11172 19012 11182
rect 18956 10610 19012 11116
rect 19068 11060 19124 11230
rect 19068 10994 19124 11004
rect 18956 10558 18958 10610
rect 19010 10558 19012 10610
rect 18956 10546 19012 10558
rect 17276 3502 17278 3554
rect 17330 3502 17332 3554
rect 17276 3490 17332 3502
rect 17948 4956 18564 5012
rect 18732 7980 18900 8036
rect 18956 10164 19012 10174
rect 18956 9042 19012 10108
rect 18956 8990 18958 9042
rect 19010 8990 19012 9042
rect 17948 3554 18004 4956
rect 17948 3502 17950 3554
rect 18002 3502 18004 3554
rect 17948 3490 18004 3502
rect 18508 3554 18564 3566
rect 18508 3502 18510 3554
rect 18562 3502 18564 3554
rect 16380 3442 16436 3454
rect 16380 3390 16382 3442
rect 16434 3390 16436 3442
rect 16380 3388 16436 3390
rect 16380 3332 16884 3388
rect 16828 800 16884 3332
rect 17500 3330 17556 3342
rect 17500 3278 17502 3330
rect 17554 3278 17556 3330
rect 17500 800 17556 3278
rect 18172 3330 18228 3342
rect 18172 3278 18174 3330
rect 18226 3278 18228 3330
rect 18172 800 18228 3278
rect 18508 3332 18564 3502
rect 18732 3332 18788 7980
rect 18956 7476 19012 8990
rect 18956 7382 19012 7420
rect 19292 3554 19348 14028
rect 19516 13972 19572 13982
rect 19516 13878 19572 13916
rect 19628 13858 19684 14140
rect 19628 13806 19630 13858
rect 19682 13806 19684 13858
rect 19628 13748 19684 13806
rect 19516 13692 19684 13748
rect 19404 11620 19460 11630
rect 19404 11282 19460 11564
rect 19404 11230 19406 11282
rect 19458 11230 19460 11282
rect 19404 11218 19460 11230
rect 19404 10836 19460 10846
rect 19404 9938 19460 10780
rect 19404 9886 19406 9938
rect 19458 9886 19460 9938
rect 19404 9874 19460 9886
rect 19516 9156 19572 13692
rect 19740 12964 19796 16044
rect 20076 15876 20132 15886
rect 20188 15876 20244 16830
rect 20636 16994 20692 17006
rect 20636 16942 20638 16994
rect 20690 16942 20692 16994
rect 20636 16772 20692 16942
rect 20636 16100 20692 16716
rect 20636 16034 20692 16044
rect 20076 15874 20244 15876
rect 20076 15822 20078 15874
rect 20130 15822 20244 15874
rect 20076 15820 20244 15822
rect 20076 15810 20132 15820
rect 19860 15708 20124 15718
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 19860 15642 20124 15652
rect 20188 15204 20244 15820
rect 20188 15138 20244 15148
rect 20524 15652 20580 15662
rect 20524 15148 20580 15596
rect 20748 15148 20804 18956
rect 20860 18676 20916 19966
rect 20972 19012 21028 20636
rect 21084 19684 21140 21980
rect 21308 21700 21364 21710
rect 21308 21606 21364 21644
rect 21644 21588 21700 22316
rect 21868 22258 21924 22540
rect 22428 22372 22484 22382
rect 22428 22278 22484 22316
rect 22652 22370 22708 22540
rect 22876 22372 22932 24332
rect 22652 22318 22654 22370
rect 22706 22318 22708 22370
rect 22652 22306 22708 22318
rect 22764 22370 22932 22372
rect 22764 22318 22878 22370
rect 22930 22318 22932 22370
rect 22764 22316 22932 22318
rect 21868 22206 21870 22258
rect 21922 22206 21924 22258
rect 21868 22194 21924 22206
rect 22540 22260 22596 22270
rect 22540 22166 22596 22204
rect 22764 22036 22820 22316
rect 22876 22306 22932 22316
rect 22988 23828 23044 23838
rect 21980 21980 22820 22036
rect 21980 21810 22036 21980
rect 21980 21758 21982 21810
rect 22034 21758 22036 21810
rect 21980 21746 22036 21758
rect 21644 21522 21700 21532
rect 21756 21586 21812 21598
rect 21756 21534 21758 21586
rect 21810 21534 21812 21586
rect 21756 20916 21812 21534
rect 22876 21588 22932 21598
rect 22428 21474 22484 21486
rect 22428 21422 22430 21474
rect 22482 21422 22484 21474
rect 22428 20916 22484 21422
rect 21756 20860 22484 20916
rect 22876 21474 22932 21532
rect 22876 21422 22878 21474
rect 22930 21422 22932 21474
rect 21308 20692 21364 20702
rect 21980 20692 22036 20702
rect 21308 20244 21364 20636
rect 21868 20690 22036 20692
rect 21868 20638 21982 20690
rect 22034 20638 22036 20690
rect 21868 20636 22036 20638
rect 21644 20580 21700 20590
rect 21644 20486 21700 20524
rect 21308 20178 21364 20188
rect 21196 20132 21252 20142
rect 21196 20038 21252 20076
rect 21644 20132 21700 20142
rect 21868 20132 21924 20636
rect 21980 20626 22036 20636
rect 21644 20130 21924 20132
rect 21644 20078 21646 20130
rect 21698 20078 21924 20130
rect 21644 20076 21924 20078
rect 21644 20020 21700 20076
rect 21644 19954 21700 19964
rect 21980 20020 22036 20030
rect 22092 20020 22148 20860
rect 22764 20692 22820 20702
rect 22764 20598 22820 20636
rect 22316 20580 22372 20590
rect 22316 20578 22484 20580
rect 22316 20526 22318 20578
rect 22370 20526 22484 20578
rect 22316 20524 22484 20526
rect 22316 20514 22372 20524
rect 21980 20018 22148 20020
rect 21980 19966 21982 20018
rect 22034 19966 22148 20018
rect 21980 19964 22148 19966
rect 22316 20130 22372 20142
rect 22316 20078 22318 20130
rect 22370 20078 22372 20130
rect 22316 20020 22372 20078
rect 21980 19908 22036 19964
rect 22316 19954 22372 19964
rect 21980 19842 22036 19852
rect 22428 19796 22484 20524
rect 22876 20468 22932 21422
rect 22764 20412 22932 20468
rect 22764 20018 22820 20412
rect 22988 20356 23044 23772
rect 23100 23716 23156 24556
rect 23212 24052 23268 25452
rect 23436 25396 23492 25406
rect 23772 25396 23828 25406
rect 23436 25394 23828 25396
rect 23436 25342 23438 25394
rect 23490 25342 23774 25394
rect 23826 25342 23828 25394
rect 23436 25340 23828 25342
rect 23436 25330 23492 25340
rect 23772 25330 23828 25340
rect 23324 24052 23380 24062
rect 23212 23996 23324 24052
rect 23324 23826 23380 23996
rect 23324 23774 23326 23826
rect 23378 23774 23380 23826
rect 23324 23762 23380 23774
rect 23548 23938 23604 23950
rect 23548 23886 23550 23938
rect 23602 23886 23604 23938
rect 23100 23650 23156 23660
rect 23212 23604 23268 23614
rect 23212 22596 23268 23548
rect 23548 23604 23604 23886
rect 23548 23538 23604 23548
rect 23772 23268 23828 23278
rect 23772 23174 23828 23212
rect 23436 23156 23492 23166
rect 22764 19966 22766 20018
rect 22818 19966 22820 20018
rect 22540 19796 22596 19806
rect 22428 19740 22540 19796
rect 22540 19730 22596 19740
rect 21084 19628 21700 19684
rect 21532 19234 21588 19246
rect 21532 19182 21534 19234
rect 21586 19182 21588 19234
rect 21308 19012 21364 19022
rect 20972 19010 21476 19012
rect 20972 18958 21310 19010
rect 21362 18958 21476 19010
rect 20972 18956 21476 18958
rect 21308 18946 21364 18956
rect 20860 18610 20916 18620
rect 21420 18450 21476 18956
rect 21420 18398 21422 18450
rect 21474 18398 21476 18450
rect 21420 18386 21476 18398
rect 21084 18340 21140 18350
rect 21084 18246 21140 18284
rect 21532 16996 21588 19182
rect 21644 18562 21700 19628
rect 22652 19460 22708 19470
rect 22428 19234 22484 19246
rect 22428 19182 22430 19234
rect 22482 19182 22484 19234
rect 22428 18674 22484 19182
rect 22652 19122 22708 19404
rect 22652 19070 22654 19122
rect 22706 19070 22708 19122
rect 22652 19058 22708 19070
rect 22428 18622 22430 18674
rect 22482 18622 22484 18674
rect 22428 18610 22484 18622
rect 21644 18510 21646 18562
rect 21698 18510 21700 18562
rect 21644 18498 21700 18510
rect 22652 18562 22708 18574
rect 22652 18510 22654 18562
rect 22706 18510 22708 18562
rect 21756 18452 21812 18462
rect 22204 18452 22260 18462
rect 22652 18452 22708 18510
rect 21756 18450 21924 18452
rect 21756 18398 21758 18450
rect 21810 18398 21924 18450
rect 21756 18396 21924 18398
rect 21756 18386 21812 18396
rect 21756 17668 21812 17678
rect 21644 17612 21756 17668
rect 21644 17106 21700 17612
rect 21756 17574 21812 17612
rect 21868 17444 21924 18396
rect 22204 18450 22708 18452
rect 22204 18398 22206 18450
rect 22258 18398 22708 18450
rect 22204 18396 22708 18398
rect 22092 17444 22148 17454
rect 21868 17442 22148 17444
rect 21868 17390 22094 17442
rect 22146 17390 22148 17442
rect 21868 17388 22148 17390
rect 21644 17054 21646 17106
rect 21698 17054 21700 17106
rect 21644 17042 21700 17054
rect 21532 16930 21588 16940
rect 21980 16996 22036 17006
rect 21980 16902 22036 16940
rect 20972 16884 21028 16894
rect 21420 16884 21476 16894
rect 21868 16884 21924 16894
rect 20972 16882 21476 16884
rect 20972 16830 20974 16882
rect 21026 16830 21422 16882
rect 21474 16830 21476 16882
rect 20972 16828 21476 16830
rect 20972 16818 21028 16828
rect 21308 15986 21364 15998
rect 21308 15934 21310 15986
rect 21362 15934 21364 15986
rect 20972 15314 21028 15326
rect 20972 15262 20974 15314
rect 21026 15262 21028 15314
rect 20972 15204 21028 15262
rect 20524 15092 20692 15148
rect 20748 15092 20916 15148
rect 20972 15138 21028 15148
rect 21084 15314 21140 15326
rect 21084 15262 21086 15314
rect 21138 15262 21140 15314
rect 20636 14754 20692 15092
rect 20636 14702 20638 14754
rect 20690 14702 20692 14754
rect 20636 14690 20692 14702
rect 20188 14532 20244 14542
rect 19860 14140 20124 14150
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 19860 14074 20124 14084
rect 20076 13748 20132 13758
rect 20188 13748 20244 14476
rect 20524 14530 20580 14542
rect 20524 14478 20526 14530
rect 20578 14478 20580 14530
rect 20524 14420 20580 14478
rect 20524 13858 20580 14364
rect 20524 13806 20526 13858
rect 20578 13806 20580 13858
rect 20524 13794 20580 13806
rect 20076 13746 20244 13748
rect 20076 13694 20078 13746
rect 20130 13694 20244 13746
rect 20076 13692 20244 13694
rect 20076 13682 20132 13692
rect 19516 9090 19572 9100
rect 19628 12908 19796 12964
rect 20412 12964 20468 12974
rect 19628 7588 19684 12908
rect 20412 12870 20468 12908
rect 20748 12964 20804 12974
rect 20748 12850 20804 12908
rect 20748 12798 20750 12850
rect 20802 12798 20804 12850
rect 20748 12786 20804 12798
rect 19740 12740 19796 12750
rect 19740 12646 19796 12684
rect 20076 12740 20132 12750
rect 20188 12740 20244 12750
rect 20076 12738 20188 12740
rect 20076 12686 20078 12738
rect 20130 12686 20188 12738
rect 20076 12684 20188 12686
rect 20076 12674 20132 12684
rect 19860 12572 20124 12582
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 19860 12506 20124 12516
rect 20076 12180 20132 12190
rect 19740 11282 19796 11294
rect 19740 11230 19742 11282
rect 19794 11230 19796 11282
rect 19740 10836 19796 11230
rect 20076 11282 20132 12124
rect 20188 11396 20244 12684
rect 20412 11396 20468 11406
rect 20188 11340 20412 11396
rect 20076 11230 20078 11282
rect 20130 11230 20132 11282
rect 20076 11218 20132 11230
rect 20412 11282 20468 11340
rect 20412 11230 20414 11282
rect 20466 11230 20468 11282
rect 20412 11218 20468 11230
rect 20748 11282 20804 11294
rect 20748 11230 20750 11282
rect 20802 11230 20804 11282
rect 19860 11004 20124 11014
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 19860 10938 20124 10948
rect 19740 10770 19796 10780
rect 20636 10724 20692 10734
rect 20524 9716 20580 9726
rect 20524 9622 20580 9660
rect 20636 9714 20692 10668
rect 20748 10276 20804 11230
rect 20748 10210 20804 10220
rect 20860 9828 20916 15092
rect 21084 14980 21140 15262
rect 21196 15316 21252 15354
rect 21196 15250 21252 15260
rect 21308 15148 21364 15934
rect 21420 15876 21476 16828
rect 21756 16828 21868 16884
rect 21644 15988 21700 15998
rect 21756 15988 21812 16828
rect 21868 16818 21924 16828
rect 22092 16212 22148 17388
rect 21980 16156 22148 16212
rect 21980 16100 22036 16156
rect 21644 15986 21812 15988
rect 21644 15934 21646 15986
rect 21698 15934 21812 15986
rect 21644 15932 21812 15934
rect 21868 16044 22036 16100
rect 21644 15922 21700 15932
rect 21420 15810 21476 15820
rect 20972 14924 21140 14980
rect 21196 15092 21364 15148
rect 21644 15316 21700 15326
rect 21644 15202 21700 15260
rect 21644 15150 21646 15202
rect 21698 15150 21700 15202
rect 21644 15138 21700 15150
rect 21756 15204 21812 15214
rect 20972 14308 21028 14924
rect 20972 12740 21028 14252
rect 20972 12674 21028 12684
rect 21196 12292 21252 15092
rect 21308 14532 21364 14542
rect 21308 14438 21364 14476
rect 21756 13746 21812 15148
rect 21868 15148 21924 16044
rect 22092 15986 22148 15998
rect 22092 15934 22094 15986
rect 22146 15934 22148 15986
rect 21980 15876 22036 15886
rect 21980 15782 22036 15820
rect 21868 15092 22036 15148
rect 21980 14420 22036 15092
rect 21980 14354 22036 14364
rect 21868 14308 21924 14318
rect 21868 14214 21924 14252
rect 21756 13694 21758 13746
rect 21810 13694 21812 13746
rect 21756 13682 21812 13694
rect 22092 13636 22148 15934
rect 22204 14532 22260 18396
rect 22764 18340 22820 19966
rect 22652 18284 22820 18340
rect 22876 20300 23044 20356
rect 23100 22540 23268 22596
rect 23324 23154 23492 23156
rect 23324 23102 23438 23154
rect 23490 23102 23492 23154
rect 23324 23100 23492 23102
rect 23324 22594 23380 23100
rect 23436 23090 23492 23100
rect 23324 22542 23326 22594
rect 23378 22542 23380 22594
rect 22876 18450 22932 20300
rect 22988 20132 23044 20142
rect 22988 20038 23044 20076
rect 23100 19348 23156 22540
rect 23324 22530 23380 22542
rect 23212 22372 23268 22382
rect 23212 21586 23268 22316
rect 23548 22372 23604 22382
rect 23548 22258 23604 22316
rect 23548 22206 23550 22258
rect 23602 22206 23604 22258
rect 23548 22194 23604 22206
rect 23884 22370 23940 26236
rect 24108 25732 24164 26350
rect 24108 25666 24164 25676
rect 24220 26516 24276 26526
rect 24108 25396 24164 25406
rect 24220 25396 24276 26460
rect 24108 25394 24276 25396
rect 24108 25342 24110 25394
rect 24162 25342 24276 25394
rect 24108 25340 24276 25342
rect 24332 25732 24388 28476
rect 24780 28466 24836 28476
rect 24892 28642 25060 28644
rect 24892 28590 25006 28642
rect 25058 28590 25060 28642
rect 24892 28588 25060 28590
rect 25116 28644 25172 29036
rect 25228 28868 25284 28878
rect 25340 28868 25396 29148
rect 25452 29110 25508 29148
rect 25228 28866 25396 28868
rect 25228 28814 25230 28866
rect 25282 28814 25396 28866
rect 25228 28812 25396 28814
rect 25564 28866 25620 29260
rect 25564 28814 25566 28866
rect 25618 28814 25620 28866
rect 25228 28802 25284 28812
rect 25564 28802 25620 28814
rect 25116 28588 25508 28644
rect 24522 27468 24786 27478
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24522 27402 24786 27412
rect 24668 27076 24724 27086
rect 24668 26982 24724 27020
rect 24892 27074 24948 28588
rect 25004 28578 25060 28588
rect 25452 27972 25508 28588
rect 26012 28642 26068 28654
rect 26012 28590 26014 28642
rect 26066 28590 26068 28642
rect 25452 27878 25508 27916
rect 25900 28532 25956 28542
rect 25340 27860 25396 27870
rect 25340 27766 25396 27804
rect 25564 27858 25620 27870
rect 25564 27806 25566 27858
rect 25618 27806 25620 27858
rect 25564 27412 25620 27806
rect 25340 27356 25620 27412
rect 24892 27022 24894 27074
rect 24946 27022 24948 27074
rect 24892 26404 24948 27022
rect 25004 27076 25060 27086
rect 25340 27076 25396 27356
rect 25004 27074 25340 27076
rect 25004 27022 25006 27074
rect 25058 27022 25340 27074
rect 25004 27020 25340 27022
rect 25004 27010 25060 27020
rect 25340 26982 25396 27020
rect 25452 26964 25508 26974
rect 25788 26964 25844 26974
rect 25452 26962 25844 26964
rect 25452 26910 25454 26962
rect 25506 26910 25790 26962
rect 25842 26910 25844 26962
rect 25452 26908 25844 26910
rect 25452 26898 25508 26908
rect 25788 26898 25844 26908
rect 24892 26338 24948 26348
rect 24522 25900 24786 25910
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24522 25834 24786 25844
rect 24668 25732 24724 25742
rect 24332 25730 24724 25732
rect 24332 25678 24670 25730
rect 24722 25678 24724 25730
rect 24332 25676 24724 25678
rect 24108 25330 24164 25340
rect 24332 24500 24388 25676
rect 24668 25666 24724 25676
rect 24444 25508 24500 25518
rect 24444 25414 24500 25452
rect 25004 25396 25060 25406
rect 25340 25396 25396 25406
rect 25004 25394 25396 25396
rect 25004 25342 25006 25394
rect 25058 25342 25342 25394
rect 25394 25342 25396 25394
rect 25004 25340 25396 25342
rect 25004 25330 25060 25340
rect 25340 25330 25396 25340
rect 25676 25396 25732 25406
rect 25900 25396 25956 28476
rect 26012 28082 26068 28590
rect 26012 28030 26014 28082
rect 26066 28030 26068 28082
rect 26012 28018 26068 28030
rect 26124 26962 26180 29708
rect 26236 28530 26292 33852
rect 26460 33684 26516 33694
rect 26236 28478 26238 28530
rect 26290 28478 26292 28530
rect 26236 28466 26292 28478
rect 26348 32564 26404 32574
rect 26124 26910 26126 26962
rect 26178 26910 26180 26962
rect 26124 26898 26180 26910
rect 26348 26908 26404 32508
rect 26460 30098 26516 33628
rect 26460 30046 26462 30098
rect 26514 30046 26516 30098
rect 26460 30034 26516 30046
rect 26796 29764 26852 36204
rect 27132 35922 27188 37436
rect 28140 37156 28196 37772
rect 28252 37268 28308 39200
rect 28924 37828 28980 39200
rect 29596 37828 29652 39200
rect 30268 37828 30324 39200
rect 30940 37828 30996 39200
rect 28924 37772 29540 37828
rect 29596 37772 29876 37828
rect 30268 37772 30884 37828
rect 30940 37772 31220 37828
rect 29484 37716 29540 37772
rect 29484 37660 29764 37716
rect 28252 37212 28532 37268
rect 28140 37100 28420 37156
rect 27244 36932 27300 36942
rect 27244 36370 27300 36876
rect 27468 36484 27524 36494
rect 27468 36390 27524 36428
rect 27244 36318 27246 36370
rect 27298 36318 27300 36370
rect 27244 36306 27300 36318
rect 27692 36372 27748 36382
rect 27132 35870 27134 35922
rect 27186 35870 27188 35922
rect 27132 35858 27188 35870
rect 27356 35698 27412 35710
rect 27356 35646 27358 35698
rect 27410 35646 27412 35698
rect 27356 33572 27412 35646
rect 27356 33506 27412 33516
rect 27580 35364 27636 35374
rect 26796 29698 26852 29708
rect 27244 30098 27300 30110
rect 27244 30046 27246 30098
rect 27298 30046 27300 30098
rect 27132 29652 27188 29662
rect 27244 29652 27300 30046
rect 27580 30098 27636 35308
rect 27580 30046 27582 30098
rect 27634 30046 27636 30098
rect 27580 30034 27636 30046
rect 27132 29650 27300 29652
rect 27132 29598 27134 29650
rect 27186 29598 27300 29650
rect 27132 29596 27300 29598
rect 27132 29586 27188 29596
rect 27692 29540 27748 36316
rect 28364 36370 28420 37100
rect 28364 36318 28366 36370
rect 28418 36318 28420 36370
rect 28364 36306 28420 36318
rect 28476 36260 28532 37212
rect 29260 36484 29316 36494
rect 28924 36482 29316 36484
rect 28924 36430 29262 36482
rect 29314 36430 29316 36482
rect 28924 36428 29316 36430
rect 28700 36372 28756 36382
rect 28700 36278 28756 36316
rect 28476 36194 28532 36204
rect 28252 33572 28308 33582
rect 28028 30210 28084 30222
rect 28028 30158 28030 30210
rect 28082 30158 28084 30210
rect 28028 29650 28084 30158
rect 28252 30098 28308 33516
rect 28812 30996 28868 31006
rect 28252 30046 28254 30098
rect 28306 30046 28308 30098
rect 28252 30034 28308 30046
rect 28700 30940 28812 30996
rect 28028 29598 28030 29650
rect 28082 29598 28084 29650
rect 28028 29586 28084 29598
rect 27244 29484 27748 29540
rect 26572 29316 26628 29326
rect 26572 27970 26628 29260
rect 26796 29204 26852 29214
rect 26796 29110 26852 29148
rect 26572 27918 26574 27970
rect 26626 27918 26628 27970
rect 26572 27906 26628 27918
rect 26460 27860 26516 27870
rect 26460 27766 26516 27804
rect 26684 27860 26740 27870
rect 25676 25394 25956 25396
rect 25676 25342 25678 25394
rect 25730 25342 25956 25394
rect 25676 25340 25956 25342
rect 26236 26852 26404 26908
rect 26460 27076 26516 27086
rect 26684 27076 26740 27804
rect 27132 27636 27188 27646
rect 26516 27020 26740 27076
rect 26908 27634 27188 27636
rect 26908 27582 27134 27634
rect 27186 27582 27188 27634
rect 26908 27580 27188 27582
rect 26908 27074 26964 27580
rect 27132 27570 27188 27580
rect 26908 27022 26910 27074
rect 26962 27022 26964 27074
rect 25676 25330 25732 25340
rect 24668 24836 24724 24846
rect 26236 24836 26292 26852
rect 26460 26514 26516 27020
rect 26908 27010 26964 27022
rect 27132 26964 27188 26974
rect 27244 26964 27300 29484
rect 27468 29316 27524 29326
rect 27524 29260 27636 29316
rect 27468 29222 27524 29260
rect 27356 29204 27412 29214
rect 27356 28530 27412 29148
rect 27356 28478 27358 28530
rect 27410 28478 27412 28530
rect 27356 28466 27412 28478
rect 27580 27972 27636 29260
rect 27692 29204 27748 29214
rect 27692 29110 27748 29148
rect 27692 28532 27748 28542
rect 27692 28530 27972 28532
rect 27692 28478 27694 28530
rect 27746 28478 27972 28530
rect 27692 28476 27972 28478
rect 27692 28466 27748 28476
rect 27692 27972 27748 27982
rect 27580 27970 27748 27972
rect 27580 27918 27694 27970
rect 27746 27918 27748 27970
rect 27580 27916 27748 27918
rect 27692 27906 27748 27916
rect 27132 26962 27300 26964
rect 27132 26910 27134 26962
rect 27186 26910 27300 26962
rect 27132 26908 27300 26910
rect 27468 27858 27524 27870
rect 27468 27806 27470 27858
rect 27522 27806 27524 27858
rect 27132 26898 27188 26908
rect 26460 26462 26462 26514
rect 26514 26462 26516 26514
rect 26460 26450 26516 26462
rect 26796 26292 26852 26302
rect 26796 26290 26964 26292
rect 26796 26238 26798 26290
rect 26850 26238 26964 26290
rect 26796 26236 26964 26238
rect 26796 26226 26852 26236
rect 26572 25508 26628 25518
rect 24668 24742 24724 24780
rect 25452 24780 26292 24836
rect 26460 25506 26628 25508
rect 26460 25454 26574 25506
rect 26626 25454 26628 25506
rect 26460 25452 26628 25454
rect 24444 24724 24500 24734
rect 24444 24630 24500 24668
rect 25228 24724 25284 24734
rect 25228 24630 25284 24668
rect 24332 24164 24388 24444
rect 25228 24388 25284 24398
rect 24522 24332 24786 24342
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24522 24266 24786 24276
rect 24444 24164 24500 24174
rect 24108 24162 24500 24164
rect 24108 24110 24446 24162
rect 24498 24110 24500 24162
rect 24108 24108 24500 24110
rect 24108 23378 24164 24108
rect 24444 24098 24500 24108
rect 24220 23940 24276 23950
rect 24220 23846 24276 23884
rect 24780 23828 24836 23838
rect 25116 23828 25172 23838
rect 24780 23826 25172 23828
rect 24780 23774 24782 23826
rect 24834 23774 25118 23826
rect 25170 23774 25172 23826
rect 24780 23772 25172 23774
rect 24780 23762 24836 23772
rect 25116 23762 25172 23772
rect 24108 23326 24110 23378
rect 24162 23326 24164 23378
rect 24108 23314 24164 23326
rect 25228 23380 25284 24332
rect 25452 23826 25508 24780
rect 26348 24724 26404 24734
rect 26460 24724 26516 25452
rect 26572 25442 26628 25452
rect 26796 25508 26852 25518
rect 26796 25414 26852 25452
rect 26908 25506 26964 26236
rect 26908 25454 26910 25506
rect 26962 25454 26964 25506
rect 26908 25172 26964 25454
rect 26684 25116 26964 25172
rect 27020 26068 27076 26078
rect 26684 24834 26740 25116
rect 26684 24782 26686 24834
rect 26738 24782 26740 24834
rect 26348 24722 26516 24724
rect 26348 24670 26350 24722
rect 26402 24670 26516 24722
rect 26348 24668 26516 24670
rect 26572 24722 26628 24734
rect 26572 24670 26574 24722
rect 26626 24670 26628 24722
rect 25788 24612 25844 24622
rect 25788 24518 25844 24556
rect 25564 24500 25620 24510
rect 25564 24406 25620 24444
rect 25452 23774 25454 23826
rect 25506 23774 25508 23826
rect 25452 23762 25508 23774
rect 25676 24276 25732 24286
rect 25228 23314 25284 23324
rect 24444 23156 24500 23166
rect 24444 23062 24500 23100
rect 24522 22764 24786 22774
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24522 22698 24786 22708
rect 23884 22318 23886 22370
rect 23938 22318 23940 22370
rect 23324 21700 23380 21710
rect 23324 21606 23380 21644
rect 23660 21698 23716 21710
rect 23660 21646 23662 21698
rect 23714 21646 23716 21698
rect 23212 21534 23214 21586
rect 23266 21534 23268 21586
rect 23212 20916 23268 21534
rect 23324 20916 23380 20926
rect 23212 20914 23380 20916
rect 23212 20862 23326 20914
rect 23378 20862 23380 20914
rect 23212 20860 23380 20862
rect 22876 18398 22878 18450
rect 22930 18398 22932 18450
rect 22316 16994 22372 17006
rect 22316 16942 22318 16994
rect 22370 16942 22372 16994
rect 22316 16324 22372 16942
rect 22652 16772 22708 18284
rect 22764 17668 22820 17678
rect 22764 17574 22820 17612
rect 22876 16994 22932 18398
rect 22988 19292 23156 19348
rect 23212 20244 23268 20254
rect 22988 17668 23044 19292
rect 23212 19234 23268 20188
rect 23324 20018 23380 20860
rect 23548 20690 23604 20702
rect 23548 20638 23550 20690
rect 23602 20638 23604 20690
rect 23548 20580 23604 20638
rect 23660 20692 23716 21646
rect 23772 20692 23828 20702
rect 23660 20690 23828 20692
rect 23660 20638 23774 20690
rect 23826 20638 23828 20690
rect 23660 20636 23828 20638
rect 23548 20514 23604 20524
rect 23772 20132 23828 20636
rect 23884 20244 23940 22318
rect 24668 22484 24724 22494
rect 24332 22258 24388 22270
rect 24332 22206 24334 22258
rect 24386 22206 24388 22258
rect 24220 21812 24276 21822
rect 24332 21812 24388 22206
rect 24668 22258 24724 22428
rect 24668 22206 24670 22258
rect 24722 22206 24724 22258
rect 24668 22194 24724 22206
rect 25676 22370 25732 24220
rect 26348 23940 26404 24668
rect 26572 24612 26628 24670
rect 26572 24546 26628 24556
rect 26236 23938 26404 23940
rect 26236 23886 26350 23938
rect 26402 23886 26404 23938
rect 26236 23884 26404 23886
rect 26124 23154 26180 23166
rect 26124 23102 26126 23154
rect 26178 23102 26180 23154
rect 25676 22318 25678 22370
rect 25730 22318 25732 22370
rect 24220 21810 24388 21812
rect 24220 21758 24222 21810
rect 24274 21758 24388 21810
rect 24220 21756 24388 21758
rect 25676 21812 25732 22318
rect 25900 22708 25956 22718
rect 25900 22260 25956 22652
rect 25900 22166 25956 22204
rect 26012 22258 26068 22270
rect 26012 22206 26014 22258
rect 26066 22206 26068 22258
rect 24220 21746 24276 21756
rect 25676 21746 25732 21756
rect 25564 21698 25620 21710
rect 25564 21646 25566 21698
rect 25618 21646 25620 21698
rect 23996 21586 24052 21598
rect 23996 21534 23998 21586
rect 24050 21534 24052 21586
rect 23996 20804 24052 21534
rect 24332 21588 24388 21598
rect 24332 21026 24388 21532
rect 25228 21588 25284 21598
rect 25228 21494 25284 21532
rect 25564 21364 25620 21646
rect 26012 21700 26068 22206
rect 26012 21634 26068 21644
rect 25564 21298 25620 21308
rect 25228 21252 25284 21262
rect 24522 21196 24786 21206
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24522 21130 24786 21140
rect 24332 20974 24334 21026
rect 24386 20974 24388 21026
rect 24332 20962 24388 20974
rect 24108 20804 24164 20814
rect 23996 20802 24164 20804
rect 23996 20750 24110 20802
rect 24162 20750 24164 20802
rect 23996 20748 24164 20750
rect 23884 20178 23940 20188
rect 23324 19966 23326 20018
rect 23378 19966 23380 20018
rect 23324 19954 23380 19966
rect 23548 20018 23604 20030
rect 23548 19966 23550 20018
rect 23602 19966 23604 20018
rect 23548 19796 23604 19966
rect 23772 19796 23828 20076
rect 24108 20020 24164 20748
rect 24892 20692 24948 20702
rect 24444 20690 24948 20692
rect 24444 20638 24894 20690
rect 24946 20638 24948 20690
rect 24444 20636 24948 20638
rect 24332 20244 24388 20254
rect 24444 20244 24500 20636
rect 24892 20626 24948 20636
rect 25228 20690 25284 21196
rect 25228 20638 25230 20690
rect 25282 20638 25284 20690
rect 25228 20626 25284 20638
rect 26012 20692 26068 20702
rect 26124 20692 26180 23102
rect 26012 20690 26180 20692
rect 26012 20638 26014 20690
rect 26066 20638 26180 20690
rect 26012 20636 26180 20638
rect 24332 20242 24500 20244
rect 24332 20190 24334 20242
rect 24386 20190 24500 20242
rect 24332 20188 24500 20190
rect 24332 20178 24388 20188
rect 25564 20132 25620 20142
rect 25564 20038 25620 20076
rect 25228 20020 25284 20030
rect 24164 19964 24276 20020
rect 24108 19926 24164 19964
rect 23772 19740 24164 19796
rect 23548 19730 23604 19740
rect 23212 19182 23214 19234
rect 23266 19182 23268 19234
rect 23212 19170 23268 19182
rect 23772 19234 23828 19246
rect 23996 19236 24052 19246
rect 23772 19182 23774 19234
rect 23826 19182 23828 19234
rect 23436 19124 23492 19134
rect 23772 19124 23828 19182
rect 23436 19122 23828 19124
rect 23436 19070 23438 19122
rect 23490 19070 23828 19122
rect 23436 19068 23828 19070
rect 23884 19180 23996 19236
rect 23436 19058 23492 19068
rect 23324 18450 23380 18462
rect 23324 18398 23326 18450
rect 23378 18398 23380 18450
rect 23324 18340 23380 18398
rect 23324 18274 23380 18284
rect 23548 17780 23604 19068
rect 23884 19012 23940 19180
rect 23996 19142 24052 19180
rect 24108 19234 24164 19740
rect 24108 19182 24110 19234
rect 24162 19182 24164 19234
rect 24108 19170 24164 19182
rect 24220 19236 24276 19964
rect 24892 20018 25284 20020
rect 24892 19966 25230 20018
rect 25282 19966 25284 20018
rect 24892 19964 25284 19966
rect 24522 19628 24786 19638
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24522 19562 24786 19572
rect 24780 19460 24836 19470
rect 24892 19460 24948 19964
rect 25228 19954 25284 19964
rect 24780 19458 24948 19460
rect 24780 19406 24782 19458
rect 24834 19406 24948 19458
rect 24780 19404 24948 19406
rect 24780 19394 24836 19404
rect 25900 19348 25956 19358
rect 24332 19236 24388 19246
rect 24220 19234 24388 19236
rect 24220 19182 24334 19234
rect 24386 19182 24388 19234
rect 24220 19180 24388 19182
rect 24332 19170 24388 19180
rect 25900 19234 25956 19292
rect 25900 19182 25902 19234
rect 25954 19182 25956 19234
rect 25900 19170 25956 19182
rect 23660 18956 23940 19012
rect 25228 19010 25284 19022
rect 25228 18958 25230 19010
rect 25282 18958 25284 19010
rect 23660 18674 23716 18956
rect 23660 18622 23662 18674
rect 23714 18622 23716 18674
rect 23660 18610 23716 18622
rect 24332 18562 24388 18574
rect 24332 18510 24334 18562
rect 24386 18510 24388 18562
rect 24108 18452 24164 18462
rect 24108 18358 24164 18396
rect 24332 18340 24388 18510
rect 23548 17714 23604 17724
rect 24220 17780 24276 17790
rect 22988 17602 23044 17612
rect 23436 17556 23492 17566
rect 23772 17556 23828 17566
rect 23436 17554 23716 17556
rect 23436 17502 23438 17554
rect 23490 17502 23716 17554
rect 23436 17500 23716 17502
rect 23436 17490 23492 17500
rect 23100 17444 23156 17454
rect 23324 17444 23380 17454
rect 23100 17442 23324 17444
rect 23100 17390 23102 17442
rect 23154 17390 23324 17442
rect 23100 17388 23324 17390
rect 23100 17378 23156 17388
rect 22876 16942 22878 16994
rect 22930 16942 22932 16994
rect 22876 16884 22932 16942
rect 22876 16818 22932 16828
rect 23212 16994 23268 17006
rect 23212 16942 23214 16994
rect 23266 16942 23268 16994
rect 22652 16706 22708 16716
rect 22316 16268 23044 16324
rect 22316 15428 22372 15438
rect 22316 15316 22372 15372
rect 22652 15316 22708 15326
rect 22316 15314 22708 15316
rect 22316 15262 22318 15314
rect 22370 15262 22654 15314
rect 22706 15262 22708 15314
rect 22316 15260 22708 15262
rect 22316 15250 22372 15260
rect 22652 15250 22708 15260
rect 22204 14466 22260 14476
rect 22876 14530 22932 16268
rect 22988 16210 23044 16268
rect 22988 16158 22990 16210
rect 23042 16158 23044 16210
rect 22988 16146 23044 16158
rect 23212 16212 23268 16942
rect 23212 16146 23268 16156
rect 23324 16098 23380 17388
rect 23660 17108 23716 17500
rect 23772 17462 23828 17500
rect 23660 17014 23716 17052
rect 23884 16884 23940 16894
rect 23324 16046 23326 16098
rect 23378 16046 23380 16098
rect 23324 16034 23380 16046
rect 23772 16100 23828 16110
rect 23772 16006 23828 16044
rect 23100 15986 23156 15998
rect 23100 15934 23102 15986
rect 23154 15934 23156 15986
rect 22988 15428 23044 15438
rect 23100 15428 23156 15934
rect 22988 15426 23156 15428
rect 22988 15374 22990 15426
rect 23042 15374 23156 15426
rect 22988 15372 23156 15374
rect 23660 15540 23716 15550
rect 22988 15204 23044 15372
rect 22988 15138 23044 15148
rect 23660 15314 23716 15484
rect 23884 15538 23940 16828
rect 24220 16212 24276 17724
rect 24332 17554 24388 18284
rect 25228 18452 25284 18958
rect 25788 18562 25844 18574
rect 25788 18510 25790 18562
rect 25842 18510 25844 18562
rect 25452 18452 25508 18462
rect 24522 18060 24786 18070
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24522 17994 24786 18004
rect 25228 18004 25284 18396
rect 25228 17938 25284 17948
rect 25340 18450 25508 18452
rect 25340 18398 25454 18450
rect 25506 18398 25508 18450
rect 25340 18396 25508 18398
rect 25340 17890 25396 18396
rect 25452 18386 25508 18396
rect 25340 17838 25342 17890
rect 25394 17838 25396 17890
rect 25340 17826 25396 17838
rect 25788 17780 25844 18510
rect 25788 17714 25844 17724
rect 24892 17668 24948 17678
rect 25564 17668 25620 17678
rect 24948 17612 25060 17668
rect 24892 17574 24948 17612
rect 24332 17502 24334 17554
rect 24386 17502 24388 17554
rect 24332 17490 24388 17502
rect 24668 17554 24724 17566
rect 24668 17502 24670 17554
rect 24722 17502 24724 17554
rect 24668 17444 24724 17502
rect 24668 17378 24724 17388
rect 24892 16884 24948 16894
rect 24522 16492 24786 16502
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24522 16426 24786 16436
rect 24444 16212 24500 16222
rect 24892 16212 24948 16828
rect 24220 16210 24500 16212
rect 24220 16158 24446 16210
rect 24498 16158 24500 16210
rect 24220 16156 24500 16158
rect 24444 16146 24500 16156
rect 24668 16156 24948 16212
rect 24668 16098 24724 16156
rect 24668 16046 24670 16098
rect 24722 16046 24724 16098
rect 24668 16034 24724 16046
rect 25004 16100 25060 17612
rect 25564 17574 25620 17612
rect 25900 17554 25956 17566
rect 25900 17502 25902 17554
rect 25954 17502 25956 17554
rect 25004 16006 25060 16044
rect 25116 17444 25172 17454
rect 24556 15988 24612 15998
rect 23996 15876 24052 15886
rect 23996 15874 24276 15876
rect 23996 15822 23998 15874
rect 24050 15822 24276 15874
rect 23996 15820 24276 15822
rect 23996 15810 24052 15820
rect 23884 15486 23886 15538
rect 23938 15486 23940 15538
rect 23884 15474 23940 15486
rect 24220 15426 24276 15820
rect 24556 15538 24612 15932
rect 24892 15986 24948 15998
rect 24892 15934 24894 15986
rect 24946 15934 24948 15986
rect 24892 15876 24948 15934
rect 25116 15876 25172 17388
rect 25228 17444 25284 17454
rect 25900 17444 25956 17502
rect 25228 17442 25396 17444
rect 25228 17390 25230 17442
rect 25282 17390 25396 17442
rect 25228 17388 25396 17390
rect 25228 17378 25284 17388
rect 25340 16994 25396 17388
rect 25900 17378 25956 17388
rect 25788 17220 25844 17230
rect 25676 17108 25732 17118
rect 25676 17014 25732 17052
rect 25340 16942 25342 16994
rect 25394 16942 25396 16994
rect 25340 16930 25396 16942
rect 25452 15988 25508 15998
rect 25676 15988 25732 15998
rect 25452 15986 25732 15988
rect 25452 15934 25454 15986
rect 25506 15934 25678 15986
rect 25730 15934 25732 15986
rect 25452 15932 25732 15934
rect 25452 15922 25508 15932
rect 25676 15922 25732 15932
rect 24892 15820 25172 15876
rect 24556 15486 24558 15538
rect 24610 15486 24612 15538
rect 24556 15474 24612 15486
rect 25564 15652 25620 15662
rect 24220 15374 24222 15426
rect 24274 15374 24276 15426
rect 24220 15362 24276 15374
rect 25564 15426 25620 15596
rect 25564 15374 25566 15426
rect 25618 15374 25620 15426
rect 25564 15362 25620 15374
rect 23660 15262 23662 15314
rect 23714 15262 23716 15314
rect 23660 15148 23716 15262
rect 25676 15316 25732 15326
rect 25788 15316 25844 17164
rect 26012 16884 26068 20636
rect 26124 19348 26180 19358
rect 26124 18562 26180 19292
rect 26124 18510 26126 18562
rect 26178 18510 26180 18562
rect 26124 18498 26180 18510
rect 26236 19010 26292 23884
rect 26348 23874 26404 23884
rect 26572 23940 26628 23950
rect 26572 23846 26628 23884
rect 26684 23938 26740 24782
rect 26796 24948 26852 24958
rect 26796 24276 26852 24892
rect 26796 24210 26852 24220
rect 26684 23886 26686 23938
rect 26738 23886 26740 23938
rect 26460 23380 26516 23390
rect 26684 23380 26740 23886
rect 26460 23378 26740 23380
rect 26460 23326 26462 23378
rect 26514 23326 26740 23378
rect 26460 23324 26740 23326
rect 26460 23314 26516 23324
rect 26460 22260 26516 22270
rect 26796 22260 26852 22270
rect 26460 22258 26852 22260
rect 26460 22206 26462 22258
rect 26514 22206 26798 22258
rect 26850 22206 26852 22258
rect 26460 22204 26852 22206
rect 26460 22194 26516 22204
rect 26796 22194 26852 22204
rect 26572 22036 26628 22046
rect 26460 21812 26516 21822
rect 26348 21700 26404 21710
rect 26348 20692 26404 21644
rect 26460 21698 26516 21756
rect 26460 21646 26462 21698
rect 26514 21646 26516 21698
rect 26460 21634 26516 21646
rect 26572 21588 26628 21980
rect 26684 21700 26740 21710
rect 26684 21606 26740 21644
rect 26572 21494 26628 21532
rect 27020 21476 27076 26012
rect 27468 25620 27524 27806
rect 27804 27860 27860 27870
rect 27804 27766 27860 27804
rect 27804 26292 27860 26302
rect 27916 26292 27972 28476
rect 28252 27860 28308 27870
rect 28588 27860 28644 27870
rect 28252 27858 28644 27860
rect 28252 27806 28254 27858
rect 28306 27806 28590 27858
rect 28642 27806 28644 27858
rect 28252 27804 28644 27806
rect 28252 27794 28308 27804
rect 28588 27794 28644 27804
rect 28252 26962 28308 26974
rect 28252 26910 28254 26962
rect 28306 26910 28308 26962
rect 28140 26516 28196 26526
rect 28252 26516 28308 26910
rect 28588 26964 28644 26974
rect 28700 26964 28756 30940
rect 28812 30930 28868 30940
rect 28924 28082 28980 36428
rect 29260 36418 29316 36428
rect 29708 36370 29764 37660
rect 29708 36318 29710 36370
rect 29762 36318 29764 36370
rect 29708 36306 29764 36318
rect 29036 36260 29092 36270
rect 29036 36166 29092 36204
rect 29820 36260 29876 37772
rect 30828 37716 30884 37772
rect 30828 37660 31108 37716
rect 29820 36194 29876 36204
rect 30044 36370 30100 36382
rect 30044 36318 30046 36370
rect 30098 36318 30100 36370
rect 29184 36092 29448 36102
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29184 36026 29448 36036
rect 29184 34524 29448 34534
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29184 34458 29448 34468
rect 30044 33572 30100 36318
rect 30716 36370 30772 36382
rect 30716 36318 30718 36370
rect 30770 36318 30772 36370
rect 30380 36260 30436 36270
rect 30380 36166 30436 36204
rect 30716 35364 30772 36318
rect 31052 36370 31108 37660
rect 31052 36318 31054 36370
rect 31106 36318 31108 36370
rect 31052 36306 31108 36318
rect 31164 36372 31220 37772
rect 31612 36932 31668 39200
rect 32284 37826 32340 39200
rect 32284 37774 32286 37826
rect 32338 37774 32340 37826
rect 32284 37762 32340 37774
rect 31612 36866 31668 36876
rect 32844 36932 32900 36942
rect 32396 36484 32452 36494
rect 32284 36482 32452 36484
rect 32284 36430 32398 36482
rect 32450 36430 32452 36482
rect 32284 36428 32452 36430
rect 31164 36306 31220 36316
rect 31388 36370 31444 36382
rect 31388 36318 31390 36370
rect 31442 36318 31444 36370
rect 30716 35298 30772 35308
rect 30044 33506 30100 33516
rect 29184 32956 29448 32966
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29184 32890 29448 32900
rect 30380 31668 30436 31678
rect 29184 31388 29448 31398
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29184 31322 29448 31332
rect 29932 30324 29988 30334
rect 29820 30268 29932 30324
rect 29184 29820 29448 29830
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29184 29754 29448 29764
rect 29184 28252 29448 28262
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29184 28186 29448 28196
rect 28924 28030 28926 28082
rect 28978 28030 28980 28082
rect 28924 28018 28980 28030
rect 28588 26962 28756 26964
rect 28588 26910 28590 26962
rect 28642 26910 28756 26962
rect 28588 26908 28756 26910
rect 28588 26898 28644 26908
rect 29708 26852 29764 26862
rect 29184 26684 29448 26694
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29184 26618 29448 26628
rect 28140 26514 28308 26516
rect 28140 26462 28142 26514
rect 28194 26462 28308 26514
rect 28140 26460 28308 26462
rect 28140 26450 28196 26460
rect 27804 26290 28420 26292
rect 27804 26238 27806 26290
rect 27858 26238 28420 26290
rect 27804 26236 28420 26238
rect 27804 26226 27860 26236
rect 27244 25564 27524 25620
rect 27580 26178 27636 26190
rect 27580 26126 27582 26178
rect 27634 26126 27636 26178
rect 27580 25620 27636 26126
rect 27132 24948 27188 24958
rect 27244 24948 27300 25564
rect 27580 25554 27636 25564
rect 27356 25396 27412 25406
rect 27692 25396 27748 25406
rect 27356 25394 27748 25396
rect 27356 25342 27358 25394
rect 27410 25342 27694 25394
rect 27746 25342 27748 25394
rect 27356 25340 27748 25342
rect 27356 25330 27412 25340
rect 27692 25330 27748 25340
rect 28028 25396 28084 25406
rect 28028 25302 28084 25340
rect 27188 24892 27300 24948
rect 27132 24882 27188 24892
rect 27804 24834 27860 24846
rect 27804 24782 27806 24834
rect 27858 24782 27860 24834
rect 27132 24724 27188 24734
rect 27468 24724 27524 24734
rect 27132 24722 27524 24724
rect 27132 24670 27134 24722
rect 27186 24670 27470 24722
rect 27522 24670 27524 24722
rect 27132 24668 27524 24670
rect 27132 24658 27188 24668
rect 27468 24658 27524 24668
rect 27804 24164 27860 24782
rect 28364 24724 28420 26236
rect 29184 25116 29448 25126
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29184 25050 29448 25060
rect 29372 24948 29428 24958
rect 29708 24948 29764 26796
rect 29372 24946 29764 24948
rect 29372 24894 29374 24946
rect 29426 24894 29764 24946
rect 29372 24892 29764 24894
rect 29372 24882 29428 24892
rect 29820 24836 29876 30268
rect 29932 30258 29988 30268
rect 30268 29428 30324 29438
rect 29484 24780 29876 24836
rect 29932 27188 29988 27198
rect 28252 24722 28420 24724
rect 28252 24670 28366 24722
rect 28418 24670 28420 24722
rect 28252 24668 28420 24670
rect 28140 24612 28196 24622
rect 28140 24518 28196 24556
rect 28140 24164 28196 24174
rect 28252 24164 28308 24668
rect 28364 24658 28420 24668
rect 28700 24724 28756 24734
rect 29036 24724 29092 24734
rect 28700 24722 29092 24724
rect 28700 24670 28702 24722
rect 28754 24670 29038 24722
rect 29090 24670 29092 24722
rect 28700 24668 29092 24670
rect 28700 24658 28756 24668
rect 29036 24658 29092 24668
rect 27804 24098 27860 24108
rect 28028 24162 28308 24164
rect 28028 24110 28142 24162
rect 28194 24110 28308 24162
rect 28028 24108 28308 24110
rect 27916 23938 27972 23950
rect 27916 23886 27918 23938
rect 27970 23886 27972 23938
rect 27132 23716 27188 23726
rect 27132 23714 27300 23716
rect 27132 23662 27134 23714
rect 27186 23662 27300 23714
rect 27132 23660 27300 23662
rect 27132 23650 27188 23660
rect 27244 23266 27300 23660
rect 27916 23604 27972 23886
rect 27916 23538 27972 23548
rect 27580 23380 27636 23390
rect 27580 23286 27636 23324
rect 27916 23380 27972 23390
rect 28028 23380 28084 24108
rect 28140 24098 28196 24108
rect 28476 23828 28532 23838
rect 28476 23734 28532 23772
rect 29148 23828 29204 23838
rect 29148 23734 29204 23772
rect 29484 23826 29540 24780
rect 29484 23774 29486 23826
rect 29538 23774 29540 23826
rect 29484 23762 29540 23774
rect 29184 23548 29448 23558
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29184 23482 29448 23492
rect 27916 23378 28084 23380
rect 27916 23326 27918 23378
rect 27970 23326 28084 23378
rect 27916 23324 28084 23326
rect 27916 23314 27972 23324
rect 27244 23214 27246 23266
rect 27298 23214 27300 23266
rect 27244 23202 27300 23214
rect 29372 23266 29428 23278
rect 29372 23214 29374 23266
rect 29426 23214 29428 23266
rect 28252 23154 28308 23166
rect 28252 23102 28254 23154
rect 28306 23102 28308 23154
rect 27804 22596 27860 22606
rect 27132 22260 27188 22270
rect 27468 22260 27524 22270
rect 27132 22166 27188 22204
rect 27244 22258 27524 22260
rect 27244 22206 27470 22258
rect 27522 22206 27524 22258
rect 27244 22204 27524 22206
rect 27132 21812 27188 21822
rect 27244 21812 27300 22204
rect 27468 22194 27524 22204
rect 27804 22258 27860 22540
rect 28252 22260 28308 23102
rect 28700 23156 28756 23166
rect 27804 22206 27806 22258
rect 27858 22206 27860 22258
rect 27804 22194 27860 22206
rect 28140 22258 28308 22260
rect 28140 22206 28254 22258
rect 28306 22206 28308 22258
rect 28140 22204 28308 22206
rect 27132 21810 27300 21812
rect 27132 21758 27134 21810
rect 27186 21758 27300 21810
rect 27132 21756 27300 21758
rect 27468 21812 27524 21822
rect 27132 21746 27188 21756
rect 27468 21586 27524 21756
rect 27804 21700 27860 21710
rect 27804 21606 27860 21644
rect 27468 21534 27470 21586
rect 27522 21534 27524 21586
rect 27468 21522 27524 21534
rect 27692 21586 27748 21598
rect 27692 21534 27694 21586
rect 27746 21534 27748 21586
rect 27020 21410 27076 21420
rect 27692 20916 27748 21534
rect 27468 20860 27748 20916
rect 26348 20598 26404 20636
rect 27132 20692 27188 20702
rect 27132 20130 27188 20636
rect 27468 20580 27524 20860
rect 27692 20692 27748 20702
rect 27468 20514 27524 20524
rect 27580 20690 27748 20692
rect 27580 20638 27694 20690
rect 27746 20638 27748 20690
rect 27580 20636 27748 20638
rect 27580 20242 27636 20636
rect 27692 20626 27748 20636
rect 28028 20692 28084 20702
rect 28028 20598 28084 20636
rect 27580 20190 27582 20242
rect 27634 20190 27636 20242
rect 27580 20178 27636 20190
rect 28140 20188 28196 22204
rect 28252 22194 28308 22204
rect 28588 22372 28644 22382
rect 28588 22258 28644 22316
rect 28588 22206 28590 22258
rect 28642 22206 28644 22258
rect 28588 22194 28644 22206
rect 28252 21588 28308 21598
rect 28588 21588 28644 21598
rect 28252 21586 28644 21588
rect 28252 21534 28254 21586
rect 28306 21534 28590 21586
rect 28642 21534 28644 21586
rect 28252 21532 28644 21534
rect 28252 21522 28308 21532
rect 28588 21522 28644 21532
rect 28140 20132 28420 20188
rect 27132 20078 27134 20130
rect 27186 20078 27188 20130
rect 27132 20066 27188 20078
rect 26908 20018 26964 20030
rect 26908 19966 26910 20018
rect 26962 19966 26964 20018
rect 26572 19348 26628 19358
rect 26572 19234 26628 19292
rect 26572 19182 26574 19234
rect 26626 19182 26628 19234
rect 26572 19170 26628 19182
rect 26908 19236 26964 19966
rect 27020 20020 27076 20030
rect 27020 19796 27076 19964
rect 27020 19730 27076 19740
rect 28252 20018 28308 20030
rect 28252 19966 28254 20018
rect 28306 19966 28308 20018
rect 27356 19236 27412 19246
rect 26908 19234 27412 19236
rect 26908 19182 27358 19234
rect 27410 19182 27412 19234
rect 26908 19180 27412 19182
rect 26908 19122 26964 19180
rect 26908 19070 26910 19122
rect 26962 19070 26964 19122
rect 26908 19058 26964 19070
rect 26236 18958 26238 19010
rect 26290 18958 26292 19010
rect 26124 17556 26180 17566
rect 26124 17462 26180 17500
rect 26236 17444 26292 18958
rect 26460 18562 26516 18574
rect 27356 18564 27412 19180
rect 27580 19236 27636 19246
rect 27580 19142 27636 19180
rect 27692 19122 27748 19134
rect 27692 19070 27694 19122
rect 27746 19070 27748 19122
rect 26460 18510 26462 18562
rect 26514 18510 26516 18562
rect 26348 17892 26404 17902
rect 26348 17778 26404 17836
rect 26348 17726 26350 17778
rect 26402 17726 26404 17778
rect 26348 17714 26404 17726
rect 26236 17388 26404 17444
rect 26236 16884 26292 16894
rect 26012 16882 26292 16884
rect 26012 16830 26238 16882
rect 26290 16830 26292 16882
rect 26012 16828 26292 16830
rect 26012 15874 26068 15886
rect 26012 15822 26014 15874
rect 26066 15822 26068 15874
rect 25900 15428 25956 15438
rect 25900 15334 25956 15372
rect 25732 15260 25844 15316
rect 24892 15204 24948 15214
rect 23660 15092 24276 15148
rect 23100 14588 23380 14644
rect 22876 14478 22878 14530
rect 22930 14478 22932 14530
rect 22316 14420 22372 14430
rect 22372 14364 22484 14420
rect 22316 14354 22372 14364
rect 22316 13972 22372 13982
rect 22316 13878 22372 13916
rect 22428 13748 22484 14364
rect 21868 13580 22148 13636
rect 22316 13692 22484 13748
rect 21420 13076 21476 13086
rect 21420 12982 21476 13020
rect 21196 12236 21476 12292
rect 21308 12066 21364 12078
rect 21308 12014 21310 12066
rect 21362 12014 21364 12066
rect 21308 11394 21364 12014
rect 21308 11342 21310 11394
rect 21362 11342 21364 11394
rect 21308 10164 21364 11342
rect 21308 10098 21364 10108
rect 21420 11284 21476 12236
rect 20860 9772 21364 9828
rect 20636 9662 20638 9714
rect 20690 9662 20692 9714
rect 20636 9650 20692 9662
rect 20860 9602 20916 9614
rect 20860 9550 20862 9602
rect 20914 9550 20916 9602
rect 19860 9436 20124 9446
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 19860 9370 20124 9380
rect 19740 9156 19796 9166
rect 19740 9062 19796 9100
rect 19860 7868 20124 7878
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 19860 7802 20124 7812
rect 19628 7586 19796 7588
rect 19628 7534 19630 7586
rect 19682 7534 19796 7586
rect 19628 7532 19796 7534
rect 19628 7522 19684 7532
rect 19292 3502 19294 3554
rect 19346 3502 19348 3554
rect 19292 3490 19348 3502
rect 19740 3444 19796 7532
rect 19860 6300 20124 6310
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 19860 6234 20124 6244
rect 20860 5908 20916 9550
rect 20860 5842 20916 5852
rect 19860 4732 20124 4742
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 19860 4666 20124 4676
rect 20412 4228 20468 4238
rect 20188 4226 20468 4228
rect 20188 4174 20414 4226
rect 20466 4174 20468 4226
rect 20188 4172 20468 4174
rect 20188 3554 20244 4172
rect 20412 4162 20468 4172
rect 20188 3502 20190 3554
rect 20242 3502 20244 3554
rect 19852 3444 19908 3454
rect 19740 3442 19908 3444
rect 19740 3390 19854 3442
rect 19906 3390 19908 3442
rect 19740 3388 19908 3390
rect 19852 3378 19908 3388
rect 18508 3276 18788 3332
rect 18844 3330 18900 3342
rect 18844 3278 18846 3330
rect 18898 3278 18900 3330
rect 18844 800 18900 3278
rect 19516 3330 19572 3342
rect 19516 3278 19518 3330
rect 19570 3278 19572 3330
rect 19516 800 19572 3278
rect 19860 3164 20124 3174
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 19860 3098 20124 3108
rect 20188 800 20244 3502
rect 21308 3554 21364 9772
rect 21308 3502 21310 3554
rect 21362 3502 21364 3554
rect 21308 3490 21364 3502
rect 21420 3388 21476 11228
rect 21756 11284 21812 11294
rect 21756 10724 21812 11228
rect 21756 10630 21812 10668
rect 21868 10500 21924 13580
rect 21980 12962 22036 12974
rect 21980 12910 21982 12962
rect 22034 12910 22036 12962
rect 21980 12740 22036 12910
rect 22092 12964 22148 12974
rect 22092 12870 22148 12908
rect 22204 12964 22260 12974
rect 22316 12964 22372 13692
rect 22876 13634 22932 14478
rect 22876 13582 22878 13634
rect 22930 13582 22932 13634
rect 22876 13524 22932 13582
rect 22204 12962 22372 12964
rect 22204 12910 22206 12962
rect 22258 12910 22372 12962
rect 22204 12908 22372 12910
rect 22540 13468 22932 13524
rect 22988 14532 23044 14542
rect 22204 12898 22260 12908
rect 22540 12740 22596 13468
rect 22988 13412 23044 14476
rect 23100 14530 23156 14588
rect 23100 14478 23102 14530
rect 23154 14478 23156 14530
rect 23100 14466 23156 14478
rect 23212 14420 23268 14458
rect 23212 13858 23268 14364
rect 23212 13806 23214 13858
rect 23266 13806 23268 13858
rect 23212 13794 23268 13806
rect 22652 13356 23044 13412
rect 23100 13746 23156 13758
rect 23100 13694 23102 13746
rect 23154 13694 23156 13746
rect 23100 13524 23156 13694
rect 22652 12962 22708 13356
rect 23100 13076 23156 13468
rect 23100 13020 23268 13076
rect 22652 12910 22654 12962
rect 22706 12910 22708 12962
rect 22652 12898 22708 12910
rect 22876 12852 22932 12862
rect 23100 12852 23156 12862
rect 22876 12850 23156 12852
rect 22876 12798 22878 12850
rect 22930 12798 23102 12850
rect 23154 12798 23156 12850
rect 22876 12796 23156 12798
rect 22876 12786 22932 12796
rect 23100 12786 23156 12796
rect 21980 12684 22596 12740
rect 23100 12180 23156 12190
rect 23212 12180 23268 13020
rect 23156 12124 23268 12180
rect 23100 12114 23156 12124
rect 23212 11732 23268 11742
rect 22092 11396 22148 11406
rect 22092 11302 22148 11340
rect 21756 10444 21924 10500
rect 21756 10276 21812 10444
rect 21756 10210 21812 10220
rect 22540 10276 22596 10286
rect 21868 10164 21924 10174
rect 21868 8930 21924 10108
rect 22316 9716 22372 9726
rect 22316 9156 22372 9660
rect 22316 9042 22372 9100
rect 22316 8990 22318 9042
rect 22370 8990 22372 9042
rect 22316 8978 22372 8990
rect 21868 8878 21870 8930
rect 21922 8878 21924 8930
rect 21868 8866 21924 8878
rect 22428 8820 22484 8830
rect 22092 8146 22148 8158
rect 22092 8094 22094 8146
rect 22146 8094 22148 8146
rect 22092 8036 22148 8094
rect 22428 8146 22484 8764
rect 22428 8094 22430 8146
rect 22482 8094 22484 8146
rect 22428 8082 22484 8094
rect 21756 7364 21812 7374
rect 22092 7364 22148 7980
rect 21756 7362 22148 7364
rect 21756 7310 21758 7362
rect 21810 7310 22148 7362
rect 21756 7308 22148 7310
rect 21756 7298 21812 7308
rect 21532 4228 21588 4238
rect 21532 4226 21924 4228
rect 21532 4174 21534 4226
rect 21586 4174 21924 4226
rect 21532 4172 21924 4174
rect 21532 4162 21588 4172
rect 21084 3332 21140 3342
rect 20860 3330 21140 3332
rect 20860 3278 21086 3330
rect 21138 3278 21140 3330
rect 20860 3276 21140 3278
rect 21308 3332 21476 3388
rect 21868 3556 21924 4172
rect 22204 4226 22260 4238
rect 22204 4174 22206 4226
rect 22258 4174 22260 4226
rect 21980 3556 22036 3566
rect 21868 3554 22036 3556
rect 21868 3502 21982 3554
rect 22034 3502 22036 3554
rect 21868 3500 22036 3502
rect 21756 3332 21812 3342
rect 21308 3330 21812 3332
rect 21308 3278 21758 3330
rect 21810 3278 21812 3330
rect 21308 3276 21812 3278
rect 20860 800 20916 3276
rect 21084 3266 21140 3276
rect 21756 3266 21812 3276
rect 21868 3108 21924 3500
rect 21980 3490 22036 3500
rect 21756 3052 21924 3108
rect 21756 2772 21812 3052
rect 21532 2716 21812 2772
rect 21532 800 21588 2716
rect 22204 2548 22260 4174
rect 22428 3444 22484 3454
rect 22540 3444 22596 10220
rect 23212 10164 23268 11676
rect 23324 11620 23380 14588
rect 24220 14642 24276 15092
rect 24522 14924 24786 14934
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24522 14858 24786 14868
rect 24892 14756 24948 15148
rect 24220 14590 24222 14642
rect 24274 14590 24276 14642
rect 24220 14578 24276 14590
rect 24556 14700 24948 14756
rect 24556 14642 24612 14700
rect 24556 14590 24558 14642
rect 24610 14590 24612 14642
rect 24556 14578 24612 14590
rect 23436 14532 23492 14542
rect 23492 14476 23604 14532
rect 23436 14438 23492 14476
rect 23548 13746 23604 14476
rect 24780 14530 24836 14542
rect 24780 14478 24782 14530
rect 24834 14478 24836 14530
rect 24780 14420 24836 14478
rect 25676 14530 25732 15260
rect 25676 14478 25678 14530
rect 25730 14478 25732 14530
rect 25676 14466 25732 14478
rect 25452 14420 25508 14430
rect 24836 14364 24948 14420
rect 24780 14354 24836 14364
rect 23884 14308 23940 14318
rect 23884 14306 24164 14308
rect 23884 14254 23886 14306
rect 23938 14254 24164 14306
rect 23884 14252 24164 14254
rect 23884 14242 23940 14252
rect 24108 13858 24164 14252
rect 24444 13860 24500 13870
rect 24108 13806 24110 13858
rect 24162 13806 24164 13858
rect 24108 13794 24164 13806
rect 24332 13858 24500 13860
rect 24332 13806 24446 13858
rect 24498 13806 24500 13858
rect 24332 13804 24500 13806
rect 23548 13694 23550 13746
rect 23602 13694 23604 13746
rect 23548 13682 23604 13694
rect 23884 13522 23940 13534
rect 23884 13470 23886 13522
rect 23938 13470 23940 13522
rect 23884 12962 23940 13470
rect 23884 12910 23886 12962
rect 23938 12910 23940 12962
rect 23884 12898 23940 12910
rect 23436 12738 23492 12750
rect 24108 12740 24164 12750
rect 23436 12686 23438 12738
rect 23490 12686 23492 12738
rect 23436 12404 23492 12686
rect 23996 12738 24164 12740
rect 23996 12686 24110 12738
rect 24162 12686 24164 12738
rect 23996 12684 24164 12686
rect 23436 12348 23604 12404
rect 23324 11554 23380 11564
rect 23436 12178 23492 12190
rect 23436 12126 23438 12178
rect 23490 12126 23492 12178
rect 22876 9154 22932 9166
rect 22876 9102 22878 9154
rect 22930 9102 22932 9154
rect 22652 9044 22708 9054
rect 22652 9042 22820 9044
rect 22652 8990 22654 9042
rect 22706 8990 22820 9042
rect 22652 8988 22820 8990
rect 22652 8978 22708 8988
rect 22764 7700 22820 8988
rect 22876 8820 22932 9102
rect 23212 9154 23268 10108
rect 23436 9716 23492 12126
rect 23436 9650 23492 9660
rect 23548 9268 23604 12348
rect 23996 10388 24052 12684
rect 24108 12674 24164 12684
rect 24220 12178 24276 12190
rect 24220 12126 24222 12178
rect 24274 12126 24276 12178
rect 24220 11732 24276 12126
rect 24332 11956 24388 13804
rect 24444 13794 24500 13804
rect 24522 13356 24786 13366
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24522 13290 24786 13300
rect 24780 13188 24836 13198
rect 24892 13188 24948 14364
rect 25452 14326 25508 14364
rect 25116 14306 25172 14318
rect 25116 14254 25118 14306
rect 25170 14254 25172 14306
rect 25116 13972 25172 14254
rect 25116 13916 25396 13972
rect 25228 13748 25284 13758
rect 25116 13746 25284 13748
rect 25116 13694 25230 13746
rect 25282 13694 25284 13746
rect 25116 13692 25284 13694
rect 24780 13186 25060 13188
rect 24780 13134 24782 13186
rect 24834 13134 25060 13186
rect 24780 13132 25060 13134
rect 24780 13122 24836 13132
rect 24556 12964 24612 12974
rect 24556 12870 24612 12908
rect 24556 12292 24612 12302
rect 24556 12290 24948 12292
rect 24556 12238 24558 12290
rect 24610 12238 24948 12290
rect 24556 12236 24948 12238
rect 24556 12226 24612 12236
rect 24332 11890 24388 11900
rect 24522 11788 24786 11798
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24522 11722 24786 11732
rect 24220 11666 24276 11676
rect 24220 11508 24276 11518
rect 23996 10322 24052 10332
rect 24108 11452 24220 11508
rect 24108 10164 24164 11452
rect 24220 11414 24276 11452
rect 24892 11396 24948 12236
rect 25004 12180 25060 13132
rect 25116 13186 25172 13692
rect 25228 13682 25284 13692
rect 25116 13134 25118 13186
rect 25170 13134 25172 13186
rect 25116 13122 25172 13134
rect 25228 13524 25284 13534
rect 25004 12114 25060 12124
rect 25228 12178 25284 13468
rect 25340 12964 25396 13916
rect 25564 13860 25620 13870
rect 25564 13766 25620 13804
rect 26012 13412 26068 15822
rect 26236 15652 26292 16828
rect 26236 15586 26292 15596
rect 26348 15426 26404 17388
rect 26460 17220 26516 18510
rect 27244 18562 27412 18564
rect 27244 18510 27358 18562
rect 27410 18510 27412 18562
rect 27244 18508 27412 18510
rect 27244 17666 27300 18508
rect 27356 18498 27412 18508
rect 27580 18564 27636 18574
rect 27692 18564 27748 19070
rect 28140 19124 28196 19134
rect 28140 19030 28196 19068
rect 28028 18676 28084 18686
rect 28252 18676 28308 19966
rect 28028 18674 28308 18676
rect 28028 18622 28030 18674
rect 28082 18622 28308 18674
rect 28028 18620 28308 18622
rect 28028 18610 28084 18620
rect 27580 18562 27748 18564
rect 27580 18510 27582 18562
rect 27634 18510 27748 18562
rect 27580 18508 27748 18510
rect 27468 18450 27524 18462
rect 27468 18398 27470 18450
rect 27522 18398 27524 18450
rect 27468 18340 27524 18398
rect 27468 18274 27524 18284
rect 27244 17614 27246 17666
rect 27298 17614 27300 17666
rect 27244 17602 27300 17614
rect 27468 17668 27524 17678
rect 27580 17668 27636 18508
rect 27468 17666 27636 17668
rect 27468 17614 27470 17666
rect 27522 17614 27636 17666
rect 27468 17612 27636 17614
rect 27356 17554 27412 17566
rect 27356 17502 27358 17554
rect 27410 17502 27412 17554
rect 27132 17444 27188 17454
rect 27356 17444 27412 17502
rect 27188 17388 27412 17444
rect 27132 17378 27188 17388
rect 27468 17332 27524 17612
rect 27916 17556 27972 17566
rect 28252 17556 28308 17566
rect 27916 17554 28308 17556
rect 27916 17502 27918 17554
rect 27970 17502 28254 17554
rect 28306 17502 28308 17554
rect 27916 17500 28308 17502
rect 27916 17490 27972 17500
rect 28252 17490 28308 17500
rect 27244 17276 27524 17332
rect 26460 17164 26964 17220
rect 26572 16996 26628 17006
rect 26572 16902 26628 16940
rect 26908 16884 26964 17164
rect 27244 16996 27300 17276
rect 28364 17220 28420 20132
rect 28588 20132 28644 20142
rect 28588 20038 28644 20076
rect 28588 17668 28644 17678
rect 28588 17554 28644 17612
rect 28588 17502 28590 17554
rect 28642 17502 28644 17554
rect 28588 17490 28644 17502
rect 28364 17154 28420 17164
rect 27244 16902 27300 16940
rect 28364 16994 28420 17006
rect 28364 16942 28366 16994
rect 28418 16942 28420 16994
rect 27132 16884 27188 16894
rect 26908 16882 27076 16884
rect 26908 16830 26910 16882
rect 26962 16830 27076 16882
rect 26908 16828 27076 16830
rect 26908 16818 26964 16828
rect 27020 15652 27076 16828
rect 27132 16790 27188 16828
rect 27692 16884 27748 16894
rect 28028 16884 28084 16894
rect 27692 16882 28084 16884
rect 27692 16830 27694 16882
rect 27746 16830 28030 16882
rect 28082 16830 28084 16882
rect 27692 16828 28084 16830
rect 27692 16818 27748 16828
rect 28028 16818 28084 16828
rect 28364 15876 28420 16942
rect 28700 16884 28756 23100
rect 29036 23156 29092 23166
rect 29036 23062 29092 23100
rect 29372 22820 29428 23214
rect 29372 22148 29428 22764
rect 29596 22708 29652 22718
rect 29596 22482 29652 22652
rect 29596 22430 29598 22482
rect 29650 22430 29652 22482
rect 29596 22418 29652 22430
rect 29820 22372 29876 22382
rect 29820 22278 29876 22316
rect 29932 22260 29988 27132
rect 30268 23380 30324 29372
rect 30380 26852 30436 31612
rect 31388 28532 31444 36318
rect 32172 36372 32228 36382
rect 32172 36278 32228 36316
rect 31388 28466 31444 28476
rect 31500 34804 31556 34814
rect 30380 26786 30436 26796
rect 30492 27748 30548 27758
rect 30492 23380 30548 27692
rect 30268 23314 30324 23324
rect 30380 23324 30548 23380
rect 31276 24724 31332 24734
rect 31276 23378 31332 24668
rect 31276 23326 31278 23378
rect 31330 23326 31332 23378
rect 30380 23268 30436 23324
rect 31276 23314 31332 23326
rect 30380 23202 30436 23212
rect 30604 23268 30660 23278
rect 30604 23174 30660 23212
rect 30268 23156 30324 23166
rect 30156 23154 30324 23156
rect 30156 23102 30270 23154
rect 30322 23102 30324 23154
rect 30156 23100 30324 23102
rect 30156 22594 30212 23100
rect 30268 23090 30324 23100
rect 31052 23154 31108 23166
rect 31052 23102 31054 23154
rect 31106 23102 31108 23154
rect 30716 22820 30772 22830
rect 30156 22542 30158 22594
rect 30210 22542 30212 22594
rect 30156 22530 30212 22542
rect 30492 22708 30548 22718
rect 30492 22482 30548 22652
rect 30716 22594 30772 22764
rect 30716 22542 30718 22594
rect 30770 22542 30772 22594
rect 30716 22530 30772 22542
rect 31052 22594 31108 23102
rect 31388 22820 31444 22830
rect 31052 22542 31054 22594
rect 31106 22542 31108 22594
rect 31052 22530 31108 22542
rect 31276 22764 31388 22820
rect 30492 22430 30494 22482
rect 30546 22430 30548 22482
rect 30492 22418 30548 22430
rect 29932 22194 29988 22204
rect 29372 22092 29652 22148
rect 29184 21980 29448 21990
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29184 21914 29448 21924
rect 28924 21812 28980 21822
rect 28924 21718 28980 21756
rect 29484 21028 29540 21038
rect 29596 21028 29652 22092
rect 30156 21700 30212 21710
rect 30156 21606 30212 21644
rect 29932 21588 29988 21598
rect 29932 21586 30100 21588
rect 29932 21534 29934 21586
rect 29986 21534 30100 21586
rect 29932 21532 30100 21534
rect 29932 21522 29988 21532
rect 29484 21026 29652 21028
rect 29484 20974 29486 21026
rect 29538 20974 29652 21026
rect 29484 20972 29652 20974
rect 29932 21028 29988 21038
rect 30044 21028 30100 21532
rect 30156 21028 30212 21038
rect 30044 21026 30212 21028
rect 30044 20974 30158 21026
rect 30210 20974 30212 21026
rect 30044 20972 30212 20974
rect 31276 21028 31332 22764
rect 31388 22754 31444 22764
rect 31388 22370 31444 22382
rect 31388 22318 31390 22370
rect 31442 22318 31444 22370
rect 31388 22148 31444 22318
rect 31388 22082 31444 22092
rect 31500 21252 31556 34748
rect 32284 33684 32340 36428
rect 32396 36418 32452 36428
rect 32844 36370 32900 36876
rect 32844 36318 32846 36370
rect 32898 36318 32900 36370
rect 32844 36306 32900 36318
rect 32956 36372 33012 39200
rect 33516 37826 33572 37838
rect 33516 37774 33518 37826
rect 33570 37774 33572 37826
rect 32956 36306 33012 36316
rect 33068 36482 33124 36494
rect 33068 36430 33070 36482
rect 33122 36430 33124 36482
rect 32284 33618 32340 33628
rect 32508 35588 32564 35598
rect 33068 35588 33124 36430
rect 33516 36370 33572 37774
rect 33628 37714 33684 39200
rect 33628 37662 33630 37714
rect 33682 37662 33684 37714
rect 33628 37650 33684 37662
rect 33846 36876 34110 36886
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 33846 36810 34110 36820
rect 33516 36318 33518 36370
rect 33570 36318 33572 36370
rect 33516 36306 33572 36318
rect 33852 36370 33908 36382
rect 33852 36318 33854 36370
rect 33906 36318 33908 36370
rect 33740 35924 33796 35934
rect 33740 35830 33796 35868
rect 32508 35586 33124 35588
rect 32508 35534 32510 35586
rect 32562 35534 33124 35586
rect 32508 35532 33124 35534
rect 33180 35588 33236 35598
rect 32172 33124 32228 33134
rect 32060 23156 32116 23166
rect 31948 23154 32116 23156
rect 31948 23102 32062 23154
rect 32114 23102 32116 23154
rect 31948 23100 32116 23102
rect 31948 22594 32004 23100
rect 32060 23090 32116 23100
rect 31948 22542 31950 22594
rect 32002 22542 32004 22594
rect 31948 22530 32004 22542
rect 31500 21186 31556 21196
rect 31612 22372 31668 22382
rect 31388 21028 31444 21038
rect 31276 21026 31444 21028
rect 31276 20974 31390 21026
rect 31442 20974 31444 21026
rect 31276 20972 31444 20974
rect 29484 20962 29540 20972
rect 29260 20804 29316 20814
rect 29036 20748 29260 20804
rect 29036 20020 29092 20748
rect 29260 20710 29316 20748
rect 29820 20578 29876 20590
rect 29820 20526 29822 20578
rect 29874 20526 29876 20578
rect 29184 20412 29448 20422
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29184 20346 29448 20356
rect 29820 20130 29876 20526
rect 29932 20188 29988 20972
rect 30156 20962 30212 20972
rect 31388 20962 31444 20972
rect 30492 20916 30548 20926
rect 30492 20822 30548 20860
rect 31612 20916 31668 22316
rect 32172 22260 32228 33068
rect 32508 31948 32564 35532
rect 33180 35494 33236 35532
rect 33852 35588 33908 36318
rect 34188 36372 34244 36382
rect 34188 36278 34244 36316
rect 34300 35924 34356 39200
rect 34860 37714 34916 37726
rect 34860 37662 34862 37714
rect 34914 37662 34916 37714
rect 34412 36482 34468 36494
rect 34412 36430 34414 36482
rect 34466 36430 34468 36482
rect 34412 36148 34468 36430
rect 34860 36370 34916 37662
rect 34860 36318 34862 36370
rect 34914 36318 34916 36370
rect 34860 36306 34916 36318
rect 34972 36372 35028 39200
rect 35644 37828 35700 39200
rect 35644 37772 36260 37828
rect 36204 36708 36260 37772
rect 36316 36932 36372 39200
rect 36316 36866 36372 36876
rect 37324 36932 37380 36942
rect 36204 36652 36708 36708
rect 36204 36482 36260 36494
rect 36204 36430 36206 36482
rect 36258 36430 36260 36482
rect 34972 36306 35028 36316
rect 35196 36370 35252 36382
rect 35196 36318 35198 36370
rect 35250 36318 35252 36370
rect 34412 36082 34468 36092
rect 34524 35924 34580 35934
rect 34300 35922 34580 35924
rect 34300 35870 34526 35922
rect 34578 35870 34580 35922
rect 34300 35868 34580 35870
rect 34524 35858 34580 35868
rect 34748 35698 34804 35710
rect 34748 35646 34750 35698
rect 34802 35646 34804 35698
rect 33852 35522 33908 35532
rect 34188 35588 34244 35598
rect 34748 35588 34804 35646
rect 34188 35586 34804 35588
rect 34188 35534 34190 35586
rect 34242 35534 34804 35586
rect 34188 35532 34804 35534
rect 35196 35588 35252 36318
rect 35980 36372 36036 36382
rect 35980 36278 36036 36316
rect 35308 35588 35364 35598
rect 35196 35586 35364 35588
rect 35196 35534 35310 35586
rect 35362 35534 35364 35586
rect 35196 35532 35364 35534
rect 33846 35308 34110 35318
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 33846 35242 34110 35252
rect 33846 33740 34110 33750
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 33846 33674 34110 33684
rect 33846 32172 34110 32182
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 33846 32106 34110 32116
rect 32508 31892 33124 31948
rect 32956 31220 33012 31230
rect 32396 30100 32452 30110
rect 32396 23378 32452 30044
rect 32396 23326 32398 23378
rect 32450 23326 32452 23378
rect 32396 23314 32452 23326
rect 32508 22820 32564 22830
rect 32508 22594 32564 22764
rect 32508 22542 32510 22594
rect 32562 22542 32564 22594
rect 32508 22530 32564 22542
rect 32284 22372 32340 22382
rect 32284 22278 32340 22316
rect 32060 22204 32228 22260
rect 32060 21364 32116 22204
rect 32844 22148 32900 22158
rect 32172 22146 32900 22148
rect 32172 22094 32846 22146
rect 32898 22094 32900 22146
rect 32172 22092 32900 22094
rect 32172 21586 32228 22092
rect 32844 22082 32900 22092
rect 32396 21924 32452 21934
rect 32172 21534 32174 21586
rect 32226 21534 32228 21586
rect 32172 21522 32228 21534
rect 32284 21868 32396 21924
rect 32284 21364 32340 21868
rect 32396 21858 32452 21868
rect 32396 21700 32452 21710
rect 32956 21700 33012 31164
rect 33068 26516 33124 31892
rect 33846 30604 34110 30614
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 33846 30538 34110 30548
rect 33846 29036 34110 29046
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 33846 28970 34110 28980
rect 33846 27468 34110 27478
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 33846 27402 34110 27412
rect 33068 26450 33124 26460
rect 34188 26068 34244 35532
rect 35308 35476 35364 35532
rect 35308 35410 35364 35420
rect 35756 35588 35812 35598
rect 36204 35588 36260 36430
rect 36652 36370 36708 36652
rect 36876 36484 36932 36494
rect 36652 36318 36654 36370
rect 36706 36318 36708 36370
rect 36652 36306 36708 36318
rect 36764 36482 36932 36484
rect 36764 36430 36878 36482
rect 36930 36430 36932 36482
rect 36764 36428 36932 36430
rect 35756 35586 36260 35588
rect 35756 35534 35758 35586
rect 35810 35534 36260 35586
rect 35756 35532 36260 35534
rect 36316 35588 36372 35598
rect 36764 35588 36820 36428
rect 36876 36418 36932 36428
rect 37324 36370 37380 36876
rect 37548 36484 37604 36494
rect 37324 36318 37326 36370
rect 37378 36318 37380 36370
rect 37324 36306 37380 36318
rect 37436 36482 37604 36484
rect 37436 36430 37550 36482
rect 37602 36430 37604 36482
rect 37436 36428 37604 36430
rect 37212 35698 37268 35710
rect 37212 35646 37214 35698
rect 37266 35646 37268 35698
rect 36316 35586 36820 35588
rect 36316 35534 36318 35586
rect 36370 35534 36820 35586
rect 36316 35532 36820 35534
rect 36876 35588 36932 35598
rect 37212 35588 37268 35646
rect 36876 35586 37268 35588
rect 36876 35534 36878 35586
rect 36930 35534 37268 35586
rect 36876 35532 37268 35534
rect 34412 35364 34468 35374
rect 34412 30324 34468 35308
rect 34412 30258 34468 30268
rect 35756 27300 35812 35532
rect 35756 27234 35812 27244
rect 36092 34020 36148 34030
rect 34188 26002 34244 26012
rect 35308 26964 35364 26974
rect 33846 25900 34110 25910
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 33846 25834 34110 25844
rect 35308 24836 35364 26908
rect 35308 24770 35364 24780
rect 33846 24332 34110 24342
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 33846 24266 34110 24276
rect 35308 23828 35364 23838
rect 33846 22764 34110 22774
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 33846 22698 34110 22708
rect 35308 22484 35364 23772
rect 35308 22418 35364 22428
rect 32396 21698 33012 21700
rect 32396 21646 32398 21698
rect 32450 21646 33012 21698
rect 32396 21644 33012 21646
rect 32396 21634 32452 21644
rect 32060 21298 32116 21308
rect 32172 21308 32340 21364
rect 31612 20850 31668 20860
rect 30716 20804 30772 20814
rect 30716 20710 30772 20748
rect 31164 20802 31220 20814
rect 32060 20804 32116 20814
rect 31164 20750 31166 20802
rect 31218 20750 31220 20802
rect 31164 20580 31220 20750
rect 31836 20802 32116 20804
rect 31836 20750 32062 20802
rect 32114 20750 32116 20802
rect 31836 20748 32116 20750
rect 31724 20692 31780 20702
rect 31724 20598 31780 20636
rect 31164 20514 31220 20524
rect 31836 20580 31892 20748
rect 32060 20738 32116 20748
rect 31836 20514 31892 20524
rect 29932 20132 30212 20188
rect 29820 20078 29822 20130
rect 29874 20078 29876 20130
rect 29820 20066 29876 20078
rect 30156 20130 30212 20132
rect 30156 20078 30158 20130
rect 30210 20078 30212 20130
rect 30156 20066 30212 20078
rect 32172 20130 32228 21308
rect 33846 21196 34110 21206
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 33846 21130 34110 21140
rect 32284 20916 32340 20926
rect 32284 20822 32340 20860
rect 32956 20692 33012 20702
rect 32956 20598 33012 20636
rect 33292 20692 33348 20702
rect 33292 20598 33348 20636
rect 36092 20692 36148 33964
rect 36316 24612 36372 35532
rect 36316 24546 36372 24556
rect 36876 23268 36932 35532
rect 37100 34692 37156 34702
rect 37436 34692 37492 36428
rect 37548 36418 37604 36428
rect 38108 36258 38164 36270
rect 38108 36206 38110 36258
rect 38162 36206 38164 36258
rect 37548 35810 37604 35822
rect 37548 35758 37550 35810
rect 37602 35758 37604 35810
rect 37548 35700 37604 35758
rect 37548 35634 37604 35644
rect 37884 35700 37940 35710
rect 38108 35700 38164 36206
rect 38508 36092 38772 36102
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38508 36026 38772 36036
rect 37884 35698 38164 35700
rect 37884 35646 37886 35698
rect 37938 35646 38164 35698
rect 37884 35644 38164 35646
rect 38220 35810 38276 35822
rect 38220 35758 38222 35810
rect 38274 35758 38276 35810
rect 37884 35364 37940 35644
rect 37884 35298 37940 35308
rect 38220 35028 38276 35758
rect 38220 34962 38276 34972
rect 37660 34804 37716 34814
rect 37884 34804 37940 34814
rect 37716 34802 37940 34804
rect 37716 34750 37886 34802
rect 37938 34750 37940 34802
rect 37716 34748 37940 34750
rect 37660 34710 37716 34748
rect 37884 34738 37940 34748
rect 37100 34690 37492 34692
rect 37100 34638 37102 34690
rect 37154 34638 37492 34690
rect 37100 34636 37492 34638
rect 38220 34692 38276 34702
rect 38220 34690 38388 34692
rect 38220 34638 38222 34690
rect 38274 34638 38388 34690
rect 38220 34636 38388 34638
rect 37100 30436 37156 34636
rect 38220 34626 38276 34636
rect 38332 34356 38388 34636
rect 38508 34524 38772 34534
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38508 34458 38772 34468
rect 38444 34356 38500 34366
rect 38332 34300 38444 34356
rect 38444 34290 38500 34300
rect 38220 34242 38276 34254
rect 38220 34190 38222 34242
rect 38274 34190 38276 34242
rect 37996 34130 38052 34142
rect 37996 34078 37998 34130
rect 38050 34078 38052 34130
rect 37548 34020 37604 34030
rect 37548 33926 37604 33964
rect 37996 34020 38052 34078
rect 37996 33954 38052 33964
rect 38220 33684 38276 34190
rect 38220 33618 38276 33628
rect 37884 33234 37940 33246
rect 37884 33182 37886 33234
rect 37938 33182 37940 33234
rect 37660 33124 37716 33134
rect 37884 33124 37940 33182
rect 37716 33068 37940 33124
rect 38220 33124 38276 33134
rect 37660 33030 37716 33068
rect 38220 33030 38276 33068
rect 38508 32956 38772 32966
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38508 32890 38772 32900
rect 38220 32674 38276 32686
rect 38220 32622 38222 32674
rect 38274 32622 38276 32674
rect 37548 32564 37604 32574
rect 37548 32470 37604 32508
rect 37996 32564 38052 32574
rect 37996 32470 38052 32508
rect 38220 32340 38276 32622
rect 38220 32274 38276 32284
rect 37212 31668 37268 31678
rect 37212 31574 37268 31612
rect 37548 31668 37604 31678
rect 37548 31574 37604 31612
rect 37884 31666 37940 31678
rect 37884 31614 37886 31666
rect 37938 31614 37940 31666
rect 37884 31220 37940 31614
rect 38220 31556 38276 31566
rect 38220 31554 38388 31556
rect 38220 31502 38222 31554
rect 38274 31502 38388 31554
rect 38220 31500 38388 31502
rect 38220 31490 38276 31500
rect 37884 31154 37940 31164
rect 38220 31106 38276 31118
rect 38220 31054 38222 31106
rect 38274 31054 38276 31106
rect 37884 30996 37940 31006
rect 37884 30902 37940 30940
rect 37100 30370 37156 30380
rect 38220 30324 38276 31054
rect 38332 30996 38388 31500
rect 38508 31388 38772 31398
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38508 31322 38772 31332
rect 38444 30996 38500 31006
rect 38332 30940 38444 30996
rect 38444 30930 38500 30940
rect 38220 30258 38276 30268
rect 37884 30100 37940 30110
rect 37884 30006 37940 30044
rect 38220 29986 38276 29998
rect 38220 29934 38222 29986
rect 38274 29934 38276 29986
rect 38220 29764 38276 29934
rect 38508 29820 38772 29830
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38508 29754 38772 29764
rect 38220 29698 38276 29708
rect 38220 29538 38276 29550
rect 38220 29486 38222 29538
rect 38274 29486 38276 29538
rect 37884 29428 37940 29438
rect 37884 29334 37940 29372
rect 38220 28980 38276 29486
rect 38220 28914 38276 28924
rect 37884 28532 37940 28542
rect 37660 28530 37940 28532
rect 37660 28478 37886 28530
rect 37938 28478 37940 28530
rect 37660 28476 37940 28478
rect 37548 27748 37604 27758
rect 37548 27654 37604 27692
rect 37212 27188 37268 27198
rect 37212 27074 37268 27132
rect 37212 27022 37214 27074
rect 37266 27022 37268 27074
rect 37212 27010 37268 27022
rect 37548 27076 37604 27086
rect 37548 26962 37604 27020
rect 37548 26910 37550 26962
rect 37602 26910 37604 26962
rect 37548 26898 37604 26910
rect 37660 25396 37716 28476
rect 37884 28466 37940 28476
rect 38220 28420 38276 28430
rect 38220 28326 38276 28364
rect 38508 28252 38772 28262
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38508 28186 38772 28196
rect 38220 27970 38276 27982
rect 38220 27918 38222 27970
rect 38274 27918 38276 27970
rect 37996 27858 38052 27870
rect 37996 27806 37998 27858
rect 38050 27806 38052 27858
rect 37996 27748 38052 27806
rect 37996 27682 38052 27692
rect 38220 27636 38276 27918
rect 38220 27570 38276 27580
rect 37884 26964 37940 26974
rect 38220 26964 38276 26974
rect 37884 26870 37940 26908
rect 38108 26962 38276 26964
rect 38108 26910 38222 26962
rect 38274 26910 38276 26962
rect 38108 26908 38276 26910
rect 37884 26292 37940 26302
rect 37660 25330 37716 25340
rect 37772 26290 37940 26292
rect 37772 26238 37886 26290
rect 37938 26238 37940 26290
rect 37772 26236 37940 26238
rect 37772 24164 37828 26236
rect 37884 26226 37940 26236
rect 38108 26292 38164 26908
rect 38220 26898 38276 26908
rect 38508 26684 38772 26694
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38508 26618 38772 26628
rect 38108 26226 38164 26236
rect 38220 26402 38276 26414
rect 38220 26350 38222 26402
rect 38274 26350 38276 26402
rect 38220 25620 38276 26350
rect 38220 25554 38276 25564
rect 37884 25396 37940 25406
rect 37884 25394 38052 25396
rect 37884 25342 37886 25394
rect 37938 25342 38052 25394
rect 37884 25340 38052 25342
rect 37884 25330 37940 25340
rect 37884 24724 37940 24734
rect 37884 24630 37940 24668
rect 37772 24098 37828 24108
rect 37884 23828 37940 23838
rect 37884 23734 37940 23772
rect 36876 23202 36932 23212
rect 37884 23154 37940 23166
rect 37884 23102 37886 23154
rect 37938 23102 37940 23154
rect 37884 22596 37940 23102
rect 37884 22530 37940 22540
rect 37212 22258 37268 22270
rect 37884 22260 37940 22270
rect 37212 22206 37214 22258
rect 37266 22206 37268 22258
rect 37212 21028 37268 22206
rect 37772 22258 37940 22260
rect 37772 22206 37886 22258
rect 37938 22206 37940 22258
rect 37772 22204 37940 22206
rect 37548 22146 37604 22158
rect 37548 22094 37550 22146
rect 37602 22094 37604 22146
rect 37548 21588 37604 22094
rect 37772 21812 37828 22204
rect 37884 22194 37940 22204
rect 37996 21924 38052 25340
rect 38220 25284 38276 25294
rect 38220 25190 38276 25228
rect 38508 25116 38772 25126
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38508 25050 38772 25060
rect 38220 24834 38276 24846
rect 38220 24782 38222 24834
rect 38274 24782 38276 24834
rect 38220 24276 38276 24782
rect 38220 24210 38276 24220
rect 38220 23716 38276 23726
rect 38220 23622 38276 23660
rect 38508 23548 38772 23558
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38508 23482 38772 23492
rect 38220 23266 38276 23278
rect 38220 23214 38222 23266
rect 38274 23214 38276 23266
rect 38220 22932 38276 23214
rect 38220 22866 38276 22876
rect 38220 22260 38276 22270
rect 38220 22166 38276 22204
rect 38508 21980 38772 21990
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38508 21914 38772 21924
rect 37996 21858 38052 21868
rect 37772 21746 37828 21756
rect 37884 21700 37940 21710
rect 37884 21606 37940 21644
rect 38220 21698 38276 21710
rect 38220 21646 38222 21698
rect 38274 21646 38276 21698
rect 37548 21522 37604 21532
rect 37212 20962 37268 20972
rect 38220 20916 38276 21646
rect 38220 20850 38276 20860
rect 37884 20804 37940 20814
rect 37884 20710 37940 20748
rect 36092 20626 36148 20636
rect 32172 20078 32174 20130
rect 32226 20078 32228 20130
rect 32172 20066 32228 20078
rect 32620 20578 32676 20590
rect 32620 20526 32622 20578
rect 32674 20526 32676 20578
rect 29036 19954 29092 19964
rect 31948 20018 32004 20030
rect 31948 19966 31950 20018
rect 32002 19966 32004 20018
rect 31948 19908 32004 19966
rect 32620 19908 32676 20526
rect 38220 20580 38276 20590
rect 38220 20578 38388 20580
rect 38220 20526 38222 20578
rect 38274 20526 38388 20578
rect 38220 20524 38388 20526
rect 38220 20514 38276 20524
rect 38332 20244 38388 20524
rect 38508 20412 38772 20422
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38508 20346 38772 20356
rect 38444 20244 38500 20254
rect 38332 20188 38444 20244
rect 38444 20178 38500 20188
rect 31948 19852 32676 19908
rect 36540 20132 36596 20142
rect 33846 19628 34110 19638
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 33846 19562 34110 19572
rect 32956 19460 33012 19470
rect 29596 19236 29652 19246
rect 29148 19124 29204 19134
rect 29148 19030 29204 19068
rect 29484 19012 29540 19050
rect 29484 18946 29540 18956
rect 29184 18844 29448 18854
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29184 18778 29448 18788
rect 29596 18452 29652 19180
rect 30380 19236 30436 19246
rect 30380 19234 30548 19236
rect 30380 19182 30382 19234
rect 30434 19182 30548 19234
rect 30380 19180 30548 19182
rect 30380 19170 30436 19180
rect 29596 18358 29652 18396
rect 30156 19124 30212 19134
rect 30156 18450 30212 19068
rect 30492 18674 30548 19180
rect 31948 19234 32004 19246
rect 31948 19182 31950 19234
rect 32002 19182 32004 19234
rect 30940 19124 30996 19134
rect 30940 19030 30996 19068
rect 30492 18622 30494 18674
rect 30546 18622 30548 18674
rect 30492 18610 30548 18622
rect 30604 19010 30660 19022
rect 30604 18958 30606 19010
rect 30658 18958 30660 19010
rect 30156 18398 30158 18450
rect 30210 18398 30212 18450
rect 30156 18386 30212 18398
rect 29820 18228 29876 18238
rect 29708 18172 29820 18228
rect 29708 17668 29764 18172
rect 29820 18134 29876 18172
rect 29484 17612 29876 17668
rect 29148 17556 29204 17566
rect 29036 17554 29204 17556
rect 29036 17502 29150 17554
rect 29202 17502 29204 17554
rect 29036 17500 29204 17502
rect 28924 17220 28980 17230
rect 29036 17220 29092 17500
rect 29148 17490 29204 17500
rect 29484 17554 29540 17612
rect 29484 17502 29486 17554
rect 29538 17502 29540 17554
rect 29484 17490 29540 17502
rect 28980 17164 29092 17220
rect 29184 17276 29448 17286
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29184 17210 29448 17220
rect 28924 17154 28980 17164
rect 29148 16994 29204 17006
rect 29148 16942 29150 16994
rect 29202 16942 29204 16994
rect 28924 16884 28980 16894
rect 28700 16882 28980 16884
rect 28700 16830 28926 16882
rect 28978 16830 28980 16882
rect 28700 16828 28980 16830
rect 28364 15810 28420 15820
rect 27020 15596 27412 15652
rect 26348 15374 26350 15426
rect 26402 15374 26404 15426
rect 26348 15362 26404 15374
rect 26572 15428 26628 15438
rect 26012 13346 26068 13356
rect 26460 15314 26516 15326
rect 26460 15262 26462 15314
rect 26514 15262 26516 15314
rect 26460 13076 26516 15262
rect 26572 15314 26628 15372
rect 26572 15262 26574 15314
rect 26626 15262 26628 15314
rect 26572 15148 26628 15262
rect 27356 15314 27412 15596
rect 28812 15540 28868 15550
rect 28812 15446 28868 15484
rect 27356 15262 27358 15314
rect 27410 15262 27412 15314
rect 26572 15092 26852 15148
rect 26572 14532 26628 14542
rect 26572 13748 26628 14476
rect 26796 13858 26852 15092
rect 27020 15090 27076 15102
rect 27020 15038 27022 15090
rect 27074 15038 27076 15090
rect 27020 14530 27076 15038
rect 27020 14478 27022 14530
rect 27074 14478 27076 14530
rect 27020 14466 27076 14478
rect 27356 14532 27412 15262
rect 27580 15314 27636 15326
rect 27580 15262 27582 15314
rect 27634 15262 27636 15314
rect 27580 15204 27636 15262
rect 27580 15138 27636 15148
rect 27692 15314 27748 15326
rect 27692 15262 27694 15314
rect 27746 15262 27748 15314
rect 27356 14466 27412 14476
rect 27244 14306 27300 14318
rect 27244 14254 27246 14306
rect 27298 14254 27300 14306
rect 27244 13972 27300 14254
rect 27692 13972 27748 15262
rect 28140 15316 28196 15326
rect 28476 15316 28532 15326
rect 28140 15314 28532 15316
rect 28140 15262 28142 15314
rect 28194 15262 28478 15314
rect 28530 15262 28532 15314
rect 28140 15260 28532 15262
rect 28140 15250 28196 15260
rect 28476 15250 28532 15260
rect 28028 14532 28084 14542
rect 27244 13906 27300 13916
rect 27356 13916 27972 13972
rect 26796 13806 26798 13858
rect 26850 13806 26852 13858
rect 26572 13654 26628 13692
rect 26684 13746 26740 13758
rect 26684 13694 26686 13746
rect 26738 13694 26740 13746
rect 26684 13524 26740 13694
rect 26796 13748 26852 13806
rect 27356 13748 27412 13916
rect 27916 13858 27972 13916
rect 27916 13806 27918 13858
rect 27970 13806 27972 13858
rect 27916 13794 27972 13806
rect 26796 13692 27412 13748
rect 27580 13748 27636 13758
rect 27804 13748 27860 13758
rect 27580 13654 27636 13692
rect 27692 13746 27860 13748
rect 27692 13694 27806 13746
rect 27858 13694 27860 13746
rect 27692 13692 27860 13694
rect 26684 13458 26740 13468
rect 27244 13524 27300 13534
rect 27244 13522 27524 13524
rect 27244 13470 27246 13522
rect 27298 13470 27524 13522
rect 27244 13468 27524 13470
rect 27244 13458 27300 13468
rect 26236 13020 26516 13076
rect 26572 13300 26628 13310
rect 25452 12964 25508 12974
rect 25340 12962 25508 12964
rect 25340 12910 25454 12962
rect 25506 12910 25508 12962
rect 25340 12908 25508 12910
rect 25452 12898 25508 12908
rect 25788 12852 25844 12862
rect 25788 12758 25844 12796
rect 26124 12740 26180 12750
rect 25900 12738 26180 12740
rect 25900 12686 26126 12738
rect 26178 12686 26180 12738
rect 25900 12684 26180 12686
rect 25900 12628 25956 12684
rect 26124 12674 26180 12684
rect 25228 12126 25230 12178
rect 25282 12126 25284 12178
rect 25228 11732 25284 12126
rect 25228 11666 25284 11676
rect 25340 12572 25956 12628
rect 25340 11396 25396 12572
rect 26236 12516 26292 13020
rect 26124 12460 26292 12516
rect 26460 12850 26516 12862
rect 26460 12798 26462 12850
rect 26514 12798 26516 12850
rect 25788 12404 25844 12414
rect 25788 12310 25844 12348
rect 25452 12180 25508 12218
rect 25452 12114 25508 12124
rect 26124 12178 26180 12460
rect 26124 12126 26126 12178
rect 26178 12126 26180 12178
rect 25900 11956 25956 11966
rect 25956 11900 26068 11956
rect 25900 11890 25956 11900
rect 25676 11506 25732 11518
rect 25676 11454 25678 11506
rect 25730 11454 25732 11506
rect 24556 11284 24612 11294
rect 24556 11190 24612 11228
rect 24780 11170 24836 11182
rect 24780 11118 24782 11170
rect 24834 11118 24836 11170
rect 24668 10612 24724 10622
rect 24668 10518 24724 10556
rect 24780 10388 24836 11118
rect 23548 9202 23604 9212
rect 23884 10108 24164 10164
rect 24220 10332 24836 10388
rect 23212 9102 23214 9154
rect 23266 9102 23268 9154
rect 23212 8932 23268 9102
rect 23324 9156 23380 9166
rect 23324 9062 23380 9100
rect 23548 9044 23604 9054
rect 23548 8950 23604 8988
rect 23884 9044 23940 10108
rect 23884 8978 23940 8988
rect 23996 9042 24052 9054
rect 23996 8990 23998 9042
rect 24050 8990 24052 9042
rect 23212 8876 23492 8932
rect 22876 8754 22932 8764
rect 22988 8818 23044 8830
rect 22988 8766 22990 8818
rect 23042 8766 23044 8818
rect 22876 8484 22932 8494
rect 22876 8370 22932 8428
rect 22876 8318 22878 8370
rect 22930 8318 22932 8370
rect 22876 8306 22932 8318
rect 22988 8372 23044 8766
rect 22988 8316 23380 8372
rect 23100 8148 23156 8158
rect 23100 8054 23156 8092
rect 22876 8036 22932 8046
rect 22876 7942 22932 7980
rect 22876 7700 22932 7710
rect 22764 7698 22932 7700
rect 22764 7646 22878 7698
rect 22930 7646 22932 7698
rect 22764 7644 22932 7646
rect 22876 7634 22932 7644
rect 22988 7476 23044 7486
rect 22988 7382 23044 7420
rect 22428 3442 22596 3444
rect 22428 3390 22430 3442
rect 22482 3390 22596 3442
rect 22428 3388 22596 3390
rect 22652 3554 22708 3566
rect 22652 3502 22654 3554
rect 22706 3502 22708 3554
rect 22428 3378 22484 3388
rect 22652 2548 22708 3502
rect 23324 3554 23380 8316
rect 23436 7586 23492 8876
rect 23660 8260 23716 8270
rect 23548 8204 23660 8260
rect 23548 7698 23604 8204
rect 23660 8194 23716 8204
rect 23884 8258 23940 8270
rect 23884 8206 23886 8258
rect 23938 8206 23940 8258
rect 23548 7646 23550 7698
rect 23602 7646 23604 7698
rect 23548 7634 23604 7646
rect 23436 7534 23438 7586
rect 23490 7534 23492 7586
rect 23436 7522 23492 7534
rect 23884 7252 23940 8206
rect 23996 8260 24052 8990
rect 24108 9042 24164 9054
rect 24108 8990 24110 9042
rect 24162 8990 24164 9042
rect 24108 8820 24164 8990
rect 24108 8754 24164 8764
rect 24220 8260 24276 10332
rect 24522 10220 24786 10230
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24522 10154 24786 10164
rect 24892 9940 24948 11340
rect 24332 9884 24948 9940
rect 25004 11340 25396 11396
rect 25004 11282 25060 11340
rect 25004 11230 25006 11282
rect 25058 11230 25060 11282
rect 24332 9266 24388 9884
rect 24892 9716 24948 9726
rect 24892 9622 24948 9660
rect 25004 9492 25060 11230
rect 25340 11282 25396 11340
rect 25564 11396 25620 11406
rect 25564 11302 25620 11340
rect 25340 11230 25342 11282
rect 25394 11230 25396 11282
rect 25340 11218 25396 11230
rect 24332 9214 24334 9266
rect 24386 9214 24388 9266
rect 24332 9044 24388 9214
rect 24332 8978 24388 8988
rect 24556 9436 25060 9492
rect 25116 11170 25172 11182
rect 25116 11118 25118 11170
rect 25170 11118 25172 11170
rect 24556 9154 24612 9436
rect 24556 9102 24558 9154
rect 24610 9102 24612 9154
rect 24556 8820 24612 9102
rect 24668 8932 24724 8942
rect 24668 8930 24948 8932
rect 24668 8878 24670 8930
rect 24722 8878 24948 8930
rect 24668 8876 24948 8878
rect 24668 8866 24724 8876
rect 23996 8204 24164 8260
rect 23996 8034 24052 8046
rect 23996 7982 23998 8034
rect 24050 7982 24052 8034
rect 23996 7924 24052 7982
rect 23996 7858 24052 7868
rect 24108 7698 24164 8204
rect 24332 8764 24612 8820
rect 24332 8260 24388 8764
rect 24522 8652 24786 8662
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24522 8586 24786 8596
rect 24668 8372 24724 8382
rect 24444 8260 24500 8270
rect 24332 8258 24500 8260
rect 24332 8206 24446 8258
rect 24498 8206 24500 8258
rect 24332 8204 24500 8206
rect 24220 8166 24276 8204
rect 24444 8194 24500 8204
rect 24668 8148 24724 8316
rect 24780 8260 24836 8270
rect 24780 8166 24836 8204
rect 24556 8036 24612 8046
rect 24556 7942 24612 7980
rect 24108 7646 24110 7698
rect 24162 7646 24164 7698
rect 24108 7634 24164 7646
rect 24220 7588 24276 7598
rect 24668 7588 24724 8092
rect 24220 7586 24724 7588
rect 24220 7534 24222 7586
rect 24274 7534 24670 7586
rect 24722 7534 24724 7586
rect 24220 7532 24724 7534
rect 24220 7522 24276 7532
rect 24668 7522 24724 7532
rect 24556 7252 24612 7262
rect 23884 7250 24612 7252
rect 23884 7198 24558 7250
rect 24610 7198 24612 7250
rect 23884 7196 24612 7198
rect 24556 7186 24612 7196
rect 24522 7084 24786 7094
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24522 7018 24786 7028
rect 24522 5516 24786 5526
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24522 5450 24786 5460
rect 24892 4900 24948 8876
rect 25004 8820 25060 8830
rect 25004 8034 25060 8764
rect 25004 7982 25006 8034
rect 25058 7982 25060 8034
rect 25004 7924 25060 7982
rect 25004 7858 25060 7868
rect 25116 6692 25172 11118
rect 25340 10610 25396 10622
rect 25340 10558 25342 10610
rect 25394 10558 25396 10610
rect 25228 9716 25284 9726
rect 25228 9042 25284 9660
rect 25228 8990 25230 9042
rect 25282 8990 25284 9042
rect 25228 8978 25284 8990
rect 25228 8820 25284 8830
rect 25228 8258 25284 8764
rect 25340 8484 25396 10558
rect 25340 8418 25396 8428
rect 25452 9604 25508 9614
rect 25228 8206 25230 8258
rect 25282 8206 25284 8258
rect 25228 8194 25284 8206
rect 25452 8258 25508 9548
rect 25452 8206 25454 8258
rect 25506 8206 25508 8258
rect 25452 8194 25508 8206
rect 25116 6626 25172 6636
rect 25564 8034 25620 8046
rect 25564 7982 25566 8034
rect 25618 7982 25620 8034
rect 25564 5012 25620 7982
rect 25676 6580 25732 11454
rect 25788 11282 25844 11294
rect 25788 11230 25790 11282
rect 25842 11230 25844 11282
rect 25788 9716 25844 11230
rect 25788 9650 25844 9660
rect 25900 8372 25956 8382
rect 25788 8260 25844 8270
rect 25788 8166 25844 8204
rect 25900 8258 25956 8316
rect 25900 8206 25902 8258
rect 25954 8206 25956 8258
rect 25900 8194 25956 8206
rect 25676 6514 25732 6524
rect 25564 4946 25620 4956
rect 24892 4834 24948 4844
rect 26012 4788 26068 11900
rect 26124 11620 26180 12126
rect 26236 12180 26292 12190
rect 26236 12068 26292 12124
rect 26348 12068 26404 12078
rect 26236 12066 26404 12068
rect 26236 12014 26350 12066
rect 26402 12014 26404 12066
rect 26236 12012 26404 12014
rect 26348 12002 26404 12012
rect 26124 11554 26180 11564
rect 26236 11508 26292 11518
rect 26460 11508 26516 12798
rect 26292 11452 26516 11508
rect 26236 11414 26292 11452
rect 26124 11170 26180 11182
rect 26124 11118 26126 11170
rect 26178 11118 26180 11170
rect 26124 9604 26180 11118
rect 26124 9538 26180 9548
rect 26572 8260 26628 13244
rect 27468 12962 27524 13468
rect 27468 12910 27470 12962
rect 27522 12910 27524 12962
rect 27468 12898 27524 12910
rect 27692 12964 27748 13692
rect 27804 13682 27860 13692
rect 26796 12850 26852 12862
rect 26796 12798 26798 12850
rect 26850 12798 26852 12850
rect 26796 12404 26852 12798
rect 26796 12338 26852 12348
rect 27132 12738 27188 12750
rect 27132 12686 27134 12738
rect 27186 12686 27188 12738
rect 27020 12180 27076 12190
rect 26796 12178 27076 12180
rect 26796 12126 27022 12178
rect 27074 12126 27076 12178
rect 26796 12124 27076 12126
rect 26684 12068 26740 12078
rect 26796 12068 26852 12124
rect 27020 12114 27076 12124
rect 26684 12066 26852 12068
rect 26684 12014 26686 12066
rect 26738 12014 26852 12066
rect 26684 12012 26852 12014
rect 26684 12002 26740 12012
rect 26684 11620 26740 11630
rect 26684 11506 26740 11564
rect 27020 11620 27076 11630
rect 26684 11454 26686 11506
rect 26738 11454 26740 11506
rect 26684 11442 26740 11454
rect 26908 11508 26964 11518
rect 27020 11508 27076 11564
rect 26908 11506 27076 11508
rect 26908 11454 26910 11506
rect 26962 11454 27076 11506
rect 26908 11452 27076 11454
rect 26908 11442 26964 11452
rect 26572 8194 26628 8204
rect 26684 10388 26740 10398
rect 25564 4732 26068 4788
rect 26124 8036 26180 8046
rect 24892 4564 24948 4574
rect 24522 3948 24786 3958
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24522 3882 24786 3892
rect 23324 3502 23326 3554
rect 23378 3502 23380 3554
rect 23324 3490 23380 3502
rect 24220 3556 24276 3566
rect 23100 3332 23156 3342
rect 22204 2492 22708 2548
rect 22876 3330 23156 3332
rect 22876 3278 23102 3330
rect 23154 3278 23156 3330
rect 22876 3276 23156 3278
rect 22204 800 22260 2492
rect 22876 800 22932 3276
rect 23100 3266 23156 3276
rect 23772 1876 23828 1886
rect 23548 1820 23772 1876
rect 23548 800 23604 1820
rect 23772 1810 23828 1820
rect 24220 800 24276 3500
rect 24892 3554 24948 4508
rect 24892 3502 24894 3554
rect 24946 3502 24948 3554
rect 24892 3490 24948 3502
rect 25228 3556 25284 3566
rect 25004 3444 25060 3454
rect 24556 3330 24612 3342
rect 24556 3278 24558 3330
rect 24610 3278 24612 3330
rect 24556 1876 24612 3278
rect 24556 1810 24612 1820
rect 24892 3332 25060 3388
rect 25228 3442 25284 3500
rect 25564 3554 25620 4732
rect 25564 3502 25566 3554
rect 25618 3502 25620 3554
rect 25564 3490 25620 3502
rect 26124 3554 26180 7980
rect 26124 3502 26126 3554
rect 26178 3502 26180 3554
rect 26124 3490 26180 3502
rect 26684 3556 26740 10332
rect 27132 10164 27188 12686
rect 27356 12292 27412 12302
rect 27356 12290 27524 12292
rect 27356 12238 27358 12290
rect 27410 12238 27524 12290
rect 27356 12236 27524 12238
rect 27356 12226 27412 12236
rect 27244 11172 27300 11182
rect 27244 11078 27300 11116
rect 27244 10612 27300 10622
rect 27244 10498 27300 10556
rect 27244 10446 27246 10498
rect 27298 10446 27300 10498
rect 27244 10434 27300 10446
rect 27468 10388 27524 12236
rect 27692 12180 27748 12908
rect 27804 12740 27860 12750
rect 27804 12646 27860 12684
rect 27804 12180 27860 12190
rect 28028 12180 28084 14476
rect 28588 14532 28644 14542
rect 28140 14420 28196 14430
rect 28140 12852 28196 14364
rect 28252 14418 28308 14430
rect 28252 14366 28254 14418
rect 28306 14366 28308 14418
rect 28252 14084 28308 14366
rect 28588 14418 28644 14476
rect 28588 14366 28590 14418
rect 28642 14366 28644 14418
rect 28588 14354 28644 14366
rect 28252 14018 28308 14028
rect 28812 14084 28868 14094
rect 28924 14084 28980 16828
rect 29148 16772 29204 16942
rect 29484 16884 29540 16894
rect 29540 16828 29652 16884
rect 29484 16790 29540 16828
rect 29148 16706 29204 16716
rect 29596 16210 29652 16828
rect 29708 16772 29764 16782
rect 29708 16678 29764 16716
rect 29820 16322 29876 17612
rect 30044 16884 30100 16894
rect 30380 16884 30436 16894
rect 30044 16882 30436 16884
rect 30044 16830 30046 16882
rect 30098 16830 30382 16882
rect 30434 16830 30436 16882
rect 30044 16828 30436 16830
rect 30044 16818 30100 16828
rect 30380 16818 30436 16828
rect 29820 16270 29822 16322
rect 29874 16270 29876 16322
rect 29820 16258 29876 16270
rect 29596 16158 29598 16210
rect 29650 16158 29652 16210
rect 29596 16146 29652 16158
rect 30156 15988 30212 15998
rect 30492 15988 30548 15998
rect 30156 15986 30548 15988
rect 30156 15934 30158 15986
rect 30210 15934 30494 15986
rect 30546 15934 30548 15986
rect 30156 15932 30548 15934
rect 30156 15922 30212 15932
rect 30492 15922 30548 15932
rect 29184 15708 29448 15718
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29184 15642 29448 15652
rect 29148 15204 29204 15214
rect 29148 14642 29204 15148
rect 29148 14590 29150 14642
rect 29202 14590 29204 14642
rect 29148 14578 29204 14590
rect 29372 14532 29428 14542
rect 29372 14438 29428 14476
rect 29708 14420 29764 14430
rect 30044 14420 30100 14430
rect 29708 14418 30100 14420
rect 29708 14366 29710 14418
rect 29762 14366 30046 14418
rect 30098 14366 30100 14418
rect 29708 14364 30100 14366
rect 29708 14354 29764 14364
rect 30044 14354 30100 14364
rect 30380 14306 30436 14318
rect 30380 14254 30382 14306
rect 30434 14254 30436 14306
rect 28868 14028 28980 14084
rect 29184 14140 29448 14150
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29184 14074 29448 14084
rect 28812 14018 28868 14028
rect 29036 13858 29092 13870
rect 29036 13806 29038 13858
rect 29090 13806 29092 13858
rect 28364 13748 28420 13758
rect 28700 13748 28756 13758
rect 28364 13746 28756 13748
rect 28364 13694 28366 13746
rect 28418 13694 28702 13746
rect 28754 13694 28756 13746
rect 28364 13692 28756 13694
rect 28364 13682 28420 13692
rect 28700 13682 28756 13692
rect 29036 13524 29092 13806
rect 29036 13458 29092 13468
rect 30044 13636 30100 13646
rect 28140 12786 28196 12796
rect 29184 12572 29448 12582
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29184 12506 29448 12516
rect 29036 12292 29092 12302
rect 29036 12198 29092 12236
rect 27692 12178 27860 12180
rect 27692 12126 27806 12178
rect 27858 12126 27860 12178
rect 27692 12124 27860 12126
rect 27804 12114 27860 12124
rect 27916 12178 28084 12180
rect 27916 12126 28030 12178
rect 28082 12126 28084 12178
rect 27916 12124 28084 12126
rect 27580 11732 27636 11742
rect 27580 11506 27636 11676
rect 27804 11620 27860 11630
rect 27916 11620 27972 12124
rect 28028 12114 28084 12124
rect 28364 12180 28420 12190
rect 28700 12180 28756 12190
rect 28364 12178 28756 12180
rect 28364 12126 28366 12178
rect 28418 12126 28702 12178
rect 28754 12126 28756 12178
rect 28364 12124 28756 12126
rect 28364 12114 28420 12124
rect 28700 12114 28756 12124
rect 27860 11564 27972 11620
rect 27804 11526 27860 11564
rect 27580 11454 27582 11506
rect 27634 11454 27636 11506
rect 27580 11442 27636 11454
rect 28140 11284 28196 11294
rect 28140 11190 28196 11228
rect 29148 11284 29204 11294
rect 29148 11190 29204 11228
rect 27804 11172 27860 11182
rect 29484 11172 29540 11182
rect 30044 11172 30100 13580
rect 30380 13076 30436 14254
rect 30380 13010 30436 13020
rect 27860 11116 28084 11172
rect 27804 11106 27860 11116
rect 27132 10098 27188 10108
rect 27356 10332 27524 10388
rect 26796 9826 26852 9838
rect 26796 9774 26798 9826
rect 26850 9774 26852 9826
rect 26796 8036 26852 9774
rect 27244 9604 27300 9614
rect 27244 9510 27300 9548
rect 27244 8930 27300 8942
rect 27244 8878 27246 8930
rect 27298 8878 27300 8930
rect 27244 8372 27300 8878
rect 27244 8306 27300 8316
rect 26796 7970 26852 7980
rect 27132 8036 27188 8046
rect 27132 7942 27188 7980
rect 27132 4452 27188 4462
rect 26908 4450 27188 4452
rect 26908 4398 27134 4450
rect 27186 4398 27188 4450
rect 26908 4396 27188 4398
rect 26796 3556 26852 3566
rect 26684 3554 26852 3556
rect 26684 3502 26798 3554
rect 26850 3502 26852 3554
rect 26684 3500 26852 3502
rect 26796 3490 26852 3500
rect 25228 3390 25230 3442
rect 25282 3390 25284 3442
rect 25228 3378 25284 3390
rect 25900 3444 25956 3482
rect 26460 3444 26516 3454
rect 25900 3378 25956 3388
rect 26236 3332 26516 3388
rect 24892 800 24948 3332
rect 25564 980 25620 990
rect 25564 800 25620 924
rect 26236 800 26292 3332
rect 26572 3330 26628 3342
rect 26572 3278 26574 3330
rect 26626 3278 26628 3330
rect 26572 980 26628 3278
rect 26572 914 26628 924
rect 26908 800 26964 4396
rect 27132 4386 27188 4396
rect 27356 4338 27412 10332
rect 27580 9938 27636 9950
rect 27580 9886 27582 9938
rect 27634 9886 27636 9938
rect 27468 9602 27524 9614
rect 27468 9550 27470 9602
rect 27522 9550 27524 9602
rect 27468 9268 27524 9550
rect 27468 9202 27524 9212
rect 27580 6804 27636 9886
rect 27804 9826 27860 9838
rect 27804 9774 27806 9826
rect 27858 9774 27860 9826
rect 27804 9716 27860 9774
rect 28028 9826 28084 11116
rect 29484 11170 29652 11172
rect 29484 11118 29486 11170
rect 29538 11118 29652 11170
rect 29484 11116 29652 11118
rect 29484 11106 29540 11116
rect 29184 11004 29448 11014
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29184 10938 29448 10948
rect 28028 9774 28030 9826
rect 28082 9774 28084 9826
rect 28028 9762 28084 9774
rect 29148 10612 29204 10622
rect 29148 9826 29204 10556
rect 29148 9774 29150 9826
rect 29202 9774 29204 9826
rect 29148 9762 29204 9774
rect 27804 9650 27860 9660
rect 28364 9602 28420 9614
rect 28364 9550 28366 9602
rect 28418 9550 28420 9602
rect 28364 8428 28420 9550
rect 29184 9436 29448 9446
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29184 9370 29448 9380
rect 28364 8372 28644 8428
rect 27580 6738 27636 6748
rect 27356 4286 27358 4338
rect 27410 4286 27412 4338
rect 27356 4274 27412 4286
rect 27468 4900 27524 4910
rect 27468 3554 27524 4844
rect 27468 3502 27470 3554
rect 27522 3502 27524 3554
rect 27468 3490 27524 3502
rect 28588 3554 28644 8372
rect 29184 7868 29448 7878
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29184 7802 29448 7812
rect 29184 6300 29448 6310
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29184 6234 29448 6244
rect 29184 4732 29448 4742
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29184 4666 29448 4676
rect 29596 4564 29652 11116
rect 30044 11106 30100 11116
rect 30604 9268 30660 18958
rect 31276 19012 31332 19022
rect 31276 18918 31332 18956
rect 31948 18674 32004 19182
rect 32172 19012 32228 19022
rect 32172 19010 32340 19012
rect 32172 18958 32174 19010
rect 32226 18958 32340 19010
rect 32172 18956 32340 18958
rect 32172 18946 32228 18956
rect 31948 18622 31950 18674
rect 32002 18622 32004 18674
rect 31948 18610 32004 18622
rect 31052 18452 31108 18462
rect 31052 18358 31108 18396
rect 31388 18340 31444 18350
rect 30828 18226 30884 18238
rect 30828 18174 30830 18226
rect 30882 18174 30884 18226
rect 30716 16994 30772 17006
rect 30716 16942 30718 16994
rect 30770 16942 30772 16994
rect 30716 9828 30772 16942
rect 30828 16772 30884 18174
rect 31388 18004 31444 18284
rect 31164 17948 31444 18004
rect 31612 18228 31668 18238
rect 31164 17666 31220 17948
rect 31164 17614 31166 17666
rect 31218 17614 31220 17666
rect 31164 17602 31220 17614
rect 31388 17668 31444 17678
rect 31388 17666 31556 17668
rect 31388 17614 31390 17666
rect 31442 17614 31556 17666
rect 31388 17612 31556 17614
rect 31388 17602 31444 17612
rect 30828 16706 30884 16716
rect 31276 17444 31332 17454
rect 31276 16882 31332 17388
rect 31276 16830 31278 16882
rect 31330 16830 31332 16882
rect 30828 16212 30884 16222
rect 30828 15986 30884 16156
rect 31276 16210 31332 16830
rect 31500 16772 31556 17612
rect 31500 16678 31556 16716
rect 31500 16324 31556 16334
rect 31612 16324 31668 18172
rect 31724 17556 31780 17566
rect 32060 17556 32116 17566
rect 31724 17554 32116 17556
rect 31724 17502 31726 17554
rect 31778 17502 32062 17554
rect 32114 17502 32116 17554
rect 31724 17500 32116 17502
rect 31724 17490 31780 17500
rect 32060 17490 32116 17500
rect 31836 16884 31892 16894
rect 32172 16884 32228 16894
rect 31836 16882 32228 16884
rect 31836 16830 31838 16882
rect 31890 16830 32174 16882
rect 32226 16830 32228 16882
rect 31836 16828 32228 16830
rect 31836 16818 31892 16828
rect 32172 16818 32228 16828
rect 31500 16322 31668 16324
rect 31500 16270 31502 16322
rect 31554 16270 31668 16322
rect 31500 16268 31668 16270
rect 31500 16258 31556 16268
rect 31276 16158 31278 16210
rect 31330 16158 31332 16210
rect 31276 16146 31332 16158
rect 30828 15934 30830 15986
rect 30882 15934 30884 15986
rect 30828 15922 30884 15934
rect 31836 15988 31892 15998
rect 32172 15988 32228 15998
rect 31836 15986 32228 15988
rect 31836 15934 31838 15986
rect 31890 15934 32174 15986
rect 32226 15934 32228 15986
rect 31836 15932 32228 15934
rect 31836 15922 31892 15932
rect 32172 15922 32228 15932
rect 30716 9762 30772 9772
rect 31276 11172 31332 11182
rect 31164 9716 31220 9726
rect 31164 9622 31220 9660
rect 30604 9202 30660 9212
rect 28588 3502 28590 3554
rect 28642 3502 28644 3554
rect 28588 3490 28644 3502
rect 29372 4508 29652 4564
rect 29932 6692 29988 6702
rect 29372 3554 29428 4508
rect 29372 3502 29374 3554
rect 29426 3502 29428 3554
rect 29372 3490 29428 3502
rect 29932 3554 29988 6636
rect 29932 3502 29934 3554
rect 29986 3502 29988 3554
rect 29932 3490 29988 3502
rect 30604 5012 30660 5022
rect 30604 3554 30660 4956
rect 30604 3502 30606 3554
rect 30658 3502 30660 3554
rect 30604 3490 30660 3502
rect 31276 3554 31332 11116
rect 32284 7588 32340 18956
rect 32396 18452 32452 18462
rect 32396 17554 32452 18396
rect 32396 17502 32398 17554
rect 32450 17502 32452 17554
rect 32396 17490 32452 17502
rect 32508 16994 32564 17006
rect 32508 16942 32510 16994
rect 32562 16942 32564 16994
rect 32508 16100 32564 16942
rect 32508 16044 32676 16100
rect 32508 15874 32564 15886
rect 32508 15822 32510 15874
rect 32562 15822 32564 15874
rect 32508 13636 32564 15822
rect 32508 13570 32564 13580
rect 32620 12740 32676 16044
rect 32620 12674 32676 12684
rect 32284 7522 32340 7532
rect 31276 3502 31278 3554
rect 31330 3502 31332 3554
rect 31276 3490 31332 3502
rect 32396 6580 32452 6590
rect 32396 3554 32452 6524
rect 32956 6132 33012 19404
rect 36092 18676 36148 18686
rect 34860 18116 34916 18126
rect 33846 18060 34110 18070
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 33846 17994 34110 18004
rect 33846 16492 34110 16502
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 33846 16426 34110 16436
rect 33516 15876 33572 15886
rect 33516 10724 33572 15820
rect 33846 14924 34110 14934
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 33846 14858 34110 14868
rect 33846 13356 34110 13366
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 33846 13290 34110 13300
rect 34524 12740 34580 12750
rect 33846 11788 34110 11798
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 33846 11722 34110 11732
rect 33516 10658 33572 10668
rect 33846 10220 34110 10230
rect 32956 6066 33012 6076
rect 33068 10164 33124 10174
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 33846 10154 34110 10164
rect 32396 3502 32398 3554
rect 32450 3502 32452 3554
rect 32396 3490 32452 3502
rect 27244 3444 27300 3454
rect 27244 3350 27300 3388
rect 28252 3444 28308 3454
rect 27580 980 27636 990
rect 27580 800 27636 924
rect 28252 800 28308 3388
rect 29036 3444 29092 3454
rect 30380 3444 30436 3454
rect 29036 3350 29092 3388
rect 30044 3442 30436 3444
rect 30044 3390 30382 3442
rect 30434 3390 30436 3442
rect 30044 3388 30436 3390
rect 28364 3330 28420 3342
rect 28364 3278 28366 3330
rect 28418 3278 28420 3330
rect 28364 980 28420 3278
rect 29708 3330 29764 3342
rect 29708 3278 29710 3330
rect 29762 3278 29764 3330
rect 29184 3164 29448 3174
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29184 3098 29448 3108
rect 29708 1316 29764 3278
rect 28364 914 28420 924
rect 28924 1260 29764 1316
rect 28924 800 28980 1260
rect 30044 1092 30100 3388
rect 30380 3378 30436 3388
rect 30940 3444 30996 3454
rect 29596 1036 30100 1092
rect 29596 800 29652 1036
rect 30268 978 30324 990
rect 30268 926 30270 978
rect 30322 926 30324 978
rect 30268 800 30324 926
rect 30940 800 30996 3388
rect 32172 3444 32228 3454
rect 32172 3350 32228 3388
rect 32844 3442 32900 3454
rect 32844 3390 32846 3442
rect 32898 3390 32900 3442
rect 31052 3330 31108 3342
rect 31836 3332 31892 3342
rect 31052 3278 31054 3330
rect 31106 3278 31108 3330
rect 31052 978 31108 3278
rect 31052 926 31054 978
rect 31106 926 31108 978
rect 31052 914 31108 926
rect 31612 3276 31836 3332
rect 31612 800 31668 3276
rect 31836 3266 31892 3276
rect 32844 3332 32900 3390
rect 32844 3266 32900 3276
rect 32956 3444 33012 3454
rect 33068 3444 33124 10108
rect 33846 8652 34110 8662
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 33846 8586 34110 8596
rect 34524 8372 34580 12684
rect 34524 8306 34580 8316
rect 34524 8036 34580 8046
rect 33846 7084 34110 7094
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 33846 7018 34110 7028
rect 33628 6804 33684 6814
rect 33404 5908 33460 5918
rect 33404 4564 33460 5852
rect 33404 4498 33460 4508
rect 33628 3556 33684 6748
rect 33846 5516 34110 5526
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 33846 5450 34110 5460
rect 33852 4564 33908 4574
rect 33852 4470 33908 4508
rect 34412 4564 34468 4574
rect 33846 3948 34110 3958
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 33846 3882 34110 3892
rect 33740 3556 33796 3566
rect 33628 3554 33796 3556
rect 33628 3502 33742 3554
rect 33794 3502 33796 3554
rect 33628 3500 33796 3502
rect 33740 3490 33796 3500
rect 34412 3554 34468 4508
rect 34412 3502 34414 3554
rect 34466 3502 34468 3554
rect 34412 3490 34468 3502
rect 33180 3444 33236 3454
rect 33068 3442 33236 3444
rect 33068 3390 33182 3442
rect 33234 3390 33236 3442
rect 33068 3388 33236 3390
rect 32508 1988 32564 1998
rect 32284 1932 32508 1988
rect 32284 800 32340 1932
rect 32508 1922 32564 1932
rect 32956 800 33012 3388
rect 33180 3378 33236 3388
rect 34188 3444 34244 3454
rect 34188 3350 34244 3388
rect 33516 3330 33572 3342
rect 34524 3332 34580 7980
rect 33516 3278 33518 3330
rect 33570 3278 33572 3330
rect 33516 1988 33572 3278
rect 34300 3276 34580 3332
rect 34636 4226 34692 4238
rect 34636 4174 34638 4226
rect 34690 4174 34692 4226
rect 33516 1922 33572 1932
rect 33628 2546 33684 2558
rect 33628 2494 33630 2546
rect 33682 2494 33684 2546
rect 33628 800 33684 2494
rect 34300 800 34356 3276
rect 34636 2546 34692 4174
rect 34860 3442 34916 18060
rect 36092 4564 36148 18620
rect 36092 4498 36148 4508
rect 36316 18004 36372 18014
rect 36316 3668 36372 17948
rect 36428 8260 36484 8270
rect 36428 8166 36484 8204
rect 36540 6692 36596 20076
rect 38220 20130 38276 20142
rect 38220 20078 38222 20130
rect 38274 20078 38276 20130
rect 37884 20020 37940 20030
rect 37884 19926 37940 19964
rect 38220 19572 38276 20078
rect 38220 19506 38276 19516
rect 37884 19124 37940 19134
rect 37884 19030 37940 19068
rect 38220 19012 38276 19022
rect 38220 18918 38276 18956
rect 38508 18844 38772 18854
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38508 18778 38772 18788
rect 38220 18562 38276 18574
rect 38220 18510 38222 18562
rect 38274 18510 38276 18562
rect 37884 18452 37940 18462
rect 37884 18358 37940 18396
rect 38220 18228 38276 18510
rect 38220 18162 38276 18172
rect 37212 17668 37268 17678
rect 37212 17574 37268 17612
rect 37884 17554 37940 17566
rect 37884 17502 37886 17554
rect 37938 17502 37940 17554
rect 37548 17442 37604 17454
rect 37548 17390 37550 17442
rect 37602 17390 37604 17442
rect 37548 16884 37604 17390
rect 37884 17108 37940 17502
rect 38220 17556 38276 17566
rect 38220 17462 38276 17500
rect 38508 17276 38772 17286
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38508 17210 38772 17220
rect 37884 17042 37940 17052
rect 38220 16994 38276 17006
rect 38220 16942 38222 16994
rect 38274 16942 38276 16994
rect 37548 16818 37604 16828
rect 37884 16882 37940 16894
rect 37884 16830 37886 16882
rect 37938 16830 37940 16882
rect 37884 16212 37940 16830
rect 37884 16146 37940 16156
rect 38220 16212 38276 16942
rect 38220 16146 38276 16156
rect 37884 15988 37940 15998
rect 37884 15894 37940 15932
rect 38220 15876 38276 15886
rect 38220 15874 38388 15876
rect 38220 15822 38222 15874
rect 38274 15822 38388 15874
rect 38220 15820 38388 15822
rect 38220 15810 38276 15820
rect 38332 15540 38388 15820
rect 38508 15708 38772 15718
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38508 15642 38772 15652
rect 38444 15540 38500 15550
rect 38332 15484 38444 15540
rect 38444 15474 38500 15484
rect 37884 15428 37940 15438
rect 37884 15334 37940 15372
rect 38220 15426 38276 15438
rect 38220 15374 38222 15426
rect 38274 15374 38276 15426
rect 38220 14868 38276 15374
rect 38220 14802 38276 14812
rect 37884 14420 37940 14430
rect 37884 14326 37940 14364
rect 38220 14308 38276 14318
rect 38220 14214 38276 14252
rect 38508 14140 38772 14150
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38508 14074 38772 14084
rect 37660 13972 37716 13982
rect 37212 12850 37268 12862
rect 37212 12798 37214 12850
rect 37266 12798 37268 12850
rect 37212 12292 37268 12798
rect 37212 12226 37268 12236
rect 37548 12738 37604 12750
rect 37548 12686 37550 12738
rect 37602 12686 37604 12738
rect 37548 12180 37604 12686
rect 37660 12292 37716 13916
rect 38220 13858 38276 13870
rect 38220 13806 38222 13858
rect 38274 13806 38276 13858
rect 37884 13748 37940 13758
rect 37772 13746 37940 13748
rect 37772 13694 37886 13746
rect 37938 13694 37940 13746
rect 37772 13692 37940 13694
rect 37772 12964 37828 13692
rect 37884 13682 37940 13692
rect 38108 13636 38164 13646
rect 37772 12898 37828 12908
rect 37884 13524 37940 13534
rect 37884 12962 37940 13468
rect 37884 12910 37886 12962
rect 37938 12910 37940 12962
rect 37884 12898 37940 12910
rect 37996 13076 38052 13086
rect 37884 12292 37940 12302
rect 37660 12290 37940 12292
rect 37660 12238 37886 12290
rect 37938 12238 37940 12290
rect 37660 12236 37940 12238
rect 37884 12226 37940 12236
rect 37548 12114 37604 12124
rect 37996 11394 38052 13020
rect 37996 11342 37998 11394
rect 38050 11342 38052 11394
rect 37996 11330 38052 11342
rect 37884 10724 37940 10734
rect 37884 10630 37940 10668
rect 37884 9828 37940 9838
rect 37884 9734 37940 9772
rect 36540 6626 36596 6636
rect 36764 9268 36820 9278
rect 36764 5236 36820 9212
rect 37996 9044 38052 9054
rect 38108 9044 38164 13580
rect 38220 13524 38276 13806
rect 38220 13458 38276 13468
rect 38220 12852 38276 12862
rect 38220 12758 38276 12796
rect 38508 12572 38772 12582
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38508 12506 38772 12516
rect 38220 12290 38276 12302
rect 38220 12238 38222 12290
rect 38274 12238 38276 12290
rect 38220 11508 38276 12238
rect 38220 11442 38276 11452
rect 38220 11172 38276 11182
rect 38220 11170 38388 11172
rect 38220 11118 38222 11170
rect 38274 11118 38388 11170
rect 38220 11116 38388 11118
rect 38220 11106 38276 11116
rect 38332 10836 38388 11116
rect 38508 11004 38772 11014
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38508 10938 38772 10948
rect 38444 10836 38500 10846
rect 38332 10780 38444 10836
rect 38444 10770 38500 10780
rect 38220 10722 38276 10734
rect 38220 10670 38222 10722
rect 38274 10670 38276 10722
rect 38220 10164 38276 10670
rect 38220 10098 38276 10108
rect 38220 9604 38276 9614
rect 38220 9510 38276 9548
rect 38508 9436 38772 9446
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38508 9370 38772 9380
rect 37996 9042 38164 9044
rect 37996 8990 37998 9042
rect 38050 8990 38164 9042
rect 37996 8988 38164 8990
rect 38220 9154 38276 9166
rect 38220 9102 38222 9154
rect 38274 9102 38276 9154
rect 37996 8978 38052 8988
rect 38220 8820 38276 9102
rect 38220 8754 38276 8764
rect 37884 8372 37940 8382
rect 37212 8260 37268 8270
rect 37212 8166 37268 8204
rect 37884 8258 37940 8316
rect 37884 8206 37886 8258
rect 37938 8206 37940 8258
rect 37884 8194 37940 8206
rect 38220 8148 38276 8158
rect 38220 8054 38276 8092
rect 37548 8034 37604 8046
rect 37548 7982 37550 8034
rect 37602 7982 37604 8034
rect 37548 7476 37604 7982
rect 38508 7868 38772 7878
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38508 7802 38772 7812
rect 37884 7588 37940 7598
rect 37884 7494 37940 7532
rect 38220 7586 38276 7598
rect 38220 7534 38222 7586
rect 38274 7534 38276 7586
rect 37548 7410 37604 7420
rect 38220 6804 38276 7534
rect 38220 6738 38276 6748
rect 37548 6692 37604 6702
rect 37548 6598 37604 6636
rect 37996 6692 38052 6702
rect 37996 6598 38052 6636
rect 38220 6466 38276 6478
rect 38220 6414 38222 6466
rect 38274 6414 38276 6466
rect 38220 6244 38276 6414
rect 38508 6300 38772 6310
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38508 6234 38772 6244
rect 38220 6178 38276 6188
rect 37660 6132 37716 6142
rect 37716 6076 37940 6132
rect 37660 6038 37716 6076
rect 37884 6018 37940 6076
rect 37884 5966 37886 6018
rect 37938 5966 37940 6018
rect 37884 5954 37940 5966
rect 38220 6018 38276 6030
rect 38220 5966 38222 6018
rect 38274 5966 38276 6018
rect 38220 5460 38276 5966
rect 38220 5394 38276 5404
rect 36764 5170 36820 5180
rect 37548 5236 37604 5246
rect 37548 5142 37604 5180
rect 37996 5236 38052 5246
rect 37996 5122 38052 5180
rect 37996 5070 37998 5122
rect 38050 5070 38052 5122
rect 37996 5058 38052 5070
rect 38220 4900 38276 4910
rect 38220 4806 38276 4844
rect 38508 4732 38772 4742
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38508 4666 38772 4676
rect 37660 4564 37716 4574
rect 37716 4508 37940 4564
rect 37660 4470 37716 4508
rect 37884 4450 37940 4508
rect 37884 4398 37886 4450
rect 37938 4398 37940 4450
rect 37884 4386 37940 4398
rect 38220 4450 38276 4462
rect 38220 4398 38222 4450
rect 38274 4398 38276 4450
rect 38220 4116 38276 4398
rect 38220 4050 38276 4060
rect 36316 3602 36372 3612
rect 37548 3668 37604 3678
rect 37548 3574 37604 3612
rect 37996 3668 38052 3678
rect 34860 3390 34862 3442
rect 34914 3390 34916 3442
rect 34860 3378 34916 3390
rect 35084 3554 35140 3566
rect 35084 3502 35086 3554
rect 35138 3502 35140 3554
rect 34636 2494 34638 2546
rect 34690 2494 34692 2546
rect 34636 2482 34692 2494
rect 35084 2546 35140 3502
rect 37996 3554 38052 3612
rect 37996 3502 37998 3554
rect 38050 3502 38052 3554
rect 37996 3490 38052 3502
rect 38220 3444 38276 3454
rect 38220 3350 38276 3388
rect 38508 3164 38772 3174
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38508 3098 38772 3108
rect 35084 2494 35086 2546
rect 35138 2494 35140 2546
rect 35084 2482 35140 2494
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 11424 0 11536 800
rect 12096 0 12208 800
rect 12768 0 12880 800
rect 13440 0 13552 800
rect 14112 0 14224 800
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 22176 0 22288 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
rect 25536 0 25648 800
rect 26208 0 26320 800
rect 26880 0 26992 800
rect 27552 0 27664 800
rect 28224 0 28336 800
rect 28896 0 29008 800
rect 29568 0 29680 800
rect 30240 0 30352 800
rect 30912 0 31024 800
rect 31584 0 31696 800
rect 32256 0 32368 800
rect 32928 0 33040 800
rect 33600 0 33712 800
rect 34272 0 34384 800
<< via2 >>
rect 1708 32956 1764 33012
rect 1708 32284 1764 32340
rect 1708 31554 1764 31556
rect 1708 31502 1710 31554
rect 1710 31502 1762 31554
rect 1762 31502 1764 31554
rect 1708 31500 1764 31502
rect 1708 30268 1764 30324
rect 1708 29986 1764 29988
rect 1708 29934 1710 29986
rect 1710 29934 1762 29986
rect 1762 29934 1764 29986
rect 1708 29932 1764 29934
rect 2492 32956 2548 33012
rect 1932 30828 1988 30884
rect 2380 31666 2436 31668
rect 2380 31614 2382 31666
rect 2382 31614 2434 31666
rect 2434 31614 2436 31666
rect 2380 31612 2436 31614
rect 2492 30882 2548 30884
rect 2492 30830 2494 30882
rect 2494 30830 2546 30882
rect 2546 30830 2548 30882
rect 2492 30828 2548 30830
rect 2716 31500 2772 31556
rect 1708 28924 1764 28980
rect 1708 28418 1764 28420
rect 1708 28366 1710 28418
rect 1710 28366 1762 28418
rect 1762 28366 1764 28418
rect 1708 28364 1764 28366
rect 1708 27580 1764 27636
rect 1820 26236 1876 26292
rect 1708 25564 1764 25620
rect 1708 25004 1764 25060
rect 1708 24220 1764 24276
rect 1708 23714 1764 23716
rect 1708 23662 1710 23714
rect 1710 23662 1762 23714
rect 1762 23662 1764 23714
rect 1708 23660 1764 23662
rect 1708 22876 1764 22932
rect 1708 22258 1764 22260
rect 1708 22206 1710 22258
rect 1710 22206 1762 22258
rect 1762 22206 1764 22258
rect 1708 22204 1764 22206
rect 1708 20860 1764 20916
rect 2044 29260 2100 29316
rect 2492 29314 2548 29316
rect 2492 29262 2494 29314
rect 2494 29262 2546 29314
rect 2546 29262 2548 29314
rect 2492 29260 2548 29262
rect 2044 28530 2100 28532
rect 2044 28478 2046 28530
rect 2046 28478 2098 28530
rect 2098 28478 2100 28530
rect 2044 28476 2100 28478
rect 2044 27858 2100 27860
rect 2044 27806 2046 27858
rect 2046 27806 2098 27858
rect 2098 27806 2100 27858
rect 2044 27804 2100 27806
rect 2380 26962 2436 26964
rect 2380 26910 2382 26962
rect 2382 26910 2434 26962
rect 2434 26910 2436 26962
rect 2380 26908 2436 26910
rect 2044 25564 2100 25620
rect 2044 24834 2100 24836
rect 2044 24782 2046 24834
rect 2046 24782 2098 24834
rect 2098 24782 2100 24834
rect 2044 24780 2100 24782
rect 2268 25228 2324 25284
rect 2156 23660 2212 23716
rect 2044 23324 2100 23380
rect 2044 22258 2100 22260
rect 2044 22206 2046 22258
rect 2046 22206 2098 22258
rect 2098 22206 2100 22258
rect 2044 22204 2100 22206
rect 2156 22092 2212 22148
rect 2380 21756 2436 21812
rect 2716 26962 2772 26964
rect 2716 26910 2718 26962
rect 2718 26910 2770 26962
rect 2770 26910 2772 26962
rect 2716 26908 2772 26910
rect 2828 25116 2884 25172
rect 2716 22428 2772 22484
rect 2604 21756 2660 21812
rect 2044 21586 2100 21588
rect 2044 21534 2046 21586
rect 2046 21534 2098 21586
rect 2098 21534 2100 21586
rect 2044 21532 2100 21534
rect 1932 20636 1988 20692
rect 2044 20300 2100 20356
rect 1708 20188 1764 20244
rect 2044 20130 2100 20132
rect 2044 20078 2046 20130
rect 2046 20078 2098 20130
rect 2098 20078 2100 20130
rect 2044 20076 2100 20078
rect 1708 19516 1764 19572
rect 3276 31554 3332 31556
rect 3276 31502 3278 31554
rect 3278 31502 3330 31554
rect 3330 31502 3332 31554
rect 3276 31500 3332 31502
rect 3612 30044 3668 30100
rect 3052 26124 3108 26180
rect 4060 29260 4116 29316
rect 5874 36874 5930 36876
rect 5874 36822 5876 36874
rect 5876 36822 5928 36874
rect 5928 36822 5930 36874
rect 5874 36820 5930 36822
rect 5978 36874 6034 36876
rect 5978 36822 5980 36874
rect 5980 36822 6032 36874
rect 6032 36822 6034 36874
rect 5978 36820 6034 36822
rect 6082 36874 6138 36876
rect 6082 36822 6084 36874
rect 6084 36822 6136 36874
rect 6136 36822 6138 36874
rect 6082 36820 6138 36822
rect 5874 35306 5930 35308
rect 5874 35254 5876 35306
rect 5876 35254 5928 35306
rect 5928 35254 5930 35306
rect 5874 35252 5930 35254
rect 5978 35306 6034 35308
rect 5978 35254 5980 35306
rect 5980 35254 6032 35306
rect 6032 35254 6034 35306
rect 5978 35252 6034 35254
rect 6082 35306 6138 35308
rect 6082 35254 6084 35306
rect 6084 35254 6136 35306
rect 6136 35254 6138 35306
rect 6082 35252 6138 35254
rect 5874 33738 5930 33740
rect 5874 33686 5876 33738
rect 5876 33686 5928 33738
rect 5928 33686 5930 33738
rect 5874 33684 5930 33686
rect 5978 33738 6034 33740
rect 5978 33686 5980 33738
rect 5980 33686 6032 33738
rect 6032 33686 6034 33738
rect 5978 33684 6034 33686
rect 6082 33738 6138 33740
rect 6082 33686 6084 33738
rect 6084 33686 6136 33738
rect 6136 33686 6138 33738
rect 6082 33684 6138 33686
rect 5874 32170 5930 32172
rect 5874 32118 5876 32170
rect 5876 32118 5928 32170
rect 5928 32118 5930 32170
rect 5874 32116 5930 32118
rect 5978 32170 6034 32172
rect 5978 32118 5980 32170
rect 5980 32118 6032 32170
rect 6032 32118 6034 32170
rect 5978 32116 6034 32118
rect 6082 32170 6138 32172
rect 6082 32118 6084 32170
rect 6084 32118 6136 32170
rect 6136 32118 6138 32170
rect 6082 32116 6138 32118
rect 5874 30602 5930 30604
rect 5874 30550 5876 30602
rect 5876 30550 5928 30602
rect 5928 30550 5930 30602
rect 5874 30548 5930 30550
rect 5978 30602 6034 30604
rect 5978 30550 5980 30602
rect 5980 30550 6032 30602
rect 6032 30550 6034 30602
rect 5978 30548 6034 30550
rect 6082 30602 6138 30604
rect 6082 30550 6084 30602
rect 6084 30550 6136 30602
rect 6136 30550 6138 30602
rect 6082 30548 6138 30550
rect 4284 29260 4340 29316
rect 5874 29034 5930 29036
rect 5874 28982 5876 29034
rect 5876 28982 5928 29034
rect 5928 28982 5930 29034
rect 5874 28980 5930 28982
rect 5978 29034 6034 29036
rect 5978 28982 5980 29034
rect 5980 28982 6032 29034
rect 6032 28982 6034 29034
rect 5978 28980 6034 28982
rect 6082 29034 6138 29036
rect 6082 28982 6084 29034
rect 6084 28982 6136 29034
rect 6136 28982 6138 29034
rect 6082 28980 6138 28982
rect 5874 27466 5930 27468
rect 5874 27414 5876 27466
rect 5876 27414 5928 27466
rect 5928 27414 5930 27466
rect 5874 27412 5930 27414
rect 5978 27466 6034 27468
rect 5978 27414 5980 27466
rect 5980 27414 6032 27466
rect 6032 27414 6034 27466
rect 5978 27412 6034 27414
rect 6082 27466 6138 27468
rect 6082 27414 6084 27466
rect 6084 27414 6136 27466
rect 6136 27414 6138 27466
rect 6082 27412 6138 27414
rect 4172 27020 4228 27076
rect 5874 25898 5930 25900
rect 5874 25846 5876 25898
rect 5876 25846 5928 25898
rect 5928 25846 5930 25898
rect 5874 25844 5930 25846
rect 5978 25898 6034 25900
rect 5978 25846 5980 25898
rect 5980 25846 6032 25898
rect 6032 25846 6034 25898
rect 5978 25844 6034 25846
rect 6082 25898 6138 25900
rect 6082 25846 6084 25898
rect 6084 25846 6136 25898
rect 6136 25846 6138 25898
rect 6082 25844 6138 25846
rect 5068 25116 5124 25172
rect 6636 29484 6692 29540
rect 6748 29372 6804 29428
rect 6860 30828 6916 30884
rect 6524 25116 6580 25172
rect 6748 26908 6804 26964
rect 5874 24330 5930 24332
rect 5874 24278 5876 24330
rect 5876 24278 5928 24330
rect 5928 24278 5930 24330
rect 5874 24276 5930 24278
rect 5978 24330 6034 24332
rect 5978 24278 5980 24330
rect 5980 24278 6032 24330
rect 6032 24278 6034 24330
rect 5978 24276 6034 24278
rect 6082 24330 6138 24332
rect 6082 24278 6084 24330
rect 6084 24278 6136 24330
rect 6136 24278 6138 24330
rect 6082 24276 6138 24278
rect 5068 23212 5124 23268
rect 5874 22762 5930 22764
rect 5874 22710 5876 22762
rect 5876 22710 5928 22762
rect 5928 22710 5930 22762
rect 5874 22708 5930 22710
rect 5978 22762 6034 22764
rect 5978 22710 5980 22762
rect 5980 22710 6032 22762
rect 6032 22710 6034 22762
rect 5978 22708 6034 22710
rect 6082 22762 6138 22764
rect 6082 22710 6084 22762
rect 6084 22710 6136 22762
rect 6136 22710 6138 22762
rect 6082 22708 6138 22710
rect 4060 22540 4116 22596
rect 6748 22316 6804 22372
rect 7868 30156 7924 30212
rect 9996 35810 10052 35812
rect 9996 35758 9998 35810
rect 9998 35758 10050 35810
rect 10050 35758 10052 35810
rect 9996 35756 10052 35758
rect 9772 35532 9828 35588
rect 10536 36090 10592 36092
rect 10536 36038 10538 36090
rect 10538 36038 10590 36090
rect 10590 36038 10592 36090
rect 10536 36036 10592 36038
rect 10640 36090 10696 36092
rect 10640 36038 10642 36090
rect 10642 36038 10694 36090
rect 10694 36038 10696 36090
rect 10640 36036 10696 36038
rect 10744 36090 10800 36092
rect 10744 36038 10746 36090
rect 10746 36038 10798 36090
rect 10798 36038 10800 36090
rect 10744 36036 10800 36038
rect 10444 35586 10500 35588
rect 10444 35534 10446 35586
rect 10446 35534 10498 35586
rect 10498 35534 10500 35586
rect 10444 35532 10500 35534
rect 10536 34522 10592 34524
rect 10536 34470 10538 34522
rect 10538 34470 10590 34522
rect 10590 34470 10592 34522
rect 10536 34468 10592 34470
rect 10640 34522 10696 34524
rect 10640 34470 10642 34522
rect 10642 34470 10694 34522
rect 10694 34470 10696 34522
rect 10640 34468 10696 34470
rect 10744 34522 10800 34524
rect 10744 34470 10746 34522
rect 10746 34470 10798 34522
rect 10798 34470 10800 34522
rect 10744 34468 10800 34470
rect 10332 33740 10388 33796
rect 10536 32954 10592 32956
rect 10536 32902 10538 32954
rect 10538 32902 10590 32954
rect 10590 32902 10592 32954
rect 10536 32900 10592 32902
rect 10640 32954 10696 32956
rect 10640 32902 10642 32954
rect 10642 32902 10694 32954
rect 10694 32902 10696 32954
rect 10640 32900 10696 32902
rect 10744 32954 10800 32956
rect 10744 32902 10746 32954
rect 10746 32902 10798 32954
rect 10798 32902 10800 32954
rect 10744 32900 10800 32902
rect 11676 33628 11732 33684
rect 8428 27916 8484 27972
rect 9324 31500 9380 31556
rect 7084 26460 7140 26516
rect 6860 21644 6916 21700
rect 6972 25116 7028 25172
rect 9212 22258 9268 22260
rect 9212 22206 9214 22258
rect 9214 22206 9266 22258
rect 9266 22206 9268 22258
rect 9212 22204 9268 22206
rect 6972 21420 7028 21476
rect 5874 21194 5930 21196
rect 5874 21142 5876 21194
rect 5876 21142 5928 21194
rect 5928 21142 5930 21194
rect 5874 21140 5930 21142
rect 5978 21194 6034 21196
rect 5978 21142 5980 21194
rect 5980 21142 6032 21194
rect 6032 21142 6034 21194
rect 5978 21140 6034 21142
rect 6082 21194 6138 21196
rect 6082 21142 6084 21194
rect 6084 21142 6136 21194
rect 6136 21142 6138 21194
rect 6082 21140 6138 21142
rect 10536 31386 10592 31388
rect 10536 31334 10538 31386
rect 10538 31334 10590 31386
rect 10590 31334 10592 31386
rect 10536 31332 10592 31334
rect 10640 31386 10696 31388
rect 10640 31334 10642 31386
rect 10642 31334 10694 31386
rect 10694 31334 10696 31386
rect 10640 31332 10696 31334
rect 10744 31386 10800 31388
rect 10744 31334 10746 31386
rect 10746 31334 10798 31386
rect 10798 31334 10800 31386
rect 10744 31332 10800 31334
rect 10108 30044 10164 30100
rect 9436 27804 9492 27860
rect 10536 29818 10592 29820
rect 10536 29766 10538 29818
rect 10538 29766 10590 29818
rect 10590 29766 10592 29818
rect 10536 29764 10592 29766
rect 10640 29818 10696 29820
rect 10640 29766 10642 29818
rect 10642 29766 10694 29818
rect 10694 29766 10696 29818
rect 10640 29764 10696 29766
rect 10744 29818 10800 29820
rect 10744 29766 10746 29818
rect 10746 29766 10798 29818
rect 10798 29766 10800 29818
rect 10744 29764 10800 29766
rect 11564 30156 11620 30212
rect 15198 36874 15254 36876
rect 15198 36822 15200 36874
rect 15200 36822 15252 36874
rect 15252 36822 15254 36874
rect 15198 36820 15254 36822
rect 15302 36874 15358 36876
rect 15302 36822 15304 36874
rect 15304 36822 15356 36874
rect 15356 36822 15358 36874
rect 15302 36820 15358 36822
rect 15406 36874 15462 36876
rect 15406 36822 15408 36874
rect 15408 36822 15460 36874
rect 15460 36822 15462 36874
rect 15406 36820 15462 36822
rect 12236 30044 12292 30100
rect 13692 33628 13748 33684
rect 12684 28700 12740 28756
rect 11564 28364 11620 28420
rect 10536 28250 10592 28252
rect 10536 28198 10538 28250
rect 10538 28198 10590 28250
rect 10590 28198 10592 28250
rect 10536 28196 10592 28198
rect 10640 28250 10696 28252
rect 10640 28198 10642 28250
rect 10642 28198 10694 28250
rect 10694 28198 10696 28250
rect 10640 28196 10696 28198
rect 10744 28250 10800 28252
rect 10744 28198 10746 28250
rect 10746 28198 10798 28250
rect 10798 28198 10800 28250
rect 10744 28196 10800 28198
rect 10108 27356 10164 27412
rect 10444 27298 10500 27300
rect 10444 27246 10446 27298
rect 10446 27246 10498 27298
rect 10498 27246 10500 27298
rect 10444 27244 10500 27246
rect 10220 26796 10276 26852
rect 9660 26236 9716 26292
rect 9772 25676 9828 25732
rect 10892 26796 10948 26852
rect 10536 26682 10592 26684
rect 10536 26630 10538 26682
rect 10538 26630 10590 26682
rect 10590 26630 10592 26682
rect 10536 26628 10592 26630
rect 10640 26682 10696 26684
rect 10640 26630 10642 26682
rect 10642 26630 10694 26682
rect 10694 26630 10696 26682
rect 10640 26628 10696 26630
rect 10744 26682 10800 26684
rect 10744 26630 10746 26682
rect 10746 26630 10798 26682
rect 10798 26630 10800 26682
rect 10744 26628 10800 26630
rect 10668 26290 10724 26292
rect 10668 26238 10670 26290
rect 10670 26238 10722 26290
rect 10722 26238 10724 26290
rect 10668 26236 10724 26238
rect 11676 27634 11732 27636
rect 11676 27582 11678 27634
rect 11678 27582 11730 27634
rect 11730 27582 11732 27634
rect 11676 27580 11732 27582
rect 12348 28476 12404 28532
rect 13132 28588 13188 28644
rect 11564 26178 11620 26180
rect 11564 26126 11566 26178
rect 11566 26126 11618 26178
rect 11618 26126 11620 26178
rect 11564 26124 11620 26126
rect 11564 25452 11620 25508
rect 11452 25282 11508 25284
rect 11452 25230 11454 25282
rect 11454 25230 11506 25282
rect 11506 25230 11508 25282
rect 11452 25228 11508 25230
rect 10536 25114 10592 25116
rect 10536 25062 10538 25114
rect 10538 25062 10590 25114
rect 10590 25062 10592 25114
rect 10536 25060 10592 25062
rect 10640 25114 10696 25116
rect 10640 25062 10642 25114
rect 10642 25062 10694 25114
rect 10694 25062 10696 25114
rect 10640 25060 10696 25062
rect 10744 25114 10800 25116
rect 10744 25062 10746 25114
rect 10746 25062 10798 25114
rect 10798 25062 10800 25114
rect 10744 25060 10800 25062
rect 10220 24834 10276 24836
rect 10220 24782 10222 24834
rect 10222 24782 10274 24834
rect 10274 24782 10276 24834
rect 10220 24780 10276 24782
rect 10108 23378 10164 23380
rect 10108 23326 10110 23378
rect 10110 23326 10162 23378
rect 10162 23326 10164 23378
rect 10108 23324 10164 23326
rect 10444 23938 10500 23940
rect 10444 23886 10446 23938
rect 10446 23886 10498 23938
rect 10498 23886 10500 23938
rect 10444 23884 10500 23886
rect 10536 23546 10592 23548
rect 10536 23494 10538 23546
rect 10538 23494 10590 23546
rect 10590 23494 10592 23546
rect 10536 23492 10592 23494
rect 10640 23546 10696 23548
rect 10640 23494 10642 23546
rect 10642 23494 10694 23546
rect 10694 23494 10696 23546
rect 10640 23492 10696 23494
rect 10744 23546 10800 23548
rect 10744 23494 10746 23546
rect 10746 23494 10798 23546
rect 10798 23494 10800 23546
rect 10744 23492 10800 23494
rect 9324 21084 9380 21140
rect 10332 22204 10388 22260
rect 11116 23324 11172 23380
rect 10536 21978 10592 21980
rect 10536 21926 10538 21978
rect 10538 21926 10590 21978
rect 10590 21926 10592 21978
rect 10536 21924 10592 21926
rect 10640 21978 10696 21980
rect 10640 21926 10642 21978
rect 10642 21926 10694 21978
rect 10694 21926 10696 21978
rect 10640 21924 10696 21926
rect 10744 21978 10800 21980
rect 10744 21926 10746 21978
rect 10746 21926 10798 21978
rect 10798 21926 10800 21978
rect 10744 21924 10800 21926
rect 11228 22146 11284 22148
rect 11228 22094 11230 22146
rect 11230 22094 11282 22146
rect 11282 22094 11284 22146
rect 11228 22092 11284 22094
rect 12460 25116 12516 25172
rect 11676 24668 11732 24724
rect 11788 23996 11844 24052
rect 12684 25452 12740 25508
rect 13692 29202 13748 29204
rect 13692 29150 13694 29202
rect 13694 29150 13746 29202
rect 13746 29150 13748 29202
rect 13692 29148 13748 29150
rect 13580 28642 13636 28644
rect 13580 28590 13582 28642
rect 13582 28590 13634 28642
rect 13634 28590 13636 28642
rect 13580 28588 13636 28590
rect 14140 33740 14196 33796
rect 14364 30156 14420 30212
rect 13916 28754 13972 28756
rect 13916 28702 13918 28754
rect 13918 28702 13970 28754
rect 13970 28702 13972 28754
rect 13916 28700 13972 28702
rect 13804 28588 13860 28644
rect 15198 35306 15254 35308
rect 15198 35254 15200 35306
rect 15200 35254 15252 35306
rect 15252 35254 15254 35306
rect 15198 35252 15254 35254
rect 15302 35306 15358 35308
rect 15302 35254 15304 35306
rect 15304 35254 15356 35306
rect 15356 35254 15358 35306
rect 15302 35252 15358 35254
rect 15406 35306 15462 35308
rect 15406 35254 15408 35306
rect 15408 35254 15460 35306
rect 15460 35254 15462 35306
rect 15406 35252 15462 35254
rect 15198 33738 15254 33740
rect 15198 33686 15200 33738
rect 15200 33686 15252 33738
rect 15252 33686 15254 33738
rect 15198 33684 15254 33686
rect 15302 33738 15358 33740
rect 15302 33686 15304 33738
rect 15304 33686 15356 33738
rect 15356 33686 15358 33738
rect 15302 33684 15358 33686
rect 15406 33738 15462 33740
rect 15406 33686 15408 33738
rect 15408 33686 15460 33738
rect 15460 33686 15462 33738
rect 15406 33684 15462 33686
rect 15198 32170 15254 32172
rect 15198 32118 15200 32170
rect 15200 32118 15252 32170
rect 15252 32118 15254 32170
rect 15198 32116 15254 32118
rect 15302 32170 15358 32172
rect 15302 32118 15304 32170
rect 15304 32118 15356 32170
rect 15356 32118 15358 32170
rect 15302 32116 15358 32118
rect 15406 32170 15462 32172
rect 15406 32118 15408 32170
rect 15408 32118 15460 32170
rect 15460 32118 15462 32170
rect 15406 32116 15462 32118
rect 15198 30602 15254 30604
rect 15198 30550 15200 30602
rect 15200 30550 15252 30602
rect 15252 30550 15254 30602
rect 15198 30548 15254 30550
rect 15302 30602 15358 30604
rect 15302 30550 15304 30602
rect 15304 30550 15356 30602
rect 15356 30550 15358 30602
rect 15302 30548 15358 30550
rect 15406 30602 15462 30604
rect 15406 30550 15408 30602
rect 15408 30550 15460 30602
rect 15460 30550 15462 30602
rect 15406 30548 15462 30550
rect 15596 30156 15652 30212
rect 14812 30044 14868 30100
rect 14252 28588 14308 28644
rect 13580 27634 13636 27636
rect 13580 27582 13582 27634
rect 13582 27582 13634 27634
rect 13634 27582 13636 27634
rect 13580 27580 13636 27582
rect 13580 27356 13636 27412
rect 12796 25394 12852 25396
rect 12796 25342 12798 25394
rect 12798 25342 12850 25394
rect 12850 25342 12852 25394
rect 12796 25340 12852 25342
rect 13020 25564 13076 25620
rect 13356 25340 13412 25396
rect 14140 26290 14196 26292
rect 14140 26238 14142 26290
rect 14142 26238 14194 26290
rect 14194 26238 14196 26290
rect 14140 26236 14196 26238
rect 13804 26178 13860 26180
rect 13804 26126 13806 26178
rect 13806 26126 13858 26178
rect 13858 26126 13860 26178
rect 13804 26124 13860 26126
rect 14028 25564 14084 25620
rect 14476 26514 14532 26516
rect 14476 26462 14478 26514
rect 14478 26462 14530 26514
rect 14530 26462 14532 26514
rect 14476 26460 14532 26462
rect 14476 25564 14532 25620
rect 14364 25228 14420 25284
rect 12572 24668 12628 24724
rect 12348 24050 12404 24052
rect 12348 23998 12350 24050
rect 12350 23998 12402 24050
rect 12402 23998 12404 24050
rect 12348 23996 12404 23998
rect 12572 23938 12628 23940
rect 12572 23886 12574 23938
rect 12574 23886 12626 23938
rect 12626 23886 12628 23938
rect 12572 23884 12628 23886
rect 12236 23266 12292 23268
rect 12236 23214 12238 23266
rect 12238 23214 12290 23266
rect 12290 23214 12292 23266
rect 12236 23212 12292 23214
rect 12124 22092 12180 22148
rect 11004 21698 11060 21700
rect 11004 21646 11006 21698
rect 11006 21646 11058 21698
rect 11058 21646 11060 21698
rect 11004 21644 11060 21646
rect 10332 21362 10388 21364
rect 10332 21310 10334 21362
rect 10334 21310 10386 21362
rect 10386 21310 10388 21362
rect 10332 21308 10388 21310
rect 10332 20914 10388 20916
rect 10332 20862 10334 20914
rect 10334 20862 10386 20914
rect 10386 20862 10388 20914
rect 10332 20860 10388 20862
rect 10536 20410 10592 20412
rect 10536 20358 10538 20410
rect 10538 20358 10590 20410
rect 10590 20358 10592 20410
rect 10536 20356 10592 20358
rect 10640 20410 10696 20412
rect 10640 20358 10642 20410
rect 10642 20358 10694 20410
rect 10694 20358 10696 20410
rect 10640 20356 10696 20358
rect 10744 20410 10800 20412
rect 10744 20358 10746 20410
rect 10746 20358 10798 20410
rect 10798 20358 10800 20410
rect 10744 20356 10800 20358
rect 2940 19740 2996 19796
rect 2492 19516 2548 19572
rect 5874 19626 5930 19628
rect 5874 19574 5876 19626
rect 5876 19574 5928 19626
rect 5928 19574 5930 19626
rect 5874 19572 5930 19574
rect 5978 19626 6034 19628
rect 5978 19574 5980 19626
rect 5980 19574 6032 19626
rect 6032 19574 6034 19626
rect 5978 19572 6034 19574
rect 6082 19626 6138 19628
rect 6082 19574 6084 19626
rect 6084 19574 6136 19626
rect 6136 19574 6138 19626
rect 6082 19572 6138 19574
rect 9660 19516 9716 19572
rect 10556 19292 10612 19348
rect 12348 22204 12404 22260
rect 12796 23938 12852 23940
rect 12796 23886 12798 23938
rect 12798 23886 12850 23938
rect 12850 23886 12852 23938
rect 12796 23884 12852 23886
rect 13804 24722 13860 24724
rect 13804 24670 13806 24722
rect 13806 24670 13858 24722
rect 13858 24670 13860 24722
rect 13804 24668 13860 24670
rect 14252 24722 14308 24724
rect 14252 24670 14254 24722
rect 14254 24670 14306 24722
rect 14306 24670 14308 24722
rect 14252 24668 14308 24670
rect 13244 23884 13300 23940
rect 13804 23884 13860 23940
rect 13692 23154 13748 23156
rect 13692 23102 13694 23154
rect 13694 23102 13746 23154
rect 13746 23102 13748 23154
rect 13692 23100 13748 23102
rect 14364 24556 14420 24612
rect 14028 24498 14084 24500
rect 14028 24446 14030 24498
rect 14030 24446 14082 24498
rect 14082 24446 14084 24498
rect 14028 24444 14084 24446
rect 12460 21980 12516 22036
rect 12572 22092 12628 22148
rect 12348 21868 12404 21924
rect 13468 22092 13524 22148
rect 13244 21810 13300 21812
rect 13244 21758 13246 21810
rect 13246 21758 13298 21810
rect 13298 21758 13300 21810
rect 13244 21756 13300 21758
rect 12572 21362 12628 21364
rect 12572 21310 12574 21362
rect 12574 21310 12626 21362
rect 12626 21310 12628 21362
rect 12572 21308 12628 21310
rect 12908 21586 12964 21588
rect 12908 21534 12910 21586
rect 12910 21534 12962 21586
rect 12962 21534 12964 21586
rect 12908 21532 12964 21534
rect 12572 20914 12628 20916
rect 12572 20862 12574 20914
rect 12574 20862 12626 20914
rect 12626 20862 12628 20914
rect 12572 20860 12628 20862
rect 13244 21308 13300 21364
rect 13468 21586 13524 21588
rect 13468 21534 13470 21586
rect 13470 21534 13522 21586
rect 13522 21534 13524 21586
rect 13468 21532 13524 21534
rect 2044 19010 2100 19012
rect 2044 18958 2046 19010
rect 2046 18958 2098 19010
rect 2098 18958 2100 19010
rect 2044 18956 2100 18958
rect 11228 19516 11284 19572
rect 12012 20018 12068 20020
rect 12012 19966 12014 20018
rect 12014 19966 12066 20018
rect 12066 19966 12068 20018
rect 12012 19964 12068 19966
rect 12572 19740 12628 19796
rect 12684 19964 12740 20020
rect 11452 19292 11508 19348
rect 1708 18844 1764 18900
rect 2492 18844 2548 18900
rect 2044 18450 2100 18452
rect 2044 18398 2046 18450
rect 2046 18398 2098 18450
rect 2098 18398 2100 18450
rect 2044 18396 2100 18398
rect 10536 18842 10592 18844
rect 10536 18790 10538 18842
rect 10538 18790 10590 18842
rect 10590 18790 10592 18842
rect 10536 18788 10592 18790
rect 10640 18842 10696 18844
rect 10640 18790 10642 18842
rect 10642 18790 10694 18842
rect 10694 18790 10696 18842
rect 10640 18788 10696 18790
rect 10744 18842 10800 18844
rect 10744 18790 10746 18842
rect 10746 18790 10798 18842
rect 10798 18790 10800 18842
rect 10744 18788 10800 18790
rect 1708 18172 1764 18228
rect 8764 18172 8820 18228
rect 5874 18058 5930 18060
rect 5874 18006 5876 18058
rect 5876 18006 5928 18058
rect 5928 18006 5930 18058
rect 5874 18004 5930 18006
rect 5978 18058 6034 18060
rect 5978 18006 5980 18058
rect 5980 18006 6032 18058
rect 6032 18006 6034 18058
rect 5978 18004 6034 18006
rect 6082 18058 6138 18060
rect 6082 18006 6084 18058
rect 6084 18006 6136 18058
rect 6136 18006 6138 18058
rect 6082 18004 6138 18006
rect 2716 17724 2772 17780
rect 10556 18226 10612 18228
rect 10556 18174 10558 18226
rect 10558 18174 10610 18226
rect 10610 18174 10612 18226
rect 10556 18172 10612 18174
rect 10108 18060 10164 18116
rect 10332 18060 10388 18116
rect 1708 17554 1764 17556
rect 1708 17502 1710 17554
rect 1710 17502 1762 17554
rect 1762 17502 1764 17554
rect 1708 17500 1764 17502
rect 2044 17554 2100 17556
rect 2044 17502 2046 17554
rect 2046 17502 2098 17554
rect 2098 17502 2100 17554
rect 2044 17500 2100 17502
rect 8428 17554 8484 17556
rect 8428 17502 8430 17554
rect 8430 17502 8482 17554
rect 8482 17502 8484 17554
rect 8428 17500 8484 17502
rect 2044 16994 2100 16996
rect 2044 16942 2046 16994
rect 2046 16942 2098 16994
rect 2098 16942 2100 16994
rect 2044 16940 2100 16942
rect 2380 16828 2436 16884
rect 2156 16716 2212 16772
rect 1708 16156 1764 16212
rect 2044 16604 2100 16660
rect 1708 15874 1764 15876
rect 1708 15822 1710 15874
rect 1710 15822 1762 15874
rect 1762 15822 1764 15874
rect 1708 15820 1764 15822
rect 10444 17890 10500 17892
rect 10444 17838 10446 17890
rect 10446 17838 10498 17890
rect 10498 17838 10500 17890
rect 10444 17836 10500 17838
rect 10892 18060 10948 18116
rect 10668 17500 10724 17556
rect 10536 17274 10592 17276
rect 10536 17222 10538 17274
rect 10538 17222 10590 17274
rect 10590 17222 10592 17274
rect 10536 17220 10592 17222
rect 10640 17274 10696 17276
rect 10640 17222 10642 17274
rect 10642 17222 10694 17274
rect 10694 17222 10696 17274
rect 10640 17220 10696 17222
rect 10744 17274 10800 17276
rect 10744 17222 10746 17274
rect 10746 17222 10798 17274
rect 10798 17222 10800 17274
rect 10744 17220 10800 17222
rect 10780 17052 10836 17108
rect 5874 16490 5930 16492
rect 5874 16438 5876 16490
rect 5876 16438 5928 16490
rect 5928 16438 5930 16490
rect 5874 16436 5930 16438
rect 5978 16490 6034 16492
rect 5978 16438 5980 16490
rect 5980 16438 6032 16490
rect 6032 16438 6034 16490
rect 5978 16436 6034 16438
rect 6082 16490 6138 16492
rect 6082 16438 6084 16490
rect 6084 16438 6136 16490
rect 6136 16438 6138 16490
rect 6082 16436 6138 16438
rect 8876 16268 8932 16324
rect 9772 16156 9828 16212
rect 2268 15820 2324 15876
rect 1708 14812 1764 14868
rect 1708 14306 1764 14308
rect 1708 14254 1710 14306
rect 1710 14254 1762 14306
rect 1762 14254 1764 14306
rect 1708 14252 1764 14254
rect 2044 14028 2100 14084
rect 2044 13858 2100 13860
rect 2044 13806 2046 13858
rect 2046 13806 2098 13858
rect 2098 13806 2100 13858
rect 2044 13804 2100 13806
rect 1708 13468 1764 13524
rect 2044 12962 2100 12964
rect 2044 12910 2046 12962
rect 2046 12910 2098 12962
rect 2098 12910 2100 12962
rect 2044 12908 2100 12910
rect 1708 12850 1764 12852
rect 1708 12798 1710 12850
rect 1710 12798 1762 12850
rect 1762 12798 1764 12850
rect 1708 12796 1764 12798
rect 8204 15484 8260 15540
rect 6300 15260 6356 15316
rect 5874 14922 5930 14924
rect 5874 14870 5876 14922
rect 5876 14870 5928 14922
rect 5928 14870 5930 14922
rect 5874 14868 5930 14870
rect 5978 14922 6034 14924
rect 5978 14870 5980 14922
rect 5980 14870 6032 14922
rect 6032 14870 6034 14922
rect 5978 14868 6034 14870
rect 6082 14922 6138 14924
rect 6082 14870 6084 14922
rect 6084 14870 6136 14922
rect 6136 14870 6138 14922
rect 6082 14868 6138 14870
rect 5874 13354 5930 13356
rect 5874 13302 5876 13354
rect 5876 13302 5928 13354
rect 5928 13302 5930 13354
rect 5874 13300 5930 13302
rect 5978 13354 6034 13356
rect 5978 13302 5980 13354
rect 5980 13302 6032 13354
rect 6032 13302 6034 13354
rect 5978 13300 6034 13302
rect 6082 13354 6138 13356
rect 6082 13302 6084 13354
rect 6084 13302 6136 13354
rect 6136 13302 6138 13354
rect 6082 13300 6138 13302
rect 2716 13132 2772 13188
rect 2380 12124 2436 12180
rect 5874 11786 5930 11788
rect 5874 11734 5876 11786
rect 5876 11734 5928 11786
rect 5928 11734 5930 11786
rect 5874 11732 5930 11734
rect 5978 11786 6034 11788
rect 5978 11734 5980 11786
rect 5980 11734 6032 11786
rect 6032 11734 6034 11786
rect 5978 11732 6034 11734
rect 6082 11786 6138 11788
rect 6082 11734 6084 11786
rect 6084 11734 6136 11786
rect 6136 11734 6138 11786
rect 6082 11732 6138 11734
rect 1708 11452 1764 11508
rect 2044 11452 2100 11508
rect 1708 11170 1764 11172
rect 1708 11118 1710 11170
rect 1710 11118 1762 11170
rect 1762 11118 1764 11170
rect 1708 11116 1764 11118
rect 2044 10722 2100 10724
rect 2044 10670 2046 10722
rect 2046 10670 2098 10722
rect 2098 10670 2100 10722
rect 2044 10668 2100 10670
rect 1708 10108 1764 10164
rect 5874 10218 5930 10220
rect 5874 10166 5876 10218
rect 5876 10166 5928 10218
rect 5928 10166 5930 10218
rect 5874 10164 5930 10166
rect 5978 10218 6034 10220
rect 5978 10166 5980 10218
rect 5980 10166 6032 10218
rect 6032 10166 6034 10218
rect 5978 10164 6034 10166
rect 6082 10218 6138 10220
rect 6082 10166 6084 10218
rect 6084 10166 6136 10218
rect 6136 10166 6138 10218
rect 6082 10164 6138 10166
rect 2044 9826 2100 9828
rect 2044 9774 2046 9826
rect 2046 9774 2098 9826
rect 2098 9774 2100 9826
rect 2044 9772 2100 9774
rect 1708 9602 1764 9604
rect 1708 9550 1710 9602
rect 1710 9550 1762 9602
rect 1762 9550 1764 9602
rect 1708 9548 1764 9550
rect 2044 9154 2100 9156
rect 2044 9102 2046 9154
rect 2046 9102 2098 9154
rect 2098 9102 2100 9154
rect 2044 9100 2100 9102
rect 1708 8764 1764 8820
rect 5874 8650 5930 8652
rect 5874 8598 5876 8650
rect 5876 8598 5928 8650
rect 5928 8598 5930 8650
rect 5874 8596 5930 8598
rect 5978 8650 6034 8652
rect 5978 8598 5980 8650
rect 5980 8598 6032 8650
rect 6032 8598 6034 8650
rect 5978 8596 6034 8598
rect 6082 8650 6138 8652
rect 6082 8598 6084 8650
rect 6084 8598 6136 8650
rect 6136 8598 6138 8650
rect 6082 8596 6138 8598
rect 2604 8316 2660 8372
rect 3164 8370 3220 8372
rect 3164 8318 3166 8370
rect 3166 8318 3218 8370
rect 3218 8318 3220 8370
rect 3164 8316 3220 8318
rect 1708 8146 1764 8148
rect 1708 8094 1710 8146
rect 1710 8094 1762 8146
rect 1762 8094 1764 8146
rect 1708 8092 1764 8094
rect 2380 7644 2436 7700
rect 2380 7362 2436 7364
rect 2380 7310 2382 7362
rect 2382 7310 2434 7362
rect 2434 7310 2436 7362
rect 2380 7308 2436 7310
rect 5874 7082 5930 7084
rect 5874 7030 5876 7082
rect 5876 7030 5928 7082
rect 5928 7030 5930 7082
rect 5874 7028 5930 7030
rect 5978 7082 6034 7084
rect 5978 7030 5980 7082
rect 5980 7030 6032 7082
rect 6032 7030 6034 7082
rect 5978 7028 6034 7030
rect 6082 7082 6138 7084
rect 6082 7030 6084 7082
rect 6084 7030 6136 7082
rect 6136 7030 6138 7082
rect 6082 7028 6138 7030
rect 5874 5514 5930 5516
rect 5874 5462 5876 5514
rect 5876 5462 5928 5514
rect 5928 5462 5930 5514
rect 5874 5460 5930 5462
rect 5978 5514 6034 5516
rect 5978 5462 5980 5514
rect 5980 5462 6032 5514
rect 6032 5462 6034 5514
rect 5978 5460 6034 5462
rect 6082 5514 6138 5516
rect 6082 5462 6084 5514
rect 6084 5462 6136 5514
rect 6136 5462 6138 5514
rect 6082 5460 6138 5462
rect 7644 14700 7700 14756
rect 6412 14588 6468 14644
rect 5874 3946 5930 3948
rect 5874 3894 5876 3946
rect 5876 3894 5928 3946
rect 5928 3894 5930 3946
rect 5874 3892 5930 3894
rect 5978 3946 6034 3948
rect 5978 3894 5980 3946
rect 5980 3894 6032 3946
rect 6032 3894 6034 3946
rect 5978 3892 6034 3894
rect 6082 3946 6138 3948
rect 6082 3894 6084 3946
rect 6084 3894 6136 3946
rect 6136 3894 6138 3946
rect 6082 3892 6138 3894
rect 6748 13692 6804 13748
rect 9100 15986 9156 15988
rect 9100 15934 9102 15986
rect 9102 15934 9154 15986
rect 9154 15934 9156 15986
rect 9100 15932 9156 15934
rect 10444 16770 10500 16772
rect 10444 16718 10446 16770
rect 10446 16718 10498 16770
rect 10498 16718 10500 16770
rect 10444 16716 10500 16718
rect 10332 16156 10388 16212
rect 10668 16380 10724 16436
rect 10108 15932 10164 15988
rect 11228 17052 11284 17108
rect 11116 16604 11172 16660
rect 10556 16210 10612 16212
rect 10556 16158 10558 16210
rect 10558 16158 10610 16210
rect 10610 16158 10612 16210
rect 10556 16156 10612 16158
rect 10444 15820 10500 15876
rect 10536 15706 10592 15708
rect 10536 15654 10538 15706
rect 10538 15654 10590 15706
rect 10590 15654 10592 15706
rect 10536 15652 10592 15654
rect 10640 15706 10696 15708
rect 10640 15654 10642 15706
rect 10642 15654 10694 15706
rect 10694 15654 10696 15706
rect 10640 15652 10696 15654
rect 10744 15706 10800 15708
rect 10744 15654 10746 15706
rect 10746 15654 10798 15706
rect 10798 15654 10800 15706
rect 10744 15652 10800 15654
rect 9548 15372 9604 15428
rect 9996 15426 10052 15428
rect 9996 15374 9998 15426
rect 9998 15374 10050 15426
rect 10050 15374 10052 15426
rect 9996 15372 10052 15374
rect 9212 14476 9268 14532
rect 9884 14418 9940 14420
rect 9884 14366 9886 14418
rect 9886 14366 9938 14418
rect 9938 14366 9940 14418
rect 9884 14364 9940 14366
rect 9548 12908 9604 12964
rect 9996 13580 10052 13636
rect 9884 12348 9940 12404
rect 8764 11116 8820 11172
rect 9548 3442 9604 3444
rect 9548 3390 9550 3442
rect 9550 3390 9602 3442
rect 9602 3390 9604 3442
rect 9548 3388 9604 3390
rect 10444 14812 10500 14868
rect 10220 14530 10276 14532
rect 10220 14478 10222 14530
rect 10222 14478 10274 14530
rect 10274 14478 10276 14530
rect 10220 14476 10276 14478
rect 10668 14530 10724 14532
rect 10668 14478 10670 14530
rect 10670 14478 10722 14530
rect 10722 14478 10724 14530
rect 10668 14476 10724 14478
rect 10332 14364 10388 14420
rect 10536 14138 10592 14140
rect 10536 14086 10538 14138
rect 10538 14086 10590 14138
rect 10590 14086 10592 14138
rect 10536 14084 10592 14086
rect 10640 14138 10696 14140
rect 10640 14086 10642 14138
rect 10642 14086 10694 14138
rect 10694 14086 10696 14138
rect 10640 14084 10696 14086
rect 10744 14138 10800 14140
rect 10744 14086 10746 14138
rect 10746 14086 10798 14138
rect 10798 14086 10800 14138
rect 10744 14084 10800 14086
rect 10556 13916 10612 13972
rect 10780 13356 10836 13412
rect 11452 15986 11508 15988
rect 11452 15934 11454 15986
rect 11454 15934 11506 15986
rect 11506 15934 11508 15986
rect 11452 15932 11508 15934
rect 11340 15708 11396 15764
rect 11340 15426 11396 15428
rect 11340 15374 11342 15426
rect 11342 15374 11394 15426
rect 11394 15374 11396 15426
rect 11340 15372 11396 15374
rect 11452 13858 11508 13860
rect 11452 13806 11454 13858
rect 11454 13806 11506 13858
rect 11506 13806 11508 13858
rect 11452 13804 11508 13806
rect 11116 13522 11172 13524
rect 11116 13470 11118 13522
rect 11118 13470 11170 13522
rect 11170 13470 11172 13522
rect 11116 13468 11172 13470
rect 10556 12962 10612 12964
rect 10556 12910 10558 12962
rect 10558 12910 10610 12962
rect 10610 12910 10612 12962
rect 10556 12908 10612 12910
rect 10536 12570 10592 12572
rect 10536 12518 10538 12570
rect 10538 12518 10590 12570
rect 10590 12518 10592 12570
rect 10536 12516 10592 12518
rect 10640 12570 10696 12572
rect 10640 12518 10642 12570
rect 10642 12518 10694 12570
rect 10694 12518 10696 12570
rect 10640 12516 10696 12518
rect 10744 12570 10800 12572
rect 10744 12518 10746 12570
rect 10746 12518 10798 12570
rect 10798 12518 10800 12570
rect 10744 12516 10800 12518
rect 10556 12236 10612 12292
rect 10556 12066 10612 12068
rect 10556 12014 10558 12066
rect 10558 12014 10610 12066
rect 10610 12014 10612 12066
rect 10556 12012 10612 12014
rect 10108 9772 10164 9828
rect 10332 11452 10388 11508
rect 12124 17948 12180 18004
rect 13244 20412 13300 20468
rect 13244 20018 13300 20020
rect 13244 19966 13246 20018
rect 13246 19966 13298 20018
rect 13298 19966 13300 20018
rect 13244 19964 13300 19966
rect 13692 21532 13748 21588
rect 13804 20690 13860 20692
rect 13804 20638 13806 20690
rect 13806 20638 13858 20690
rect 13858 20638 13860 20690
rect 13804 20636 13860 20638
rect 13692 20300 13748 20356
rect 14700 28364 14756 28420
rect 14812 28028 14868 28084
rect 15372 29314 15428 29316
rect 15372 29262 15374 29314
rect 15374 29262 15426 29314
rect 15426 29262 15428 29314
rect 15372 29260 15428 29262
rect 15036 29148 15092 29204
rect 15198 29034 15254 29036
rect 15198 28982 15200 29034
rect 15200 28982 15252 29034
rect 15252 28982 15254 29034
rect 15198 28980 15254 28982
rect 15302 29034 15358 29036
rect 15302 28982 15304 29034
rect 15304 28982 15356 29034
rect 15356 28982 15358 29034
rect 15302 28980 15358 28982
rect 15406 29034 15462 29036
rect 15406 28982 15408 29034
rect 15408 28982 15460 29034
rect 15460 28982 15462 29034
rect 15406 28980 15462 28982
rect 16044 36370 16100 36372
rect 16044 36318 16046 36370
rect 16046 36318 16098 36370
rect 16098 36318 16100 36370
rect 16044 36316 16100 36318
rect 15820 29426 15876 29428
rect 15820 29374 15822 29426
rect 15822 29374 15874 29426
rect 15874 29374 15876 29426
rect 15820 29372 15876 29374
rect 16268 29314 16324 29316
rect 16268 29262 16270 29314
rect 16270 29262 16322 29314
rect 16322 29262 16324 29314
rect 16268 29260 16324 29262
rect 16156 29202 16212 29204
rect 16156 29150 16158 29202
rect 16158 29150 16210 29202
rect 16210 29150 16212 29202
rect 16156 29148 16212 29150
rect 15820 28866 15876 28868
rect 15820 28814 15822 28866
rect 15822 28814 15874 28866
rect 15874 28814 15876 28866
rect 15820 28812 15876 28814
rect 15708 28028 15764 28084
rect 15596 27970 15652 27972
rect 15596 27918 15598 27970
rect 15598 27918 15650 27970
rect 15650 27918 15652 27970
rect 15596 27916 15652 27918
rect 14700 26290 14756 26292
rect 14700 26238 14702 26290
rect 14702 26238 14754 26290
rect 14754 26238 14756 26290
rect 14700 26236 14756 26238
rect 14700 25788 14756 25844
rect 15198 27466 15254 27468
rect 15198 27414 15200 27466
rect 15200 27414 15252 27466
rect 15252 27414 15254 27466
rect 15198 27412 15254 27414
rect 15302 27466 15358 27468
rect 15302 27414 15304 27466
rect 15304 27414 15356 27466
rect 15356 27414 15358 27466
rect 15302 27412 15358 27414
rect 15406 27466 15462 27468
rect 15406 27414 15408 27466
rect 15408 27414 15460 27466
rect 15460 27414 15462 27466
rect 15406 27412 15462 27414
rect 15932 27634 15988 27636
rect 15932 27582 15934 27634
rect 15934 27582 15986 27634
rect 15986 27582 15988 27634
rect 15932 27580 15988 27582
rect 16156 28028 16212 28084
rect 15036 27244 15092 27300
rect 15372 27074 15428 27076
rect 15372 27022 15374 27074
rect 15374 27022 15426 27074
rect 15426 27022 15428 27074
rect 15372 27020 15428 27022
rect 15708 26460 15764 26516
rect 15596 26402 15652 26404
rect 15596 26350 15598 26402
rect 15598 26350 15650 26402
rect 15650 26350 15652 26402
rect 15596 26348 15652 26350
rect 16156 26796 16212 26852
rect 15708 26124 15764 26180
rect 15820 26012 15876 26068
rect 15036 25788 15092 25844
rect 15198 25898 15254 25900
rect 15198 25846 15200 25898
rect 15200 25846 15252 25898
rect 15252 25846 15254 25898
rect 15198 25844 15254 25846
rect 15302 25898 15358 25900
rect 15302 25846 15304 25898
rect 15304 25846 15356 25898
rect 15356 25846 15358 25898
rect 15302 25844 15358 25846
rect 15406 25898 15462 25900
rect 15406 25846 15408 25898
rect 15408 25846 15460 25898
rect 15460 25846 15462 25898
rect 15406 25844 15462 25846
rect 14924 25618 14980 25620
rect 14924 25566 14926 25618
rect 14926 25566 14978 25618
rect 14978 25566 14980 25618
rect 14924 25564 14980 25566
rect 14700 24444 14756 24500
rect 14588 23884 14644 23940
rect 14364 23826 14420 23828
rect 14364 23774 14366 23826
rect 14366 23774 14418 23826
rect 14418 23774 14420 23826
rect 14364 23772 14420 23774
rect 14812 23154 14868 23156
rect 14812 23102 14814 23154
rect 14814 23102 14866 23154
rect 14866 23102 14868 23154
rect 14812 23100 14868 23102
rect 15148 25506 15204 25508
rect 15148 25454 15150 25506
rect 15150 25454 15202 25506
rect 15202 25454 15204 25506
rect 15148 25452 15204 25454
rect 15148 25228 15204 25284
rect 16268 26572 16324 26628
rect 16268 26012 16324 26068
rect 16940 29484 16996 29540
rect 16716 29426 16772 29428
rect 16716 29374 16718 29426
rect 16718 29374 16770 29426
rect 16770 29374 16772 29426
rect 16716 29372 16772 29374
rect 16492 29148 16548 29204
rect 16604 28812 16660 28868
rect 17388 35756 17444 35812
rect 17388 29372 17444 29428
rect 17276 28588 17332 28644
rect 17500 27916 17556 27972
rect 17724 35532 17780 35588
rect 16828 27692 16884 27748
rect 17500 27746 17556 27748
rect 17500 27694 17502 27746
rect 17502 27694 17554 27746
rect 17554 27694 17556 27746
rect 17500 27692 17556 27694
rect 17388 27634 17444 27636
rect 17388 27582 17390 27634
rect 17390 27582 17442 27634
rect 17442 27582 17444 27634
rect 17388 27580 17444 27582
rect 17948 31836 18004 31892
rect 18396 29986 18452 29988
rect 18396 29934 18398 29986
rect 18398 29934 18450 29986
rect 18450 29934 18452 29986
rect 18396 29932 18452 29934
rect 17948 29426 18004 29428
rect 17948 29374 17950 29426
rect 17950 29374 18002 29426
rect 18002 29374 18004 29426
rect 17948 29372 18004 29374
rect 17948 29148 18004 29204
rect 18508 29372 18564 29428
rect 18620 36316 18676 36372
rect 18732 31836 18788 31892
rect 19292 29932 19348 29988
rect 19628 29650 19684 29652
rect 19628 29598 19630 29650
rect 19630 29598 19682 29650
rect 19682 29598 19684 29650
rect 19628 29596 19684 29598
rect 19516 29484 19572 29540
rect 18396 29148 18452 29204
rect 18956 28418 19012 28420
rect 18956 28366 18958 28418
rect 18958 28366 19010 28418
rect 19010 28366 19012 28418
rect 18956 28364 19012 28366
rect 17948 27916 18004 27972
rect 18060 27468 18116 27524
rect 18172 27692 18228 27748
rect 17836 27020 17892 27076
rect 17388 26908 17444 26964
rect 17612 26962 17668 26964
rect 17612 26910 17614 26962
rect 17614 26910 17666 26962
rect 17666 26910 17668 26962
rect 17612 26908 17668 26910
rect 16604 26514 16660 26516
rect 16604 26462 16606 26514
rect 16606 26462 16658 26514
rect 16658 26462 16660 26514
rect 16604 26460 16660 26462
rect 17948 26796 18004 26852
rect 17948 26572 18004 26628
rect 17164 26348 17220 26404
rect 16604 25676 16660 25732
rect 15820 25282 15876 25284
rect 15820 25230 15822 25282
rect 15822 25230 15874 25282
rect 15874 25230 15876 25282
rect 15820 25228 15876 25230
rect 15932 25004 15988 25060
rect 15198 24330 15254 24332
rect 15198 24278 15200 24330
rect 15200 24278 15252 24330
rect 15252 24278 15254 24330
rect 15198 24276 15254 24278
rect 15302 24330 15358 24332
rect 15302 24278 15304 24330
rect 15304 24278 15356 24330
rect 15356 24278 15358 24330
rect 15302 24276 15358 24278
rect 15406 24330 15462 24332
rect 15406 24278 15408 24330
rect 15408 24278 15460 24330
rect 15460 24278 15462 24330
rect 15406 24276 15462 24278
rect 16604 25452 16660 25508
rect 16380 25228 16436 25284
rect 16492 25004 16548 25060
rect 16268 24892 16324 24948
rect 15596 23212 15652 23268
rect 14140 22316 14196 22372
rect 14588 22540 14644 22596
rect 14476 22428 14532 22484
rect 14700 22204 14756 22260
rect 15198 22762 15254 22764
rect 15198 22710 15200 22762
rect 15200 22710 15252 22762
rect 15252 22710 15254 22762
rect 15198 22708 15254 22710
rect 15302 22762 15358 22764
rect 15302 22710 15304 22762
rect 15304 22710 15356 22762
rect 15356 22710 15358 22762
rect 15302 22708 15358 22710
rect 15406 22762 15462 22764
rect 15406 22710 15408 22762
rect 15408 22710 15460 22762
rect 15460 22710 15462 22762
rect 15406 22708 15462 22710
rect 15484 22258 15540 22260
rect 15484 22206 15486 22258
rect 15486 22206 15538 22258
rect 15538 22206 15540 22258
rect 15484 22204 15540 22206
rect 16044 24780 16100 24836
rect 16940 26012 16996 26068
rect 16716 25228 16772 25284
rect 16828 24780 16884 24836
rect 16940 25452 16996 25508
rect 16492 23772 16548 23828
rect 16380 23100 16436 23156
rect 15820 22146 15876 22148
rect 15820 22094 15822 22146
rect 15822 22094 15874 22146
rect 15874 22094 15876 22146
rect 15820 22092 15876 22094
rect 14476 21308 14532 21364
rect 15036 21532 15092 21588
rect 14364 20914 14420 20916
rect 14364 20862 14366 20914
rect 14366 20862 14418 20914
rect 14418 20862 14420 20914
rect 14364 20860 14420 20862
rect 14140 20636 14196 20692
rect 14588 20636 14644 20692
rect 14252 20578 14308 20580
rect 14252 20526 14254 20578
rect 14254 20526 14306 20578
rect 14306 20526 14308 20578
rect 14252 20524 14308 20526
rect 15260 21980 15316 22036
rect 15708 21868 15764 21924
rect 14924 21362 14980 21364
rect 14924 21310 14926 21362
rect 14926 21310 14978 21362
rect 14978 21310 14980 21362
rect 14924 21308 14980 21310
rect 14924 21084 14980 21140
rect 15198 21194 15254 21196
rect 15198 21142 15200 21194
rect 15200 21142 15252 21194
rect 15252 21142 15254 21194
rect 15198 21140 15254 21142
rect 15302 21194 15358 21196
rect 15302 21142 15304 21194
rect 15304 21142 15356 21194
rect 15356 21142 15358 21194
rect 15302 21140 15358 21142
rect 15406 21194 15462 21196
rect 15406 21142 15408 21194
rect 15408 21142 15460 21194
rect 15460 21142 15462 21194
rect 15406 21140 15462 21142
rect 15596 20748 15652 20804
rect 15148 20636 15204 20692
rect 14924 20300 14980 20356
rect 13468 18732 13524 18788
rect 13020 18450 13076 18452
rect 13020 18398 13022 18450
rect 13022 18398 13074 18450
rect 13074 18398 13076 18450
rect 13020 18396 13076 18398
rect 11676 17500 11732 17556
rect 11676 16716 11732 16772
rect 12684 17836 12740 17892
rect 12908 17948 12964 18004
rect 12572 17500 12628 17556
rect 13692 18450 13748 18452
rect 13692 18398 13694 18450
rect 13694 18398 13746 18450
rect 13746 18398 13748 18450
rect 13692 18396 13748 18398
rect 13356 18284 13412 18340
rect 12684 16492 12740 16548
rect 13020 16882 13076 16884
rect 13020 16830 13022 16882
rect 13022 16830 13074 16882
rect 13074 16830 13076 16882
rect 13020 16828 13076 16830
rect 12572 16210 12628 16212
rect 12572 16158 12574 16210
rect 12574 16158 12626 16210
rect 12626 16158 12628 16210
rect 12572 16156 12628 16158
rect 12012 15932 12068 15988
rect 11676 15708 11732 15764
rect 12796 16098 12852 16100
rect 12796 16046 12798 16098
rect 12798 16046 12850 16098
rect 12850 16046 12852 16098
rect 12796 16044 12852 16046
rect 12348 15932 12404 15988
rect 12460 15820 12516 15876
rect 11900 14418 11956 14420
rect 11900 14366 11902 14418
rect 11902 14366 11954 14418
rect 11954 14366 11956 14418
rect 11900 14364 11956 14366
rect 11676 13468 11732 13524
rect 11004 11676 11060 11732
rect 10536 11002 10592 11004
rect 10536 10950 10538 11002
rect 10538 10950 10590 11002
rect 10590 10950 10592 11002
rect 10536 10948 10592 10950
rect 10640 11002 10696 11004
rect 10640 10950 10642 11002
rect 10642 10950 10694 11002
rect 10694 10950 10696 11002
rect 10640 10948 10696 10950
rect 10744 11002 10800 11004
rect 10744 10950 10746 11002
rect 10746 10950 10798 11002
rect 10798 10950 10800 11002
rect 10744 10948 10800 10950
rect 10536 9434 10592 9436
rect 10536 9382 10538 9434
rect 10538 9382 10590 9434
rect 10590 9382 10592 9434
rect 10536 9380 10592 9382
rect 10640 9434 10696 9436
rect 10640 9382 10642 9434
rect 10642 9382 10694 9434
rect 10694 9382 10696 9434
rect 10640 9380 10696 9382
rect 10744 9434 10800 9436
rect 10744 9382 10746 9434
rect 10746 9382 10798 9434
rect 10798 9382 10800 9434
rect 10744 9380 10800 9382
rect 10332 9100 10388 9156
rect 10536 7866 10592 7868
rect 10536 7814 10538 7866
rect 10538 7814 10590 7866
rect 10590 7814 10592 7866
rect 10536 7812 10592 7814
rect 10640 7866 10696 7868
rect 10640 7814 10642 7866
rect 10642 7814 10694 7866
rect 10694 7814 10696 7866
rect 10640 7812 10696 7814
rect 10744 7866 10800 7868
rect 10744 7814 10746 7866
rect 10746 7814 10798 7866
rect 10798 7814 10800 7866
rect 10744 7812 10800 7814
rect 10536 6298 10592 6300
rect 10536 6246 10538 6298
rect 10538 6246 10590 6298
rect 10590 6246 10592 6298
rect 10536 6244 10592 6246
rect 10640 6298 10696 6300
rect 10640 6246 10642 6298
rect 10642 6246 10694 6298
rect 10694 6246 10696 6298
rect 10640 6244 10696 6246
rect 10744 6298 10800 6300
rect 10744 6246 10746 6298
rect 10746 6246 10798 6298
rect 10798 6246 10800 6298
rect 10744 6244 10800 6246
rect 10536 4730 10592 4732
rect 10536 4678 10538 4730
rect 10538 4678 10590 4730
rect 10590 4678 10592 4730
rect 10536 4676 10592 4678
rect 10640 4730 10696 4732
rect 10640 4678 10642 4730
rect 10642 4678 10694 4730
rect 10694 4678 10696 4730
rect 10640 4676 10696 4678
rect 10744 4730 10800 4732
rect 10744 4678 10746 4730
rect 10746 4678 10798 4730
rect 10798 4678 10800 4730
rect 10744 4676 10800 4678
rect 10108 3388 10164 3444
rect 11004 10668 11060 10724
rect 11340 12236 11396 12292
rect 11676 12236 11732 12292
rect 11228 8316 11284 8372
rect 12572 14306 12628 14308
rect 12572 14254 12574 14306
rect 12574 14254 12626 14306
rect 12626 14254 12628 14306
rect 12572 14252 12628 14254
rect 12460 14140 12516 14196
rect 12796 14252 12852 14308
rect 12908 14364 12964 14420
rect 12796 13916 12852 13972
rect 12236 12348 12292 12404
rect 12012 12066 12068 12068
rect 12012 12014 12014 12066
rect 12014 12014 12066 12066
rect 12066 12014 12068 12066
rect 12012 12012 12068 12014
rect 11676 11954 11732 11956
rect 11676 11902 11678 11954
rect 11678 11902 11730 11954
rect 11730 11902 11732 11954
rect 11676 11900 11732 11902
rect 12796 12684 12852 12740
rect 13244 14140 13300 14196
rect 13580 16882 13636 16884
rect 13580 16830 13582 16882
rect 13582 16830 13634 16882
rect 13634 16830 13636 16882
rect 13580 16828 13636 16830
rect 14476 19404 14532 19460
rect 14700 19516 14756 19572
rect 14364 19010 14420 19012
rect 14364 18958 14366 19010
rect 14366 18958 14418 19010
rect 14418 18958 14420 19010
rect 14364 18956 14420 18958
rect 14252 18732 14308 18788
rect 14252 18338 14308 18340
rect 14252 18286 14254 18338
rect 14254 18286 14306 18338
rect 14306 18286 14308 18338
rect 14252 18284 14308 18286
rect 13468 15986 13524 15988
rect 13468 15934 13470 15986
rect 13470 15934 13522 15986
rect 13522 15934 13524 15986
rect 13468 15932 13524 15934
rect 13804 15986 13860 15988
rect 13804 15934 13806 15986
rect 13806 15934 13858 15986
rect 13858 15934 13860 15986
rect 13804 15932 13860 15934
rect 14140 16044 14196 16100
rect 14028 15932 14084 15988
rect 13132 13356 13188 13412
rect 13132 12796 13188 12852
rect 13916 14530 13972 14532
rect 13916 14478 13918 14530
rect 13918 14478 13970 14530
rect 13970 14478 13972 14530
rect 13916 14476 13972 14478
rect 13692 14364 13748 14420
rect 13580 14306 13636 14308
rect 13580 14254 13582 14306
rect 13582 14254 13634 14306
rect 13634 14254 13636 14306
rect 13580 14252 13636 14254
rect 13468 13916 13524 13972
rect 12684 11900 12740 11956
rect 12572 11788 12628 11844
rect 12460 11676 12516 11732
rect 12348 11340 12404 11396
rect 12348 8428 12404 8484
rect 13356 13132 13412 13188
rect 15372 20524 15428 20580
rect 16380 21308 16436 21364
rect 15708 20636 15764 20692
rect 16268 20412 16324 20468
rect 15198 19626 15254 19628
rect 15198 19574 15200 19626
rect 15200 19574 15252 19626
rect 15252 19574 15254 19626
rect 15198 19572 15254 19574
rect 15302 19626 15358 19628
rect 15302 19574 15304 19626
rect 15304 19574 15356 19626
rect 15356 19574 15358 19626
rect 15302 19572 15358 19574
rect 15406 19626 15462 19628
rect 15406 19574 15408 19626
rect 15408 19574 15460 19626
rect 15460 19574 15462 19626
rect 15406 19572 15462 19574
rect 15596 19404 15652 19460
rect 14700 18620 14756 18676
rect 14812 17836 14868 17892
rect 14588 17052 14644 17108
rect 14476 15484 14532 15540
rect 14812 17666 14868 17668
rect 14812 17614 14814 17666
rect 14814 17614 14866 17666
rect 14866 17614 14868 17666
rect 14812 17612 14868 17614
rect 14812 16492 14868 16548
rect 15932 19122 15988 19124
rect 15932 19070 15934 19122
rect 15934 19070 15986 19122
rect 15986 19070 15988 19122
rect 15932 19068 15988 19070
rect 16380 20018 16436 20020
rect 16380 19966 16382 20018
rect 16382 19966 16434 20018
rect 16434 19966 16436 20018
rect 16380 19964 16436 19966
rect 15372 18956 15428 19012
rect 15372 18284 15428 18340
rect 15198 18058 15254 18060
rect 15198 18006 15200 18058
rect 15200 18006 15252 18058
rect 15252 18006 15254 18058
rect 15198 18004 15254 18006
rect 15302 18058 15358 18060
rect 15302 18006 15304 18058
rect 15304 18006 15356 18058
rect 15356 18006 15358 18058
rect 15302 18004 15358 18006
rect 15406 18058 15462 18060
rect 15406 18006 15408 18058
rect 15408 18006 15460 18058
rect 15460 18006 15462 18058
rect 15406 18004 15462 18006
rect 15148 17724 15204 17780
rect 15484 17836 15540 17892
rect 14588 14364 14644 14420
rect 14252 14252 14308 14308
rect 14028 13132 14084 13188
rect 13916 12962 13972 12964
rect 13916 12910 13918 12962
rect 13918 12910 13970 12962
rect 13970 12910 13972 12962
rect 13916 12908 13972 12910
rect 13580 12738 13636 12740
rect 13580 12686 13582 12738
rect 13582 12686 13634 12738
rect 13634 12686 13636 12738
rect 13580 12684 13636 12686
rect 14364 13634 14420 13636
rect 14364 13582 14366 13634
rect 14366 13582 14418 13634
rect 14418 13582 14420 13634
rect 14364 13580 14420 13582
rect 15148 16940 15204 16996
rect 15036 16882 15092 16884
rect 15036 16830 15038 16882
rect 15038 16830 15090 16882
rect 15090 16830 15092 16882
rect 15036 16828 15092 16830
rect 16156 18172 16212 18228
rect 16156 17724 16212 17780
rect 15708 17500 15764 17556
rect 15596 17442 15652 17444
rect 15596 17390 15598 17442
rect 15598 17390 15650 17442
rect 15650 17390 15652 17442
rect 15596 17388 15652 17390
rect 16716 21868 16772 21924
rect 16828 21308 16884 21364
rect 16604 20690 16660 20692
rect 16604 20638 16606 20690
rect 16606 20638 16658 20690
rect 16658 20638 16660 20690
rect 16604 20636 16660 20638
rect 16604 19122 16660 19124
rect 16604 19070 16606 19122
rect 16606 19070 16658 19122
rect 16658 19070 16660 19122
rect 16604 19068 16660 19070
rect 16604 18508 16660 18564
rect 15932 16882 15988 16884
rect 15932 16830 15934 16882
rect 15934 16830 15986 16882
rect 15986 16830 15988 16882
rect 15932 16828 15988 16830
rect 16492 16994 16548 16996
rect 16492 16942 16494 16994
rect 16494 16942 16546 16994
rect 16546 16942 16548 16994
rect 16492 16940 16548 16942
rect 15148 16770 15204 16772
rect 15148 16718 15150 16770
rect 15150 16718 15202 16770
rect 15202 16718 15204 16770
rect 15148 16716 15204 16718
rect 15198 16490 15254 16492
rect 15198 16438 15200 16490
rect 15200 16438 15252 16490
rect 15252 16438 15254 16490
rect 15198 16436 15254 16438
rect 15302 16490 15358 16492
rect 15302 16438 15304 16490
rect 15304 16438 15356 16490
rect 15356 16438 15358 16490
rect 15302 16436 15358 16438
rect 15406 16490 15462 16492
rect 15406 16438 15408 16490
rect 15408 16438 15460 16490
rect 15460 16438 15462 16490
rect 15406 16436 15462 16438
rect 15484 16156 15540 16212
rect 15820 15708 15876 15764
rect 15596 15484 15652 15540
rect 15198 14922 15254 14924
rect 15198 14870 15200 14922
rect 15200 14870 15252 14922
rect 15252 14870 15254 14922
rect 15198 14868 15254 14870
rect 15302 14922 15358 14924
rect 15302 14870 15304 14922
rect 15304 14870 15356 14922
rect 15356 14870 15358 14922
rect 15302 14868 15358 14870
rect 15406 14922 15462 14924
rect 15406 14870 15408 14922
rect 15408 14870 15460 14922
rect 15460 14870 15462 14922
rect 15406 14868 15462 14870
rect 14924 14530 14980 14532
rect 14924 14478 14926 14530
rect 14926 14478 14978 14530
rect 14978 14478 14980 14530
rect 14924 14476 14980 14478
rect 15596 14530 15652 14532
rect 15596 14478 15598 14530
rect 15598 14478 15650 14530
rect 15650 14478 15652 14530
rect 15596 14476 15652 14478
rect 14812 13132 14868 13188
rect 15708 14252 15764 14308
rect 15708 13634 15764 13636
rect 15708 13582 15710 13634
rect 15710 13582 15762 13634
rect 15762 13582 15764 13634
rect 15708 13580 15764 13582
rect 14924 12962 14980 12964
rect 14924 12910 14926 12962
rect 14926 12910 14978 12962
rect 14978 12910 14980 12962
rect 14924 12908 14980 12910
rect 14252 12460 14308 12516
rect 13356 12348 13412 12404
rect 13804 12290 13860 12292
rect 13804 12238 13806 12290
rect 13806 12238 13858 12290
rect 13858 12238 13860 12290
rect 13804 12236 13860 12238
rect 13468 12178 13524 12180
rect 13468 12126 13470 12178
rect 13470 12126 13522 12178
rect 13522 12126 13524 12178
rect 13468 12124 13524 12126
rect 14028 12178 14084 12180
rect 14028 12126 14030 12178
rect 14030 12126 14082 12178
rect 14082 12126 14084 12178
rect 14028 12124 14084 12126
rect 13804 11900 13860 11956
rect 13692 11394 13748 11396
rect 13692 11342 13694 11394
rect 13694 11342 13746 11394
rect 13746 11342 13748 11394
rect 13692 11340 13748 11342
rect 13468 8428 13524 8484
rect 13244 7308 13300 7364
rect 14476 3500 14532 3556
rect 10536 3162 10592 3164
rect 10536 3110 10538 3162
rect 10538 3110 10590 3162
rect 10590 3110 10592 3162
rect 10536 3108 10592 3110
rect 10640 3162 10696 3164
rect 10640 3110 10642 3162
rect 10642 3110 10694 3162
rect 10694 3110 10696 3162
rect 10640 3108 10696 3110
rect 10744 3162 10800 3164
rect 10744 3110 10746 3162
rect 10746 3110 10798 3162
rect 10798 3110 10800 3162
rect 10744 3108 10800 3110
rect 15198 13354 15254 13356
rect 15198 13302 15200 13354
rect 15200 13302 15252 13354
rect 15252 13302 15254 13354
rect 15198 13300 15254 13302
rect 15302 13354 15358 13356
rect 15302 13302 15304 13354
rect 15304 13302 15356 13354
rect 15356 13302 15358 13354
rect 15302 13300 15358 13302
rect 15406 13354 15462 13356
rect 15406 13302 15408 13354
rect 15408 13302 15460 13354
rect 15460 13302 15462 13354
rect 15406 13300 15462 13302
rect 15260 13186 15316 13188
rect 15260 13134 15262 13186
rect 15262 13134 15314 13186
rect 15314 13134 15316 13186
rect 15260 13132 15316 13134
rect 15148 12796 15204 12852
rect 15372 12908 15428 12964
rect 16380 16658 16436 16660
rect 16380 16606 16382 16658
rect 16382 16606 16434 16658
rect 16434 16606 16436 16658
rect 16380 16604 16436 16606
rect 16268 15874 16324 15876
rect 16268 15822 16270 15874
rect 16270 15822 16322 15874
rect 16322 15822 16324 15874
rect 16268 15820 16324 15822
rect 17500 26402 17556 26404
rect 17500 26350 17502 26402
rect 17502 26350 17554 26402
rect 17554 26350 17556 26402
rect 17500 26348 17556 26350
rect 17948 25564 18004 25620
rect 17388 25506 17444 25508
rect 17388 25454 17390 25506
rect 17390 25454 17442 25506
rect 17442 25454 17444 25506
rect 17388 25452 17444 25454
rect 17612 25394 17668 25396
rect 17612 25342 17614 25394
rect 17614 25342 17666 25394
rect 17666 25342 17668 25394
rect 17612 25340 17668 25342
rect 17388 24946 17444 24948
rect 17388 24894 17390 24946
rect 17390 24894 17442 24946
rect 17442 24894 17444 24946
rect 17388 24892 17444 24894
rect 17724 25116 17780 25172
rect 17948 25116 18004 25172
rect 17164 24668 17220 24724
rect 17612 24722 17668 24724
rect 17612 24670 17614 24722
rect 17614 24670 17666 24722
rect 17666 24670 17668 24722
rect 17612 24668 17668 24670
rect 17612 24332 17668 24388
rect 16828 20412 16884 20468
rect 17388 23884 17444 23940
rect 17388 23154 17444 23156
rect 17388 23102 17390 23154
rect 17390 23102 17442 23154
rect 17442 23102 17444 23154
rect 17388 23100 17444 23102
rect 17276 22146 17332 22148
rect 17276 22094 17278 22146
rect 17278 22094 17330 22146
rect 17330 22094 17332 22146
rect 17276 22092 17332 22094
rect 17388 21586 17444 21588
rect 17388 21534 17390 21586
rect 17390 21534 17442 21586
rect 17442 21534 17444 21586
rect 17388 21532 17444 21534
rect 17388 20972 17444 21028
rect 17388 20636 17444 20692
rect 17276 20578 17332 20580
rect 17276 20526 17278 20578
rect 17278 20526 17330 20578
rect 17330 20526 17332 20578
rect 17276 20524 17332 20526
rect 16940 20076 16996 20132
rect 16828 20018 16884 20020
rect 16828 19966 16830 20018
rect 16830 19966 16882 20018
rect 16882 19966 16884 20018
rect 16828 19964 16884 19966
rect 17724 23826 17780 23828
rect 17724 23774 17726 23826
rect 17726 23774 17778 23826
rect 17778 23774 17780 23826
rect 17724 23772 17780 23774
rect 18508 27074 18564 27076
rect 18508 27022 18510 27074
rect 18510 27022 18562 27074
rect 18562 27022 18564 27074
rect 18508 27020 18564 27022
rect 18396 26962 18452 26964
rect 18396 26910 18398 26962
rect 18398 26910 18450 26962
rect 18450 26910 18452 26962
rect 18396 26908 18452 26910
rect 17948 23436 18004 23492
rect 17724 21810 17780 21812
rect 17724 21758 17726 21810
rect 17726 21758 17778 21810
rect 17778 21758 17780 21810
rect 17724 21756 17780 21758
rect 18396 24610 18452 24612
rect 18396 24558 18398 24610
rect 18398 24558 18450 24610
rect 18450 24558 18452 24610
rect 18396 24556 18452 24558
rect 18284 24498 18340 24500
rect 18284 24446 18286 24498
rect 18286 24446 18338 24498
rect 18338 24446 18340 24498
rect 18284 24444 18340 24446
rect 19180 26402 19236 26404
rect 19180 26350 19182 26402
rect 19182 26350 19234 26402
rect 19234 26350 19236 26402
rect 19180 26348 19236 26350
rect 19516 26012 19572 26068
rect 18956 25730 19012 25732
rect 18956 25678 18958 25730
rect 18958 25678 19010 25730
rect 19010 25678 19012 25730
rect 18956 25676 19012 25678
rect 18844 25618 18900 25620
rect 18844 25566 18846 25618
rect 18846 25566 18898 25618
rect 18898 25566 18900 25618
rect 18844 25564 18900 25566
rect 20748 36316 20804 36372
rect 19860 36090 19916 36092
rect 19860 36038 19862 36090
rect 19862 36038 19914 36090
rect 19914 36038 19916 36090
rect 19860 36036 19916 36038
rect 19964 36090 20020 36092
rect 19964 36038 19966 36090
rect 19966 36038 20018 36090
rect 20018 36038 20020 36090
rect 19964 36036 20020 36038
rect 20068 36090 20124 36092
rect 20068 36038 20070 36090
rect 20070 36038 20122 36090
rect 20122 36038 20124 36090
rect 20068 36036 20124 36038
rect 19860 34522 19916 34524
rect 19860 34470 19862 34522
rect 19862 34470 19914 34522
rect 19914 34470 19916 34522
rect 19860 34468 19916 34470
rect 19964 34522 20020 34524
rect 19964 34470 19966 34522
rect 19966 34470 20018 34522
rect 20018 34470 20020 34522
rect 19964 34468 20020 34470
rect 20068 34522 20124 34524
rect 20068 34470 20070 34522
rect 20070 34470 20122 34522
rect 20122 34470 20124 34522
rect 20068 34468 20124 34470
rect 19860 32954 19916 32956
rect 19860 32902 19862 32954
rect 19862 32902 19914 32954
rect 19914 32902 19916 32954
rect 19860 32900 19916 32902
rect 19964 32954 20020 32956
rect 19964 32902 19966 32954
rect 19966 32902 20018 32954
rect 20018 32902 20020 32954
rect 19964 32900 20020 32902
rect 20068 32954 20124 32956
rect 20068 32902 20070 32954
rect 20070 32902 20122 32954
rect 20122 32902 20124 32954
rect 20068 32900 20124 32902
rect 19860 31386 19916 31388
rect 19860 31334 19862 31386
rect 19862 31334 19914 31386
rect 19914 31334 19916 31386
rect 19860 31332 19916 31334
rect 19964 31386 20020 31388
rect 19964 31334 19966 31386
rect 19966 31334 20018 31386
rect 20018 31334 20020 31386
rect 19964 31332 20020 31334
rect 20068 31386 20124 31388
rect 20068 31334 20070 31386
rect 20070 31334 20122 31386
rect 20122 31334 20124 31386
rect 20068 31332 20124 31334
rect 19860 29818 19916 29820
rect 19860 29766 19862 29818
rect 19862 29766 19914 29818
rect 19914 29766 19916 29818
rect 19860 29764 19916 29766
rect 19964 29818 20020 29820
rect 19964 29766 19966 29818
rect 19966 29766 20018 29818
rect 20018 29766 20020 29818
rect 19964 29764 20020 29766
rect 20068 29818 20124 29820
rect 20068 29766 20070 29818
rect 20070 29766 20122 29818
rect 20122 29766 20124 29818
rect 20068 29764 20124 29766
rect 19964 29538 20020 29540
rect 19964 29486 19966 29538
rect 19966 29486 20018 29538
rect 20018 29486 20020 29538
rect 19964 29484 20020 29486
rect 20300 29260 20356 29316
rect 19860 28250 19916 28252
rect 19860 28198 19862 28250
rect 19862 28198 19914 28250
rect 19914 28198 19916 28250
rect 19860 28196 19916 28198
rect 19964 28250 20020 28252
rect 19964 28198 19966 28250
rect 19966 28198 20018 28250
rect 20018 28198 20020 28250
rect 19964 28196 20020 28198
rect 20068 28250 20124 28252
rect 20068 28198 20070 28250
rect 20070 28198 20122 28250
rect 20122 28198 20124 28250
rect 20068 28196 20124 28198
rect 20524 27970 20580 27972
rect 20524 27918 20526 27970
rect 20526 27918 20578 27970
rect 20578 27918 20580 27970
rect 20524 27916 20580 27918
rect 20188 27692 20244 27748
rect 19740 27244 19796 27300
rect 20412 26796 20468 26852
rect 19860 26682 19916 26684
rect 19860 26630 19862 26682
rect 19862 26630 19914 26682
rect 19914 26630 19916 26682
rect 19860 26628 19916 26630
rect 19964 26682 20020 26684
rect 19964 26630 19966 26682
rect 19966 26630 20018 26682
rect 20018 26630 20020 26682
rect 19964 26628 20020 26630
rect 20068 26682 20124 26684
rect 20068 26630 20070 26682
rect 20070 26630 20122 26682
rect 20122 26630 20124 26682
rect 20068 26628 20124 26630
rect 20076 26348 20132 26404
rect 19740 26290 19796 26292
rect 19740 26238 19742 26290
rect 19742 26238 19794 26290
rect 19794 26238 19796 26290
rect 19740 26236 19796 26238
rect 19852 25788 19908 25844
rect 20076 25452 20132 25508
rect 18956 24722 19012 24724
rect 18956 24670 18958 24722
rect 18958 24670 19010 24722
rect 19010 24670 19012 24722
rect 18956 24668 19012 24670
rect 19180 24498 19236 24500
rect 19180 24446 19182 24498
rect 19182 24446 19234 24498
rect 19234 24446 19236 24498
rect 19180 24444 19236 24446
rect 18172 23884 18228 23940
rect 20300 26012 20356 26068
rect 20188 25340 20244 25396
rect 20076 25282 20132 25284
rect 20076 25230 20078 25282
rect 20078 25230 20130 25282
rect 20130 25230 20132 25282
rect 20076 25228 20132 25230
rect 19860 25114 19916 25116
rect 19860 25062 19862 25114
rect 19862 25062 19914 25114
rect 19914 25062 19916 25114
rect 19860 25060 19916 25062
rect 19964 25114 20020 25116
rect 19964 25062 19966 25114
rect 19966 25062 20018 25114
rect 20018 25062 20020 25114
rect 19964 25060 20020 25062
rect 20068 25114 20124 25116
rect 20068 25062 20070 25114
rect 20070 25062 20122 25114
rect 20122 25062 20124 25114
rect 20068 25060 20124 25062
rect 18956 23660 19012 23716
rect 18172 23266 18228 23268
rect 18172 23214 18174 23266
rect 18174 23214 18226 23266
rect 18226 23214 18228 23266
rect 18172 23212 18228 23214
rect 18284 23100 18340 23156
rect 19292 23548 19348 23604
rect 18620 22988 18676 23044
rect 19180 23042 19236 23044
rect 19180 22990 19182 23042
rect 19182 22990 19234 23042
rect 19234 22990 19236 23042
rect 19180 22988 19236 22990
rect 18956 22930 19012 22932
rect 18956 22878 18958 22930
rect 18958 22878 19010 22930
rect 19010 22878 19012 22930
rect 18956 22876 19012 22878
rect 18732 22092 18788 22148
rect 18060 21980 18116 22036
rect 20188 24556 20244 24612
rect 21196 29202 21252 29204
rect 21196 29150 21198 29202
rect 21198 29150 21250 29202
rect 21250 29150 21252 29202
rect 21196 29148 21252 29150
rect 20972 27916 21028 27972
rect 21308 26290 21364 26292
rect 21308 26238 21310 26290
rect 21310 26238 21362 26290
rect 21362 26238 21364 26290
rect 21308 26236 21364 26238
rect 21196 26124 21252 26180
rect 19860 23546 19916 23548
rect 19860 23494 19862 23546
rect 19862 23494 19914 23546
rect 19914 23494 19916 23546
rect 19860 23492 19916 23494
rect 19964 23546 20020 23548
rect 19964 23494 19966 23546
rect 19966 23494 20018 23546
rect 20018 23494 20020 23546
rect 19964 23492 20020 23494
rect 20068 23546 20124 23548
rect 20068 23494 20070 23546
rect 20070 23494 20122 23546
rect 20122 23494 20124 23546
rect 20068 23492 20124 23494
rect 19404 23154 19460 23156
rect 19404 23102 19406 23154
rect 19406 23102 19458 23154
rect 19458 23102 19460 23154
rect 19404 23100 19460 23102
rect 19628 23324 19684 23380
rect 19964 23266 20020 23268
rect 19964 23214 19966 23266
rect 19966 23214 20018 23266
rect 20018 23214 20020 23266
rect 19964 23212 20020 23214
rect 20076 22146 20132 22148
rect 20076 22094 20078 22146
rect 20078 22094 20130 22146
rect 20130 22094 20132 22146
rect 20076 22092 20132 22094
rect 19860 21978 19916 21980
rect 19860 21926 19862 21978
rect 19862 21926 19914 21978
rect 19914 21926 19916 21978
rect 19860 21924 19916 21926
rect 19964 21978 20020 21980
rect 19964 21926 19966 21978
rect 19966 21926 20018 21978
rect 20018 21926 20020 21978
rect 19964 21924 20020 21926
rect 20068 21978 20124 21980
rect 20068 21926 20070 21978
rect 20070 21926 20122 21978
rect 20122 21926 20124 21978
rect 20068 21924 20124 21926
rect 17724 20914 17780 20916
rect 17724 20862 17726 20914
rect 17726 20862 17778 20914
rect 17778 20862 17780 20914
rect 17724 20860 17780 20862
rect 17500 20130 17556 20132
rect 17500 20078 17502 20130
rect 17502 20078 17554 20130
rect 17554 20078 17556 20130
rect 17500 20076 17556 20078
rect 17612 20188 17668 20244
rect 17276 18508 17332 18564
rect 17052 17500 17108 17556
rect 17836 20130 17892 20132
rect 17836 20078 17838 20130
rect 17838 20078 17890 20130
rect 17890 20078 17892 20130
rect 17836 20076 17892 20078
rect 17948 19964 18004 20020
rect 17836 19068 17892 19124
rect 18284 21308 18340 21364
rect 18508 20690 18564 20692
rect 18508 20638 18510 20690
rect 18510 20638 18562 20690
rect 18562 20638 18564 20690
rect 18508 20636 18564 20638
rect 18508 20188 18564 20244
rect 18732 20018 18788 20020
rect 18732 19966 18734 20018
rect 18734 19966 18786 20018
rect 18786 19966 18788 20018
rect 18732 19964 18788 19966
rect 18172 19180 18228 19236
rect 18396 18450 18452 18452
rect 18396 18398 18398 18450
rect 18398 18398 18450 18450
rect 18450 18398 18452 18450
rect 18396 18396 18452 18398
rect 18844 19234 18900 19236
rect 18844 19182 18846 19234
rect 18846 19182 18898 19234
rect 18898 19182 18900 19234
rect 18844 19180 18900 19182
rect 20972 24556 21028 24612
rect 22092 36370 22148 36372
rect 22092 36318 22094 36370
rect 22094 36318 22146 36370
rect 22146 36318 22148 36370
rect 22092 36316 22148 36318
rect 22428 35420 22484 35476
rect 21756 33068 21812 33124
rect 24522 36874 24578 36876
rect 24522 36822 24524 36874
rect 24524 36822 24576 36874
rect 24576 36822 24578 36874
rect 24522 36820 24578 36822
rect 24626 36874 24682 36876
rect 24626 36822 24628 36874
rect 24628 36822 24680 36874
rect 24680 36822 24682 36874
rect 24626 36820 24682 36822
rect 24730 36874 24786 36876
rect 24730 36822 24732 36874
rect 24732 36822 24784 36874
rect 24784 36822 24786 36874
rect 24892 36876 24948 36932
rect 25900 36876 25956 36932
rect 24730 36820 24786 36822
rect 24220 36652 24276 36708
rect 25228 36652 25284 36708
rect 22652 33068 22708 33124
rect 21980 29596 22036 29652
rect 22428 29426 22484 29428
rect 22428 29374 22430 29426
rect 22430 29374 22482 29426
rect 22482 29374 22484 29426
rect 22428 29372 22484 29374
rect 21868 29260 21924 29316
rect 22764 29314 22820 29316
rect 22764 29262 22766 29314
rect 22766 29262 22818 29314
rect 22818 29262 22820 29314
rect 22764 29260 22820 29262
rect 22204 29202 22260 29204
rect 22204 29150 22206 29202
rect 22206 29150 22258 29202
rect 22258 29150 22260 29202
rect 22204 29148 22260 29150
rect 22988 29202 23044 29204
rect 22988 29150 22990 29202
rect 22990 29150 23042 29202
rect 23042 29150 23044 29202
rect 22988 29148 23044 29150
rect 21980 27916 22036 27972
rect 22652 27804 22708 27860
rect 22316 27074 22372 27076
rect 22316 27022 22318 27074
rect 22318 27022 22370 27074
rect 22370 27022 22372 27074
rect 22316 27020 22372 27022
rect 23548 36316 23604 36372
rect 23436 33852 23492 33908
rect 23212 28028 23268 28084
rect 23324 28476 23380 28532
rect 21980 26402 22036 26404
rect 21980 26350 21982 26402
rect 21982 26350 22034 26402
rect 22034 26350 22036 26402
rect 21980 26348 22036 26350
rect 21420 26012 21476 26068
rect 21420 25788 21476 25844
rect 21308 25394 21364 25396
rect 21308 25342 21310 25394
rect 21310 25342 21362 25394
rect 21362 25342 21364 25394
rect 21308 25340 21364 25342
rect 21196 24444 21252 24500
rect 21196 23884 21252 23940
rect 20300 23266 20356 23268
rect 20300 23214 20302 23266
rect 20302 23214 20354 23266
rect 20354 23214 20356 23266
rect 20300 23212 20356 23214
rect 20412 22092 20468 22148
rect 20300 21698 20356 21700
rect 20300 21646 20302 21698
rect 20302 21646 20354 21698
rect 20354 21646 20356 21698
rect 20300 21644 20356 21646
rect 20636 22204 20692 22260
rect 21980 24444 22036 24500
rect 21644 23826 21700 23828
rect 21644 23774 21646 23826
rect 21646 23774 21698 23826
rect 21698 23774 21700 23826
rect 21644 23772 21700 23774
rect 22204 23996 22260 24052
rect 23996 35532 24052 35588
rect 23660 33068 23716 33124
rect 23884 29202 23940 29204
rect 23884 29150 23886 29202
rect 23886 29150 23938 29202
rect 23938 29150 23940 29202
rect 23884 29148 23940 29150
rect 24522 35306 24578 35308
rect 24522 35254 24524 35306
rect 24524 35254 24576 35306
rect 24576 35254 24578 35306
rect 24522 35252 24578 35254
rect 24626 35306 24682 35308
rect 24626 35254 24628 35306
rect 24628 35254 24680 35306
rect 24680 35254 24682 35306
rect 24626 35252 24682 35254
rect 24730 35306 24786 35308
rect 24730 35254 24732 35306
rect 24732 35254 24784 35306
rect 24784 35254 24786 35306
rect 24730 35252 24786 35254
rect 24892 33852 24948 33908
rect 25004 35868 25060 35924
rect 24522 33738 24578 33740
rect 24522 33686 24524 33738
rect 24524 33686 24576 33738
rect 24576 33686 24578 33738
rect 24522 33684 24578 33686
rect 24626 33738 24682 33740
rect 24626 33686 24628 33738
rect 24628 33686 24680 33738
rect 24680 33686 24682 33738
rect 24626 33684 24682 33686
rect 24730 33738 24786 33740
rect 24730 33686 24732 33738
rect 24732 33686 24784 33738
rect 24784 33686 24786 33738
rect 24730 33684 24786 33686
rect 24522 32170 24578 32172
rect 24522 32118 24524 32170
rect 24524 32118 24576 32170
rect 24576 32118 24578 32170
rect 24522 32116 24578 32118
rect 24626 32170 24682 32172
rect 24626 32118 24628 32170
rect 24628 32118 24680 32170
rect 24680 32118 24682 32170
rect 24626 32116 24682 32118
rect 24730 32170 24786 32172
rect 24730 32118 24732 32170
rect 24732 32118 24784 32170
rect 24784 32118 24786 32170
rect 24730 32116 24786 32118
rect 24522 30602 24578 30604
rect 24522 30550 24524 30602
rect 24524 30550 24576 30602
rect 24576 30550 24578 30602
rect 24522 30548 24578 30550
rect 24626 30602 24682 30604
rect 24626 30550 24628 30602
rect 24628 30550 24680 30602
rect 24680 30550 24682 30602
rect 24626 30548 24682 30550
rect 24730 30602 24786 30604
rect 24730 30550 24732 30602
rect 24732 30550 24784 30602
rect 24784 30550 24786 30602
rect 24730 30548 24786 30550
rect 24332 30380 24388 30436
rect 24522 29034 24578 29036
rect 24522 28982 24524 29034
rect 24524 28982 24576 29034
rect 24576 28982 24578 29034
rect 24522 28980 24578 28982
rect 24626 29034 24682 29036
rect 24626 28982 24628 29034
rect 24628 28982 24680 29034
rect 24680 28982 24682 29034
rect 24626 28980 24682 28982
rect 24730 29034 24786 29036
rect 24730 28982 24732 29034
rect 24732 28982 24784 29034
rect 24784 28982 24786 29034
rect 24730 28980 24786 28982
rect 26236 36876 26292 36932
rect 26236 36370 26292 36372
rect 26236 36318 26238 36370
rect 26238 36318 26290 36370
rect 26290 36318 26292 36370
rect 26236 36316 26292 36318
rect 26796 36204 26852 36260
rect 25452 33068 25508 33124
rect 25788 33516 25844 33572
rect 26124 29708 26180 29764
rect 25452 29202 25508 29204
rect 25452 29150 25454 29202
rect 25454 29150 25506 29202
rect 25506 29150 25508 29202
rect 25452 29148 25508 29150
rect 23884 27858 23940 27860
rect 23884 27806 23886 27858
rect 23886 27806 23938 27858
rect 23938 27806 23940 27858
rect 23884 27804 23940 27806
rect 24108 27804 24164 27860
rect 23660 26348 23716 26404
rect 24108 27020 24164 27076
rect 23772 26290 23828 26292
rect 23772 26238 23774 26290
rect 23774 26238 23826 26290
rect 23826 26238 23828 26290
rect 23772 26236 23828 26238
rect 22764 25730 22820 25732
rect 22764 25678 22766 25730
rect 22766 25678 22818 25730
rect 22818 25678 22820 25730
rect 22764 25676 22820 25678
rect 23324 25730 23380 25732
rect 23324 25678 23326 25730
rect 23326 25678 23378 25730
rect 23378 25678 23380 25730
rect 23324 25676 23380 25678
rect 22428 25116 22484 25172
rect 22876 25116 22932 25172
rect 22428 24946 22484 24948
rect 22428 24894 22430 24946
rect 22430 24894 22482 24946
rect 22482 24894 22484 24946
rect 22428 24892 22484 24894
rect 22876 24332 22932 24388
rect 22316 23548 22372 23604
rect 22652 23714 22708 23716
rect 22652 23662 22654 23714
rect 22654 23662 22706 23714
rect 22706 23662 22708 23714
rect 22652 23660 22708 23662
rect 20972 21308 21028 21364
rect 19860 20410 19916 20412
rect 19860 20358 19862 20410
rect 19862 20358 19914 20410
rect 19914 20358 19916 20410
rect 19860 20356 19916 20358
rect 19964 20410 20020 20412
rect 19964 20358 19966 20410
rect 19966 20358 20018 20410
rect 20018 20358 20020 20410
rect 19964 20356 20020 20358
rect 20068 20410 20124 20412
rect 20068 20358 20070 20410
rect 20070 20358 20122 20410
rect 20122 20358 20124 20410
rect 20068 20356 20124 20358
rect 19852 20242 19908 20244
rect 19852 20190 19854 20242
rect 19854 20190 19906 20242
rect 19906 20190 19908 20242
rect 19852 20188 19908 20190
rect 19068 20076 19124 20132
rect 19292 19852 19348 19908
rect 19180 19068 19236 19124
rect 18844 18284 18900 18340
rect 18956 18450 19012 18452
rect 18956 18398 18958 18450
rect 18958 18398 19010 18450
rect 19010 18398 19012 18450
rect 18956 18396 19012 18398
rect 18284 17724 18340 17780
rect 17388 17052 17444 17108
rect 17612 17052 17668 17108
rect 16492 15708 16548 15764
rect 16044 15260 16100 15316
rect 17052 16380 17108 16436
rect 16940 15986 16996 15988
rect 16940 15934 16942 15986
rect 16942 15934 16994 15986
rect 16994 15934 16996 15986
rect 16940 15932 16996 15934
rect 16716 15708 16772 15764
rect 16044 14140 16100 14196
rect 16380 13916 16436 13972
rect 16156 13746 16212 13748
rect 16156 13694 16158 13746
rect 16158 13694 16210 13746
rect 16210 13694 16212 13746
rect 16156 13692 16212 13694
rect 15932 13356 15988 13412
rect 16156 13186 16212 13188
rect 16156 13134 16158 13186
rect 16158 13134 16210 13186
rect 16210 13134 16212 13186
rect 16156 13132 16212 13134
rect 15596 13020 15652 13076
rect 16044 13074 16100 13076
rect 16044 13022 16046 13074
rect 16046 13022 16098 13074
rect 16098 13022 16100 13074
rect 16044 13020 16100 13022
rect 15820 12962 15876 12964
rect 15820 12910 15822 12962
rect 15822 12910 15874 12962
rect 15874 12910 15876 12962
rect 15820 12908 15876 12910
rect 16828 15538 16884 15540
rect 16828 15486 16830 15538
rect 16830 15486 16882 15538
rect 16882 15486 16884 15538
rect 16828 15484 16884 15486
rect 16940 14028 16996 14084
rect 17276 16604 17332 16660
rect 17388 16380 17444 16436
rect 18172 17164 18228 17220
rect 17724 16604 17780 16660
rect 17612 16492 17668 16548
rect 18396 17388 18452 17444
rect 18956 16940 19012 16996
rect 20524 19906 20580 19908
rect 20524 19854 20526 19906
rect 20526 19854 20578 19906
rect 20578 19854 20580 19906
rect 20524 19852 20580 19854
rect 20524 19122 20580 19124
rect 20524 19070 20526 19122
rect 20526 19070 20578 19122
rect 20578 19070 20580 19122
rect 20524 19068 20580 19070
rect 20076 19010 20132 19012
rect 20076 18958 20078 19010
rect 20078 18958 20130 19010
rect 20130 18958 20132 19010
rect 20076 18956 20132 18958
rect 20748 18956 20804 19012
rect 19860 18842 19916 18844
rect 19860 18790 19862 18842
rect 19862 18790 19914 18842
rect 19914 18790 19916 18842
rect 19860 18788 19916 18790
rect 19964 18842 20020 18844
rect 19964 18790 19966 18842
rect 19966 18790 20018 18842
rect 20018 18790 20020 18842
rect 19964 18788 20020 18790
rect 20068 18842 20124 18844
rect 20068 18790 20070 18842
rect 20070 18790 20122 18842
rect 20122 18790 20124 18842
rect 20068 18788 20124 18790
rect 20188 18674 20244 18676
rect 20188 18622 20190 18674
rect 20190 18622 20242 18674
rect 20242 18622 20244 18674
rect 20188 18620 20244 18622
rect 19964 18508 20020 18564
rect 19404 18396 19460 18452
rect 19516 18338 19572 18340
rect 19516 18286 19518 18338
rect 19518 18286 19570 18338
rect 19570 18286 19572 18338
rect 19516 18284 19572 18286
rect 19404 17778 19460 17780
rect 19404 17726 19406 17778
rect 19406 17726 19458 17778
rect 19458 17726 19460 17778
rect 19404 17724 19460 17726
rect 17836 15932 17892 15988
rect 17276 14588 17332 14644
rect 17612 15426 17668 15428
rect 17612 15374 17614 15426
rect 17614 15374 17666 15426
rect 17666 15374 17668 15426
rect 17612 15372 17668 15374
rect 17164 14140 17220 14196
rect 17052 13916 17108 13972
rect 17276 14028 17332 14084
rect 16492 12908 16548 12964
rect 15260 12066 15316 12068
rect 15260 12014 15262 12066
rect 15262 12014 15314 12066
rect 15314 12014 15316 12066
rect 15260 12012 15316 12014
rect 16268 12796 16324 12852
rect 16828 12850 16884 12852
rect 16828 12798 16830 12850
rect 16830 12798 16882 12850
rect 16882 12798 16884 12850
rect 16828 12796 16884 12798
rect 15820 12066 15876 12068
rect 15820 12014 15822 12066
rect 15822 12014 15874 12066
rect 15874 12014 15876 12066
rect 15820 12012 15876 12014
rect 15708 11900 15764 11956
rect 15198 11786 15254 11788
rect 15198 11734 15200 11786
rect 15200 11734 15252 11786
rect 15252 11734 15254 11786
rect 15198 11732 15254 11734
rect 15302 11786 15358 11788
rect 15302 11734 15304 11786
rect 15304 11734 15356 11786
rect 15356 11734 15358 11786
rect 15302 11732 15358 11734
rect 15406 11786 15462 11788
rect 15406 11734 15408 11786
rect 15408 11734 15460 11786
rect 15460 11734 15462 11786
rect 15406 11732 15462 11734
rect 14924 11452 14980 11508
rect 16044 11452 16100 11508
rect 15036 11170 15092 11172
rect 15036 11118 15038 11170
rect 15038 11118 15090 11170
rect 15090 11118 15092 11170
rect 15036 11116 15092 11118
rect 15484 11170 15540 11172
rect 15484 11118 15486 11170
rect 15486 11118 15538 11170
rect 15538 11118 15540 11170
rect 15484 11116 15540 11118
rect 15484 10780 15540 10836
rect 16156 10780 16212 10836
rect 17052 12962 17108 12964
rect 17052 12910 17054 12962
rect 17054 12910 17106 12962
rect 17106 12910 17108 12962
rect 17052 12908 17108 12910
rect 17052 12684 17108 12740
rect 16716 11394 16772 11396
rect 16716 11342 16718 11394
rect 16718 11342 16770 11394
rect 16770 11342 16772 11394
rect 16716 11340 16772 11342
rect 17948 15484 18004 15540
rect 18620 16156 18676 16212
rect 18172 15820 18228 15876
rect 18396 15314 18452 15316
rect 18396 15262 18398 15314
rect 18398 15262 18450 15314
rect 18450 15262 18452 15314
rect 18396 15260 18452 15262
rect 17836 14588 17892 14644
rect 17724 14418 17780 14420
rect 17724 14366 17726 14418
rect 17726 14366 17778 14418
rect 17778 14366 17780 14418
rect 17724 14364 17780 14366
rect 17500 14306 17556 14308
rect 17500 14254 17502 14306
rect 17502 14254 17554 14306
rect 17554 14254 17556 14306
rect 17500 14252 17556 14254
rect 17500 14028 17556 14084
rect 17948 14476 18004 14532
rect 18508 14530 18564 14532
rect 18508 14478 18510 14530
rect 18510 14478 18562 14530
rect 18562 14478 18564 14530
rect 18508 14476 18564 14478
rect 18060 14418 18116 14420
rect 18060 14366 18062 14418
rect 18062 14366 18114 14418
rect 18114 14366 18116 14418
rect 18060 14364 18116 14366
rect 18844 15314 18900 15316
rect 18844 15262 18846 15314
rect 18846 15262 18898 15314
rect 18898 15262 18900 15314
rect 18844 15260 18900 15262
rect 19516 16268 19572 16324
rect 18956 15148 19012 15204
rect 19860 17274 19916 17276
rect 19860 17222 19862 17274
rect 19862 17222 19914 17274
rect 19914 17222 19916 17274
rect 19860 17220 19916 17222
rect 19964 17274 20020 17276
rect 19964 17222 19966 17274
rect 19966 17222 20018 17274
rect 20018 17222 20020 17274
rect 19964 17220 20020 17222
rect 20068 17274 20124 17276
rect 20068 17222 20070 17274
rect 20070 17222 20122 17274
rect 20122 17222 20124 17274
rect 20068 17220 20124 17222
rect 19964 16994 20020 16996
rect 19964 16942 19966 16994
rect 19966 16942 20018 16994
rect 20018 16942 20020 16994
rect 19964 16940 20020 16942
rect 18844 14700 18900 14756
rect 19180 15260 19236 15316
rect 19628 14364 19684 14420
rect 19180 14252 19236 14308
rect 19628 14140 19684 14196
rect 17724 13692 17780 13748
rect 17500 13580 17556 13636
rect 17724 12962 17780 12964
rect 17724 12910 17726 12962
rect 17726 12910 17778 12962
rect 17778 12910 17780 12962
rect 17724 12908 17780 12910
rect 17500 12796 17556 12852
rect 17500 12402 17556 12404
rect 17500 12350 17502 12402
rect 17502 12350 17554 12402
rect 17554 12350 17556 12402
rect 17500 12348 17556 12350
rect 17276 11452 17332 11508
rect 16380 11282 16436 11284
rect 16380 11230 16382 11282
rect 16382 11230 16434 11282
rect 16434 11230 16436 11282
rect 16380 11228 16436 11230
rect 16940 11170 16996 11172
rect 16940 11118 16942 11170
rect 16942 11118 16994 11170
rect 16994 11118 16996 11170
rect 16940 11116 16996 11118
rect 16268 11004 16324 11060
rect 17948 12850 18004 12852
rect 17948 12798 17950 12850
rect 17950 12798 18002 12850
rect 18002 12798 18004 12850
rect 17948 12796 18004 12798
rect 17724 12348 17780 12404
rect 17724 11394 17780 11396
rect 17724 11342 17726 11394
rect 17726 11342 17778 11394
rect 17778 11342 17780 11394
rect 17724 11340 17780 11342
rect 17612 11282 17668 11284
rect 17612 11230 17614 11282
rect 17614 11230 17666 11282
rect 17666 11230 17668 11282
rect 17612 11228 17668 11230
rect 18396 11282 18452 11284
rect 18396 11230 18398 11282
rect 18398 11230 18450 11282
rect 18450 11230 18452 11282
rect 18396 11228 18452 11230
rect 17276 11004 17332 11060
rect 16716 10668 16772 10724
rect 15198 10218 15254 10220
rect 15198 10166 15200 10218
rect 15200 10166 15252 10218
rect 15252 10166 15254 10218
rect 15198 10164 15254 10166
rect 15302 10218 15358 10220
rect 15302 10166 15304 10218
rect 15304 10166 15356 10218
rect 15356 10166 15358 10218
rect 15302 10164 15358 10166
rect 15406 10218 15462 10220
rect 15406 10166 15408 10218
rect 15408 10166 15460 10218
rect 15460 10166 15462 10218
rect 15406 10164 15462 10166
rect 15198 8650 15254 8652
rect 15198 8598 15200 8650
rect 15200 8598 15252 8650
rect 15252 8598 15254 8650
rect 15198 8596 15254 8598
rect 15302 8650 15358 8652
rect 15302 8598 15304 8650
rect 15304 8598 15356 8650
rect 15356 8598 15358 8650
rect 15302 8596 15358 8598
rect 15406 8650 15462 8652
rect 15406 8598 15408 8650
rect 15408 8598 15460 8650
rect 15460 8598 15462 8650
rect 15406 8596 15462 8598
rect 15198 7082 15254 7084
rect 15198 7030 15200 7082
rect 15200 7030 15252 7082
rect 15252 7030 15254 7082
rect 15198 7028 15254 7030
rect 15302 7082 15358 7084
rect 15302 7030 15304 7082
rect 15304 7030 15356 7082
rect 15356 7030 15358 7082
rect 15302 7028 15358 7030
rect 15406 7082 15462 7084
rect 15406 7030 15408 7082
rect 15408 7030 15460 7082
rect 15460 7030 15462 7082
rect 15406 7028 15462 7030
rect 15198 5514 15254 5516
rect 15198 5462 15200 5514
rect 15200 5462 15252 5514
rect 15252 5462 15254 5514
rect 15198 5460 15254 5462
rect 15302 5514 15358 5516
rect 15302 5462 15304 5514
rect 15304 5462 15356 5514
rect 15356 5462 15358 5514
rect 15302 5460 15358 5462
rect 15406 5514 15462 5516
rect 15406 5462 15408 5514
rect 15408 5462 15460 5514
rect 15460 5462 15462 5514
rect 15406 5460 15462 5462
rect 15198 3946 15254 3948
rect 15198 3894 15200 3946
rect 15200 3894 15252 3946
rect 15252 3894 15254 3946
rect 15198 3892 15254 3894
rect 15302 3946 15358 3948
rect 15302 3894 15304 3946
rect 15304 3894 15356 3946
rect 15356 3894 15358 3946
rect 15302 3892 15358 3894
rect 15406 3946 15462 3948
rect 15406 3894 15408 3946
rect 15408 3894 15460 3946
rect 15460 3894 15462 3946
rect 15406 3892 15462 3894
rect 16044 3554 16100 3556
rect 16044 3502 16046 3554
rect 16046 3502 16098 3554
rect 16098 3502 16100 3554
rect 16044 3500 16100 3502
rect 18732 10722 18788 10724
rect 18732 10670 18734 10722
rect 18734 10670 18786 10722
rect 18786 10670 18788 10722
rect 18732 10668 18788 10670
rect 18732 9100 18788 9156
rect 18956 11116 19012 11172
rect 19068 11004 19124 11060
rect 18956 10108 19012 10164
rect 18956 7474 19012 7476
rect 18956 7422 18958 7474
rect 18958 7422 19010 7474
rect 19010 7422 19012 7474
rect 18956 7420 19012 7422
rect 19516 13970 19572 13972
rect 19516 13918 19518 13970
rect 19518 13918 19570 13970
rect 19570 13918 19572 13970
rect 19516 13916 19572 13918
rect 19404 11564 19460 11620
rect 19404 10780 19460 10836
rect 20636 16716 20692 16772
rect 20636 16044 20692 16100
rect 19860 15706 19916 15708
rect 19860 15654 19862 15706
rect 19862 15654 19914 15706
rect 19914 15654 19916 15706
rect 19860 15652 19916 15654
rect 19964 15706 20020 15708
rect 19964 15654 19966 15706
rect 19966 15654 20018 15706
rect 20018 15654 20020 15706
rect 19964 15652 20020 15654
rect 20068 15706 20124 15708
rect 20068 15654 20070 15706
rect 20070 15654 20122 15706
rect 20122 15654 20124 15706
rect 20068 15652 20124 15654
rect 20188 15148 20244 15204
rect 20524 15596 20580 15652
rect 21308 21698 21364 21700
rect 21308 21646 21310 21698
rect 21310 21646 21362 21698
rect 21362 21646 21364 21698
rect 21308 21644 21364 21646
rect 22428 22370 22484 22372
rect 22428 22318 22430 22370
rect 22430 22318 22482 22370
rect 22482 22318 22484 22370
rect 22428 22316 22484 22318
rect 22540 22258 22596 22260
rect 22540 22206 22542 22258
rect 22542 22206 22594 22258
rect 22594 22206 22596 22258
rect 22540 22204 22596 22206
rect 22988 23826 23044 23828
rect 22988 23774 22990 23826
rect 22990 23774 23042 23826
rect 23042 23774 23044 23826
rect 22988 23772 23044 23774
rect 21644 21532 21700 21588
rect 22876 21532 22932 21588
rect 21308 20690 21364 20692
rect 21308 20638 21310 20690
rect 21310 20638 21362 20690
rect 21362 20638 21364 20690
rect 21308 20636 21364 20638
rect 21644 20578 21700 20580
rect 21644 20526 21646 20578
rect 21646 20526 21698 20578
rect 21698 20526 21700 20578
rect 21644 20524 21700 20526
rect 21308 20188 21364 20244
rect 21196 20130 21252 20132
rect 21196 20078 21198 20130
rect 21198 20078 21250 20130
rect 21250 20078 21252 20130
rect 21196 20076 21252 20078
rect 21644 19964 21700 20020
rect 22764 20690 22820 20692
rect 22764 20638 22766 20690
rect 22766 20638 22818 20690
rect 22818 20638 22820 20690
rect 22764 20636 22820 20638
rect 22316 19964 22372 20020
rect 21980 19852 22036 19908
rect 23324 23996 23380 24052
rect 23100 23660 23156 23716
rect 23212 23548 23268 23604
rect 23548 23548 23604 23604
rect 23772 23266 23828 23268
rect 23772 23214 23774 23266
rect 23774 23214 23826 23266
rect 23826 23214 23828 23266
rect 23772 23212 23828 23214
rect 22540 19740 22596 19796
rect 20860 18620 20916 18676
rect 21084 18338 21140 18340
rect 21084 18286 21086 18338
rect 21086 18286 21138 18338
rect 21138 18286 21140 18338
rect 21084 18284 21140 18286
rect 22652 19404 22708 19460
rect 21756 17666 21812 17668
rect 21756 17614 21758 17666
rect 21758 17614 21810 17666
rect 21810 17614 21812 17666
rect 21756 17612 21812 17614
rect 21532 16940 21588 16996
rect 21980 16994 22036 16996
rect 21980 16942 21982 16994
rect 21982 16942 22034 16994
rect 22034 16942 22036 16994
rect 21980 16940 22036 16942
rect 20972 15148 21028 15204
rect 20188 14530 20244 14532
rect 20188 14478 20190 14530
rect 20190 14478 20242 14530
rect 20242 14478 20244 14530
rect 20188 14476 20244 14478
rect 19860 14138 19916 14140
rect 19860 14086 19862 14138
rect 19862 14086 19914 14138
rect 19914 14086 19916 14138
rect 19860 14084 19916 14086
rect 19964 14138 20020 14140
rect 19964 14086 19966 14138
rect 19966 14086 20018 14138
rect 20018 14086 20020 14138
rect 19964 14084 20020 14086
rect 20068 14138 20124 14140
rect 20068 14086 20070 14138
rect 20070 14086 20122 14138
rect 20122 14086 20124 14138
rect 20068 14084 20124 14086
rect 20524 14364 20580 14420
rect 19516 9100 19572 9156
rect 20412 12962 20468 12964
rect 20412 12910 20414 12962
rect 20414 12910 20466 12962
rect 20466 12910 20468 12962
rect 20412 12908 20468 12910
rect 20748 12908 20804 12964
rect 19740 12738 19796 12740
rect 19740 12686 19742 12738
rect 19742 12686 19794 12738
rect 19794 12686 19796 12738
rect 19740 12684 19796 12686
rect 20188 12684 20244 12740
rect 19860 12570 19916 12572
rect 19860 12518 19862 12570
rect 19862 12518 19914 12570
rect 19914 12518 19916 12570
rect 19860 12516 19916 12518
rect 19964 12570 20020 12572
rect 19964 12518 19966 12570
rect 19966 12518 20018 12570
rect 20018 12518 20020 12570
rect 19964 12516 20020 12518
rect 20068 12570 20124 12572
rect 20068 12518 20070 12570
rect 20070 12518 20122 12570
rect 20122 12518 20124 12570
rect 20068 12516 20124 12518
rect 20076 12124 20132 12180
rect 20412 11340 20468 11396
rect 19860 11002 19916 11004
rect 19860 10950 19862 11002
rect 19862 10950 19914 11002
rect 19914 10950 19916 11002
rect 19860 10948 19916 10950
rect 19964 11002 20020 11004
rect 19964 10950 19966 11002
rect 19966 10950 20018 11002
rect 20018 10950 20020 11002
rect 19964 10948 20020 10950
rect 20068 11002 20124 11004
rect 20068 10950 20070 11002
rect 20070 10950 20122 11002
rect 20122 10950 20124 11002
rect 20068 10948 20124 10950
rect 19740 10780 19796 10836
rect 20636 10668 20692 10724
rect 20524 9714 20580 9716
rect 20524 9662 20526 9714
rect 20526 9662 20578 9714
rect 20578 9662 20580 9714
rect 20524 9660 20580 9662
rect 20748 10220 20804 10276
rect 21196 15314 21252 15316
rect 21196 15262 21198 15314
rect 21198 15262 21250 15314
rect 21250 15262 21252 15314
rect 21196 15260 21252 15262
rect 21868 16828 21924 16884
rect 21420 15820 21476 15876
rect 21644 15260 21700 15316
rect 21756 15148 21812 15204
rect 20972 14252 21028 14308
rect 20972 12684 21028 12740
rect 21308 14530 21364 14532
rect 21308 14478 21310 14530
rect 21310 14478 21362 14530
rect 21362 14478 21364 14530
rect 21308 14476 21364 14478
rect 21980 15874 22036 15876
rect 21980 15822 21982 15874
rect 21982 15822 22034 15874
rect 22034 15822 22036 15874
rect 21980 15820 22036 15822
rect 21980 14364 22036 14420
rect 21868 14306 21924 14308
rect 21868 14254 21870 14306
rect 21870 14254 21922 14306
rect 21922 14254 21924 14306
rect 21868 14252 21924 14254
rect 22988 20130 23044 20132
rect 22988 20078 22990 20130
rect 22990 20078 23042 20130
rect 23042 20078 23044 20130
rect 22988 20076 23044 20078
rect 23212 22316 23268 22372
rect 23548 22316 23604 22372
rect 24108 25676 24164 25732
rect 24220 26460 24276 26516
rect 24780 28476 24836 28532
rect 24522 27466 24578 27468
rect 24522 27414 24524 27466
rect 24524 27414 24576 27466
rect 24576 27414 24578 27466
rect 24522 27412 24578 27414
rect 24626 27466 24682 27468
rect 24626 27414 24628 27466
rect 24628 27414 24680 27466
rect 24680 27414 24682 27466
rect 24626 27412 24682 27414
rect 24730 27466 24786 27468
rect 24730 27414 24732 27466
rect 24732 27414 24784 27466
rect 24784 27414 24786 27466
rect 24730 27412 24786 27414
rect 24668 27074 24724 27076
rect 24668 27022 24670 27074
rect 24670 27022 24722 27074
rect 24722 27022 24724 27074
rect 24668 27020 24724 27022
rect 25452 27970 25508 27972
rect 25452 27918 25454 27970
rect 25454 27918 25506 27970
rect 25506 27918 25508 27970
rect 25452 27916 25508 27918
rect 25900 28476 25956 28532
rect 25340 27858 25396 27860
rect 25340 27806 25342 27858
rect 25342 27806 25394 27858
rect 25394 27806 25396 27858
rect 25340 27804 25396 27806
rect 25340 27020 25396 27076
rect 24892 26348 24948 26404
rect 24522 25898 24578 25900
rect 24522 25846 24524 25898
rect 24524 25846 24576 25898
rect 24576 25846 24578 25898
rect 24522 25844 24578 25846
rect 24626 25898 24682 25900
rect 24626 25846 24628 25898
rect 24628 25846 24680 25898
rect 24680 25846 24682 25898
rect 24626 25844 24682 25846
rect 24730 25898 24786 25900
rect 24730 25846 24732 25898
rect 24732 25846 24784 25898
rect 24784 25846 24786 25898
rect 24730 25844 24786 25846
rect 24444 25506 24500 25508
rect 24444 25454 24446 25506
rect 24446 25454 24498 25506
rect 24498 25454 24500 25506
rect 24444 25452 24500 25454
rect 26460 33628 26516 33684
rect 26348 32508 26404 32564
rect 27244 36876 27300 36932
rect 27468 36482 27524 36484
rect 27468 36430 27470 36482
rect 27470 36430 27522 36482
rect 27522 36430 27524 36482
rect 27468 36428 27524 36430
rect 27692 36316 27748 36372
rect 27356 33516 27412 33572
rect 27580 35308 27636 35364
rect 26796 29708 26852 29764
rect 28700 36370 28756 36372
rect 28700 36318 28702 36370
rect 28702 36318 28754 36370
rect 28754 36318 28756 36370
rect 28700 36316 28756 36318
rect 28476 36204 28532 36260
rect 28252 33516 28308 33572
rect 28812 30940 28868 30996
rect 26572 29314 26628 29316
rect 26572 29262 26574 29314
rect 26574 29262 26626 29314
rect 26626 29262 26628 29314
rect 26572 29260 26628 29262
rect 26796 29202 26852 29204
rect 26796 29150 26798 29202
rect 26798 29150 26850 29202
rect 26850 29150 26852 29202
rect 26796 29148 26852 29150
rect 26460 27858 26516 27860
rect 26460 27806 26462 27858
rect 26462 27806 26514 27858
rect 26514 27806 26516 27858
rect 26460 27804 26516 27806
rect 26684 27858 26740 27860
rect 26684 27806 26686 27858
rect 26686 27806 26738 27858
rect 26738 27806 26740 27858
rect 26684 27804 26740 27806
rect 26460 27020 26516 27076
rect 27468 29314 27524 29316
rect 27468 29262 27470 29314
rect 27470 29262 27522 29314
rect 27522 29262 27524 29314
rect 27468 29260 27524 29262
rect 27356 29148 27412 29204
rect 27692 29202 27748 29204
rect 27692 29150 27694 29202
rect 27694 29150 27746 29202
rect 27746 29150 27748 29202
rect 27692 29148 27748 29150
rect 24668 24834 24724 24836
rect 24668 24782 24670 24834
rect 24670 24782 24722 24834
rect 24722 24782 24724 24834
rect 24668 24780 24724 24782
rect 24444 24722 24500 24724
rect 24444 24670 24446 24722
rect 24446 24670 24498 24722
rect 24498 24670 24500 24722
rect 24444 24668 24500 24670
rect 25228 24722 25284 24724
rect 25228 24670 25230 24722
rect 25230 24670 25282 24722
rect 25282 24670 25284 24722
rect 25228 24668 25284 24670
rect 24332 24444 24388 24500
rect 24522 24330 24578 24332
rect 24522 24278 24524 24330
rect 24524 24278 24576 24330
rect 24576 24278 24578 24330
rect 24522 24276 24578 24278
rect 24626 24330 24682 24332
rect 24626 24278 24628 24330
rect 24628 24278 24680 24330
rect 24680 24278 24682 24330
rect 24626 24276 24682 24278
rect 24730 24330 24786 24332
rect 24730 24278 24732 24330
rect 24732 24278 24784 24330
rect 24784 24278 24786 24330
rect 24730 24276 24786 24278
rect 25228 24332 25284 24388
rect 24220 23938 24276 23940
rect 24220 23886 24222 23938
rect 24222 23886 24274 23938
rect 24274 23886 24276 23938
rect 24220 23884 24276 23886
rect 26796 25506 26852 25508
rect 26796 25454 26798 25506
rect 26798 25454 26850 25506
rect 26850 25454 26852 25506
rect 26796 25452 26852 25454
rect 27020 26012 27076 26068
rect 25788 24610 25844 24612
rect 25788 24558 25790 24610
rect 25790 24558 25842 24610
rect 25842 24558 25844 24610
rect 25788 24556 25844 24558
rect 25564 24498 25620 24500
rect 25564 24446 25566 24498
rect 25566 24446 25618 24498
rect 25618 24446 25620 24498
rect 25564 24444 25620 24446
rect 25676 24220 25732 24276
rect 25228 23324 25284 23380
rect 24444 23154 24500 23156
rect 24444 23102 24446 23154
rect 24446 23102 24498 23154
rect 24498 23102 24500 23154
rect 24444 23100 24500 23102
rect 24522 22762 24578 22764
rect 24522 22710 24524 22762
rect 24524 22710 24576 22762
rect 24576 22710 24578 22762
rect 24522 22708 24578 22710
rect 24626 22762 24682 22764
rect 24626 22710 24628 22762
rect 24628 22710 24680 22762
rect 24680 22710 24682 22762
rect 24626 22708 24682 22710
rect 24730 22762 24786 22764
rect 24730 22710 24732 22762
rect 24732 22710 24784 22762
rect 24784 22710 24786 22762
rect 24730 22708 24786 22710
rect 23324 21698 23380 21700
rect 23324 21646 23326 21698
rect 23326 21646 23378 21698
rect 23378 21646 23380 21698
rect 23324 21644 23380 21646
rect 22764 17666 22820 17668
rect 22764 17614 22766 17666
rect 22766 17614 22818 17666
rect 22818 17614 22820 17666
rect 22764 17612 22820 17614
rect 23212 20188 23268 20244
rect 23548 20524 23604 20580
rect 24668 22428 24724 22484
rect 26572 24556 26628 24612
rect 25900 22652 25956 22708
rect 25900 22258 25956 22260
rect 25900 22206 25902 22258
rect 25902 22206 25954 22258
rect 25954 22206 25956 22258
rect 25900 22204 25956 22206
rect 25676 21756 25732 21812
rect 24332 21532 24388 21588
rect 25228 21586 25284 21588
rect 25228 21534 25230 21586
rect 25230 21534 25282 21586
rect 25282 21534 25284 21586
rect 25228 21532 25284 21534
rect 26012 21644 26068 21700
rect 25564 21308 25620 21364
rect 24522 21194 24578 21196
rect 24522 21142 24524 21194
rect 24524 21142 24576 21194
rect 24576 21142 24578 21194
rect 24522 21140 24578 21142
rect 24626 21194 24682 21196
rect 24626 21142 24628 21194
rect 24628 21142 24680 21194
rect 24680 21142 24682 21194
rect 24626 21140 24682 21142
rect 24730 21194 24786 21196
rect 24730 21142 24732 21194
rect 24732 21142 24784 21194
rect 24784 21142 24786 21194
rect 24730 21140 24786 21142
rect 25228 21196 25284 21252
rect 23884 20188 23940 20244
rect 23772 20130 23828 20132
rect 23772 20078 23774 20130
rect 23774 20078 23826 20130
rect 23826 20078 23828 20130
rect 23772 20076 23828 20078
rect 23548 19740 23604 19796
rect 25564 20130 25620 20132
rect 25564 20078 25566 20130
rect 25566 20078 25618 20130
rect 25618 20078 25620 20130
rect 25564 20076 25620 20078
rect 24108 20018 24164 20020
rect 24108 19966 24110 20018
rect 24110 19966 24162 20018
rect 24162 19966 24164 20018
rect 24108 19964 24164 19966
rect 23996 19234 24052 19236
rect 23996 19182 23998 19234
rect 23998 19182 24050 19234
rect 24050 19182 24052 19234
rect 23996 19180 24052 19182
rect 23324 18284 23380 18340
rect 24522 19626 24578 19628
rect 24522 19574 24524 19626
rect 24524 19574 24576 19626
rect 24576 19574 24578 19626
rect 24522 19572 24578 19574
rect 24626 19626 24682 19628
rect 24626 19574 24628 19626
rect 24628 19574 24680 19626
rect 24680 19574 24682 19626
rect 24626 19572 24682 19574
rect 24730 19626 24786 19628
rect 24730 19574 24732 19626
rect 24732 19574 24784 19626
rect 24784 19574 24786 19626
rect 24730 19572 24786 19574
rect 25900 19292 25956 19348
rect 24108 18450 24164 18452
rect 24108 18398 24110 18450
rect 24110 18398 24162 18450
rect 24162 18398 24164 18450
rect 24108 18396 24164 18398
rect 24332 18284 24388 18340
rect 23548 17724 23604 17780
rect 24220 17778 24276 17780
rect 24220 17726 24222 17778
rect 24222 17726 24274 17778
rect 24274 17726 24276 17778
rect 24220 17724 24276 17726
rect 22988 17612 23044 17668
rect 23324 17388 23380 17444
rect 22876 16828 22932 16884
rect 22652 16716 22708 16772
rect 22316 15372 22372 15428
rect 22204 14476 22260 14532
rect 23212 16156 23268 16212
rect 23772 17554 23828 17556
rect 23772 17502 23774 17554
rect 23774 17502 23826 17554
rect 23826 17502 23828 17554
rect 23772 17500 23828 17502
rect 23660 17106 23716 17108
rect 23660 17054 23662 17106
rect 23662 17054 23714 17106
rect 23714 17054 23716 17106
rect 23660 17052 23716 17054
rect 23884 16828 23940 16884
rect 23772 16098 23828 16100
rect 23772 16046 23774 16098
rect 23774 16046 23826 16098
rect 23826 16046 23828 16098
rect 23772 16044 23828 16046
rect 23660 15484 23716 15540
rect 22988 15148 23044 15204
rect 25228 18396 25284 18452
rect 24522 18058 24578 18060
rect 24522 18006 24524 18058
rect 24524 18006 24576 18058
rect 24576 18006 24578 18058
rect 24522 18004 24578 18006
rect 24626 18058 24682 18060
rect 24626 18006 24628 18058
rect 24628 18006 24680 18058
rect 24680 18006 24682 18058
rect 24626 18004 24682 18006
rect 24730 18058 24786 18060
rect 24730 18006 24732 18058
rect 24732 18006 24784 18058
rect 24784 18006 24786 18058
rect 24730 18004 24786 18006
rect 25228 17948 25284 18004
rect 25788 17724 25844 17780
rect 24892 17666 24948 17668
rect 24892 17614 24894 17666
rect 24894 17614 24946 17666
rect 24946 17614 24948 17666
rect 24892 17612 24948 17614
rect 24668 17388 24724 17444
rect 24892 16828 24948 16884
rect 24522 16490 24578 16492
rect 24522 16438 24524 16490
rect 24524 16438 24576 16490
rect 24576 16438 24578 16490
rect 24522 16436 24578 16438
rect 24626 16490 24682 16492
rect 24626 16438 24628 16490
rect 24628 16438 24680 16490
rect 24680 16438 24682 16490
rect 24626 16436 24682 16438
rect 24730 16490 24786 16492
rect 24730 16438 24732 16490
rect 24732 16438 24784 16490
rect 24784 16438 24786 16490
rect 24730 16436 24786 16438
rect 25564 17666 25620 17668
rect 25564 17614 25566 17666
rect 25566 17614 25618 17666
rect 25618 17614 25620 17666
rect 25564 17612 25620 17614
rect 25004 16098 25060 16100
rect 25004 16046 25006 16098
rect 25006 16046 25058 16098
rect 25058 16046 25060 16098
rect 25004 16044 25060 16046
rect 25116 17388 25172 17444
rect 24556 15932 24612 15988
rect 25900 17388 25956 17444
rect 25788 17164 25844 17220
rect 25676 17106 25732 17108
rect 25676 17054 25678 17106
rect 25678 17054 25730 17106
rect 25730 17054 25732 17106
rect 25676 17052 25732 17054
rect 25564 15596 25620 15652
rect 26124 19292 26180 19348
rect 26572 23938 26628 23940
rect 26572 23886 26574 23938
rect 26574 23886 26626 23938
rect 26626 23886 26628 23938
rect 26572 23884 26628 23886
rect 26796 24892 26852 24948
rect 26796 24220 26852 24276
rect 26572 21980 26628 22036
rect 26460 21756 26516 21812
rect 26348 21644 26404 21700
rect 26684 21698 26740 21700
rect 26684 21646 26686 21698
rect 26686 21646 26738 21698
rect 26738 21646 26740 21698
rect 26684 21644 26740 21646
rect 26572 21586 26628 21588
rect 26572 21534 26574 21586
rect 26574 21534 26626 21586
rect 26626 21534 26628 21586
rect 26572 21532 26628 21534
rect 27804 27858 27860 27860
rect 27804 27806 27806 27858
rect 27806 27806 27858 27858
rect 27858 27806 27860 27858
rect 27804 27804 27860 27806
rect 29036 36258 29092 36260
rect 29036 36206 29038 36258
rect 29038 36206 29090 36258
rect 29090 36206 29092 36258
rect 29036 36204 29092 36206
rect 29820 36204 29876 36260
rect 29184 36090 29240 36092
rect 29184 36038 29186 36090
rect 29186 36038 29238 36090
rect 29238 36038 29240 36090
rect 29184 36036 29240 36038
rect 29288 36090 29344 36092
rect 29288 36038 29290 36090
rect 29290 36038 29342 36090
rect 29342 36038 29344 36090
rect 29288 36036 29344 36038
rect 29392 36090 29448 36092
rect 29392 36038 29394 36090
rect 29394 36038 29446 36090
rect 29446 36038 29448 36090
rect 29392 36036 29448 36038
rect 29184 34522 29240 34524
rect 29184 34470 29186 34522
rect 29186 34470 29238 34522
rect 29238 34470 29240 34522
rect 29184 34468 29240 34470
rect 29288 34522 29344 34524
rect 29288 34470 29290 34522
rect 29290 34470 29342 34522
rect 29342 34470 29344 34522
rect 29288 34468 29344 34470
rect 29392 34522 29448 34524
rect 29392 34470 29394 34522
rect 29394 34470 29446 34522
rect 29446 34470 29448 34522
rect 29392 34468 29448 34470
rect 30380 36258 30436 36260
rect 30380 36206 30382 36258
rect 30382 36206 30434 36258
rect 30434 36206 30436 36258
rect 30380 36204 30436 36206
rect 31612 36876 31668 36932
rect 32844 36876 32900 36932
rect 31164 36316 31220 36372
rect 30716 35308 30772 35364
rect 30044 33516 30100 33572
rect 29184 32954 29240 32956
rect 29184 32902 29186 32954
rect 29186 32902 29238 32954
rect 29238 32902 29240 32954
rect 29184 32900 29240 32902
rect 29288 32954 29344 32956
rect 29288 32902 29290 32954
rect 29290 32902 29342 32954
rect 29342 32902 29344 32954
rect 29288 32900 29344 32902
rect 29392 32954 29448 32956
rect 29392 32902 29394 32954
rect 29394 32902 29446 32954
rect 29446 32902 29448 32954
rect 29392 32900 29448 32902
rect 30380 31612 30436 31668
rect 29184 31386 29240 31388
rect 29184 31334 29186 31386
rect 29186 31334 29238 31386
rect 29238 31334 29240 31386
rect 29184 31332 29240 31334
rect 29288 31386 29344 31388
rect 29288 31334 29290 31386
rect 29290 31334 29342 31386
rect 29342 31334 29344 31386
rect 29288 31332 29344 31334
rect 29392 31386 29448 31388
rect 29392 31334 29394 31386
rect 29394 31334 29446 31386
rect 29446 31334 29448 31386
rect 29392 31332 29448 31334
rect 29932 30268 29988 30324
rect 29184 29818 29240 29820
rect 29184 29766 29186 29818
rect 29186 29766 29238 29818
rect 29238 29766 29240 29818
rect 29184 29764 29240 29766
rect 29288 29818 29344 29820
rect 29288 29766 29290 29818
rect 29290 29766 29342 29818
rect 29342 29766 29344 29818
rect 29288 29764 29344 29766
rect 29392 29818 29448 29820
rect 29392 29766 29394 29818
rect 29394 29766 29446 29818
rect 29446 29766 29448 29818
rect 29392 29764 29448 29766
rect 29184 28250 29240 28252
rect 29184 28198 29186 28250
rect 29186 28198 29238 28250
rect 29238 28198 29240 28250
rect 29184 28196 29240 28198
rect 29288 28250 29344 28252
rect 29288 28198 29290 28250
rect 29290 28198 29342 28250
rect 29342 28198 29344 28250
rect 29288 28196 29344 28198
rect 29392 28250 29448 28252
rect 29392 28198 29394 28250
rect 29394 28198 29446 28250
rect 29446 28198 29448 28250
rect 29392 28196 29448 28198
rect 29708 26796 29764 26852
rect 29184 26682 29240 26684
rect 29184 26630 29186 26682
rect 29186 26630 29238 26682
rect 29238 26630 29240 26682
rect 29184 26628 29240 26630
rect 29288 26682 29344 26684
rect 29288 26630 29290 26682
rect 29290 26630 29342 26682
rect 29342 26630 29344 26682
rect 29288 26628 29344 26630
rect 29392 26682 29448 26684
rect 29392 26630 29394 26682
rect 29394 26630 29446 26682
rect 29446 26630 29448 26682
rect 29392 26628 29448 26630
rect 27580 25564 27636 25620
rect 28028 25394 28084 25396
rect 28028 25342 28030 25394
rect 28030 25342 28082 25394
rect 28082 25342 28084 25394
rect 28028 25340 28084 25342
rect 27132 24892 27188 24948
rect 29184 25114 29240 25116
rect 29184 25062 29186 25114
rect 29186 25062 29238 25114
rect 29238 25062 29240 25114
rect 29184 25060 29240 25062
rect 29288 25114 29344 25116
rect 29288 25062 29290 25114
rect 29290 25062 29342 25114
rect 29342 25062 29344 25114
rect 29288 25060 29344 25062
rect 29392 25114 29448 25116
rect 29392 25062 29394 25114
rect 29394 25062 29446 25114
rect 29446 25062 29448 25114
rect 29392 25060 29448 25062
rect 30268 29372 30324 29428
rect 29932 27132 29988 27188
rect 28140 24610 28196 24612
rect 28140 24558 28142 24610
rect 28142 24558 28194 24610
rect 28194 24558 28196 24610
rect 28140 24556 28196 24558
rect 27804 24108 27860 24164
rect 27916 23548 27972 23604
rect 27580 23378 27636 23380
rect 27580 23326 27582 23378
rect 27582 23326 27634 23378
rect 27634 23326 27636 23378
rect 27580 23324 27636 23326
rect 28476 23826 28532 23828
rect 28476 23774 28478 23826
rect 28478 23774 28530 23826
rect 28530 23774 28532 23826
rect 28476 23772 28532 23774
rect 29148 23826 29204 23828
rect 29148 23774 29150 23826
rect 29150 23774 29202 23826
rect 29202 23774 29204 23826
rect 29148 23772 29204 23774
rect 29184 23546 29240 23548
rect 29184 23494 29186 23546
rect 29186 23494 29238 23546
rect 29238 23494 29240 23546
rect 29184 23492 29240 23494
rect 29288 23546 29344 23548
rect 29288 23494 29290 23546
rect 29290 23494 29342 23546
rect 29342 23494 29344 23546
rect 29288 23492 29344 23494
rect 29392 23546 29448 23548
rect 29392 23494 29394 23546
rect 29394 23494 29446 23546
rect 29446 23494 29448 23546
rect 29392 23492 29448 23494
rect 27804 22540 27860 22596
rect 27132 22258 27188 22260
rect 27132 22206 27134 22258
rect 27134 22206 27186 22258
rect 27186 22206 27188 22258
rect 27132 22204 27188 22206
rect 28700 23100 28756 23156
rect 27468 21756 27524 21812
rect 27804 21698 27860 21700
rect 27804 21646 27806 21698
rect 27806 21646 27858 21698
rect 27858 21646 27860 21698
rect 27804 21644 27860 21646
rect 27020 21420 27076 21476
rect 26348 20690 26404 20692
rect 26348 20638 26350 20690
rect 26350 20638 26402 20690
rect 26402 20638 26404 20690
rect 26348 20636 26404 20638
rect 27132 20636 27188 20692
rect 27468 20524 27524 20580
rect 28028 20690 28084 20692
rect 28028 20638 28030 20690
rect 28030 20638 28082 20690
rect 28082 20638 28084 20690
rect 28028 20636 28084 20638
rect 28588 22316 28644 22372
rect 26572 19292 26628 19348
rect 27020 20018 27076 20020
rect 27020 19966 27022 20018
rect 27022 19966 27074 20018
rect 27074 19966 27076 20018
rect 27020 19964 27076 19966
rect 27020 19740 27076 19796
rect 26124 17554 26180 17556
rect 26124 17502 26126 17554
rect 26126 17502 26178 17554
rect 26178 17502 26180 17554
rect 26124 17500 26180 17502
rect 27580 19234 27636 19236
rect 27580 19182 27582 19234
rect 27582 19182 27634 19234
rect 27634 19182 27636 19234
rect 27580 19180 27636 19182
rect 26348 17836 26404 17892
rect 25900 15426 25956 15428
rect 25900 15374 25902 15426
rect 25902 15374 25954 15426
rect 25954 15374 25956 15426
rect 25900 15372 25956 15374
rect 25676 15260 25732 15316
rect 24892 15148 24948 15204
rect 22316 14364 22372 14420
rect 22316 13970 22372 13972
rect 22316 13918 22318 13970
rect 22318 13918 22370 13970
rect 22370 13918 22372 13970
rect 22316 13916 22372 13918
rect 21420 13074 21476 13076
rect 21420 13022 21422 13074
rect 21422 13022 21474 13074
rect 21474 13022 21476 13074
rect 21420 13020 21476 13022
rect 21308 10108 21364 10164
rect 21420 11228 21476 11284
rect 19860 9434 19916 9436
rect 19860 9382 19862 9434
rect 19862 9382 19914 9434
rect 19914 9382 19916 9434
rect 19860 9380 19916 9382
rect 19964 9434 20020 9436
rect 19964 9382 19966 9434
rect 19966 9382 20018 9434
rect 20018 9382 20020 9434
rect 19964 9380 20020 9382
rect 20068 9434 20124 9436
rect 20068 9382 20070 9434
rect 20070 9382 20122 9434
rect 20122 9382 20124 9434
rect 20068 9380 20124 9382
rect 19740 9154 19796 9156
rect 19740 9102 19742 9154
rect 19742 9102 19794 9154
rect 19794 9102 19796 9154
rect 19740 9100 19796 9102
rect 19860 7866 19916 7868
rect 19860 7814 19862 7866
rect 19862 7814 19914 7866
rect 19914 7814 19916 7866
rect 19860 7812 19916 7814
rect 19964 7866 20020 7868
rect 19964 7814 19966 7866
rect 19966 7814 20018 7866
rect 20018 7814 20020 7866
rect 19964 7812 20020 7814
rect 20068 7866 20124 7868
rect 20068 7814 20070 7866
rect 20070 7814 20122 7866
rect 20122 7814 20124 7866
rect 20068 7812 20124 7814
rect 19860 6298 19916 6300
rect 19860 6246 19862 6298
rect 19862 6246 19914 6298
rect 19914 6246 19916 6298
rect 19860 6244 19916 6246
rect 19964 6298 20020 6300
rect 19964 6246 19966 6298
rect 19966 6246 20018 6298
rect 20018 6246 20020 6298
rect 19964 6244 20020 6246
rect 20068 6298 20124 6300
rect 20068 6246 20070 6298
rect 20070 6246 20122 6298
rect 20122 6246 20124 6298
rect 20068 6244 20124 6246
rect 20860 5852 20916 5908
rect 19860 4730 19916 4732
rect 19860 4678 19862 4730
rect 19862 4678 19914 4730
rect 19914 4678 19916 4730
rect 19860 4676 19916 4678
rect 19964 4730 20020 4732
rect 19964 4678 19966 4730
rect 19966 4678 20018 4730
rect 20018 4678 20020 4730
rect 19964 4676 20020 4678
rect 20068 4730 20124 4732
rect 20068 4678 20070 4730
rect 20070 4678 20122 4730
rect 20122 4678 20124 4730
rect 20068 4676 20124 4678
rect 19860 3162 19916 3164
rect 19860 3110 19862 3162
rect 19862 3110 19914 3162
rect 19914 3110 19916 3162
rect 19860 3108 19916 3110
rect 19964 3162 20020 3164
rect 19964 3110 19966 3162
rect 19966 3110 20018 3162
rect 20018 3110 20020 3162
rect 19964 3108 20020 3110
rect 20068 3162 20124 3164
rect 20068 3110 20070 3162
rect 20070 3110 20122 3162
rect 20122 3110 20124 3162
rect 20068 3108 20124 3110
rect 21756 11228 21812 11284
rect 21756 10722 21812 10724
rect 21756 10670 21758 10722
rect 21758 10670 21810 10722
rect 21810 10670 21812 10722
rect 21756 10668 21812 10670
rect 22092 12962 22148 12964
rect 22092 12910 22094 12962
rect 22094 12910 22146 12962
rect 22146 12910 22148 12962
rect 22092 12908 22148 12910
rect 22988 14476 23044 14532
rect 23212 14418 23268 14420
rect 23212 14366 23214 14418
rect 23214 14366 23266 14418
rect 23266 14366 23268 14418
rect 23212 14364 23268 14366
rect 23100 13468 23156 13524
rect 23100 12124 23156 12180
rect 23212 11676 23268 11732
rect 22092 11394 22148 11396
rect 22092 11342 22094 11394
rect 22094 11342 22146 11394
rect 22146 11342 22148 11394
rect 22092 11340 22148 11342
rect 21756 10220 21812 10276
rect 22540 10220 22596 10276
rect 21868 10108 21924 10164
rect 22316 9660 22372 9716
rect 22316 9100 22372 9156
rect 22428 8764 22484 8820
rect 22092 7980 22148 8036
rect 24522 14922 24578 14924
rect 24522 14870 24524 14922
rect 24524 14870 24576 14922
rect 24576 14870 24578 14922
rect 24522 14868 24578 14870
rect 24626 14922 24682 14924
rect 24626 14870 24628 14922
rect 24628 14870 24680 14922
rect 24680 14870 24682 14922
rect 24626 14868 24682 14870
rect 24730 14922 24786 14924
rect 24730 14870 24732 14922
rect 24732 14870 24784 14922
rect 24784 14870 24786 14922
rect 24730 14868 24786 14870
rect 23436 14530 23492 14532
rect 23436 14478 23438 14530
rect 23438 14478 23490 14530
rect 23490 14478 23492 14530
rect 23436 14476 23492 14478
rect 24780 14364 24836 14420
rect 23324 11564 23380 11620
rect 23212 10108 23268 10164
rect 23436 9660 23492 9716
rect 24522 13354 24578 13356
rect 24522 13302 24524 13354
rect 24524 13302 24576 13354
rect 24576 13302 24578 13354
rect 24522 13300 24578 13302
rect 24626 13354 24682 13356
rect 24626 13302 24628 13354
rect 24628 13302 24680 13354
rect 24680 13302 24682 13354
rect 24626 13300 24682 13302
rect 24730 13354 24786 13356
rect 24730 13302 24732 13354
rect 24732 13302 24784 13354
rect 24784 13302 24786 13354
rect 24730 13300 24786 13302
rect 25452 14418 25508 14420
rect 25452 14366 25454 14418
rect 25454 14366 25506 14418
rect 25506 14366 25508 14418
rect 25452 14364 25508 14366
rect 24556 12962 24612 12964
rect 24556 12910 24558 12962
rect 24558 12910 24610 12962
rect 24610 12910 24612 12962
rect 24556 12908 24612 12910
rect 24332 11900 24388 11956
rect 24220 11676 24276 11732
rect 24522 11786 24578 11788
rect 24522 11734 24524 11786
rect 24524 11734 24576 11786
rect 24576 11734 24578 11786
rect 24522 11732 24578 11734
rect 24626 11786 24682 11788
rect 24626 11734 24628 11786
rect 24628 11734 24680 11786
rect 24680 11734 24682 11786
rect 24626 11732 24682 11734
rect 24730 11786 24786 11788
rect 24730 11734 24732 11786
rect 24732 11734 24784 11786
rect 24784 11734 24786 11786
rect 24730 11732 24786 11734
rect 23996 10332 24052 10388
rect 24220 11506 24276 11508
rect 24220 11454 24222 11506
rect 24222 11454 24274 11506
rect 24274 11454 24276 11506
rect 24220 11452 24276 11454
rect 25228 13468 25284 13524
rect 25004 12124 25060 12180
rect 25564 13858 25620 13860
rect 25564 13806 25566 13858
rect 25566 13806 25618 13858
rect 25618 13806 25620 13858
rect 25564 13804 25620 13806
rect 26236 15596 26292 15652
rect 28140 19122 28196 19124
rect 28140 19070 28142 19122
rect 28142 19070 28194 19122
rect 28194 19070 28196 19122
rect 28140 19068 28196 19070
rect 27468 18284 27524 18340
rect 27132 17388 27188 17444
rect 26572 16994 26628 16996
rect 26572 16942 26574 16994
rect 26574 16942 26626 16994
rect 26626 16942 26628 16994
rect 26572 16940 26628 16942
rect 28588 20130 28644 20132
rect 28588 20078 28590 20130
rect 28590 20078 28642 20130
rect 28642 20078 28644 20130
rect 28588 20076 28644 20078
rect 28588 17612 28644 17668
rect 28364 17164 28420 17220
rect 27244 16994 27300 16996
rect 27244 16942 27246 16994
rect 27246 16942 27298 16994
rect 27298 16942 27300 16994
rect 27244 16940 27300 16942
rect 27132 16882 27188 16884
rect 27132 16830 27134 16882
rect 27134 16830 27186 16882
rect 27186 16830 27188 16882
rect 27132 16828 27188 16830
rect 29036 23154 29092 23156
rect 29036 23102 29038 23154
rect 29038 23102 29090 23154
rect 29090 23102 29092 23154
rect 29036 23100 29092 23102
rect 29372 22764 29428 22820
rect 29596 22652 29652 22708
rect 29820 22370 29876 22372
rect 29820 22318 29822 22370
rect 29822 22318 29874 22370
rect 29874 22318 29876 22370
rect 29820 22316 29876 22318
rect 32172 36370 32228 36372
rect 32172 36318 32174 36370
rect 32174 36318 32226 36370
rect 32226 36318 32228 36370
rect 32172 36316 32228 36318
rect 31388 28476 31444 28532
rect 31500 34748 31556 34804
rect 30380 26796 30436 26852
rect 30492 27692 30548 27748
rect 30268 23324 30324 23380
rect 31276 24668 31332 24724
rect 30380 23212 30436 23268
rect 30604 23266 30660 23268
rect 30604 23214 30606 23266
rect 30606 23214 30658 23266
rect 30658 23214 30660 23266
rect 30604 23212 30660 23214
rect 30716 22764 30772 22820
rect 30492 22652 30548 22708
rect 31388 22764 31444 22820
rect 29932 22204 29988 22260
rect 29184 21978 29240 21980
rect 29184 21926 29186 21978
rect 29186 21926 29238 21978
rect 29238 21926 29240 21978
rect 29184 21924 29240 21926
rect 29288 21978 29344 21980
rect 29288 21926 29290 21978
rect 29290 21926 29342 21978
rect 29342 21926 29344 21978
rect 29288 21924 29344 21926
rect 29392 21978 29448 21980
rect 29392 21926 29394 21978
rect 29394 21926 29446 21978
rect 29446 21926 29448 21978
rect 29392 21924 29448 21926
rect 28924 21810 28980 21812
rect 28924 21758 28926 21810
rect 28926 21758 28978 21810
rect 28978 21758 28980 21810
rect 28924 21756 28980 21758
rect 30156 21698 30212 21700
rect 30156 21646 30158 21698
rect 30158 21646 30210 21698
rect 30210 21646 30212 21698
rect 30156 21644 30212 21646
rect 29932 20972 29988 21028
rect 31388 22092 31444 22148
rect 32956 36316 33012 36372
rect 32284 33628 32340 33684
rect 33846 36874 33902 36876
rect 33846 36822 33848 36874
rect 33848 36822 33900 36874
rect 33900 36822 33902 36874
rect 33846 36820 33902 36822
rect 33950 36874 34006 36876
rect 33950 36822 33952 36874
rect 33952 36822 34004 36874
rect 34004 36822 34006 36874
rect 33950 36820 34006 36822
rect 34054 36874 34110 36876
rect 34054 36822 34056 36874
rect 34056 36822 34108 36874
rect 34108 36822 34110 36874
rect 34054 36820 34110 36822
rect 33740 35922 33796 35924
rect 33740 35870 33742 35922
rect 33742 35870 33794 35922
rect 33794 35870 33796 35922
rect 33740 35868 33796 35870
rect 33180 35586 33236 35588
rect 33180 35534 33182 35586
rect 33182 35534 33234 35586
rect 33234 35534 33236 35586
rect 33180 35532 33236 35534
rect 32172 33068 32228 33124
rect 31500 21196 31556 21252
rect 31612 22370 31668 22372
rect 31612 22318 31614 22370
rect 31614 22318 31666 22370
rect 31666 22318 31668 22370
rect 31612 22316 31668 22318
rect 29260 20802 29316 20804
rect 29260 20750 29262 20802
rect 29262 20750 29314 20802
rect 29314 20750 29316 20802
rect 29260 20748 29316 20750
rect 29184 20410 29240 20412
rect 29184 20358 29186 20410
rect 29186 20358 29238 20410
rect 29238 20358 29240 20410
rect 29184 20356 29240 20358
rect 29288 20410 29344 20412
rect 29288 20358 29290 20410
rect 29290 20358 29342 20410
rect 29342 20358 29344 20410
rect 29288 20356 29344 20358
rect 29392 20410 29448 20412
rect 29392 20358 29394 20410
rect 29394 20358 29446 20410
rect 29446 20358 29448 20410
rect 29392 20356 29448 20358
rect 30492 20914 30548 20916
rect 30492 20862 30494 20914
rect 30494 20862 30546 20914
rect 30546 20862 30548 20914
rect 30492 20860 30548 20862
rect 34188 36370 34244 36372
rect 34188 36318 34190 36370
rect 34190 36318 34242 36370
rect 34242 36318 34244 36370
rect 34188 36316 34244 36318
rect 36316 36876 36372 36932
rect 37324 36876 37380 36932
rect 34972 36316 35028 36372
rect 34412 36092 34468 36148
rect 33852 35532 33908 35588
rect 35980 36370 36036 36372
rect 35980 36318 35982 36370
rect 35982 36318 36034 36370
rect 36034 36318 36036 36370
rect 35980 36316 36036 36318
rect 33846 35306 33902 35308
rect 33846 35254 33848 35306
rect 33848 35254 33900 35306
rect 33900 35254 33902 35306
rect 33846 35252 33902 35254
rect 33950 35306 34006 35308
rect 33950 35254 33952 35306
rect 33952 35254 34004 35306
rect 34004 35254 34006 35306
rect 33950 35252 34006 35254
rect 34054 35306 34110 35308
rect 34054 35254 34056 35306
rect 34056 35254 34108 35306
rect 34108 35254 34110 35306
rect 34054 35252 34110 35254
rect 33846 33738 33902 33740
rect 33846 33686 33848 33738
rect 33848 33686 33900 33738
rect 33900 33686 33902 33738
rect 33846 33684 33902 33686
rect 33950 33738 34006 33740
rect 33950 33686 33952 33738
rect 33952 33686 34004 33738
rect 34004 33686 34006 33738
rect 33950 33684 34006 33686
rect 34054 33738 34110 33740
rect 34054 33686 34056 33738
rect 34056 33686 34108 33738
rect 34108 33686 34110 33738
rect 34054 33684 34110 33686
rect 33846 32170 33902 32172
rect 33846 32118 33848 32170
rect 33848 32118 33900 32170
rect 33900 32118 33902 32170
rect 33846 32116 33902 32118
rect 33950 32170 34006 32172
rect 33950 32118 33952 32170
rect 33952 32118 34004 32170
rect 34004 32118 34006 32170
rect 33950 32116 34006 32118
rect 34054 32170 34110 32172
rect 34054 32118 34056 32170
rect 34056 32118 34108 32170
rect 34108 32118 34110 32170
rect 34054 32116 34110 32118
rect 32956 31164 33012 31220
rect 32396 30044 32452 30100
rect 32508 22764 32564 22820
rect 32284 22370 32340 22372
rect 32284 22318 32286 22370
rect 32286 22318 32338 22370
rect 32338 22318 32340 22370
rect 32284 22316 32340 22318
rect 32396 21868 32452 21924
rect 33846 30602 33902 30604
rect 33846 30550 33848 30602
rect 33848 30550 33900 30602
rect 33900 30550 33902 30602
rect 33846 30548 33902 30550
rect 33950 30602 34006 30604
rect 33950 30550 33952 30602
rect 33952 30550 34004 30602
rect 34004 30550 34006 30602
rect 33950 30548 34006 30550
rect 34054 30602 34110 30604
rect 34054 30550 34056 30602
rect 34056 30550 34108 30602
rect 34108 30550 34110 30602
rect 34054 30548 34110 30550
rect 33846 29034 33902 29036
rect 33846 28982 33848 29034
rect 33848 28982 33900 29034
rect 33900 28982 33902 29034
rect 33846 28980 33902 28982
rect 33950 29034 34006 29036
rect 33950 28982 33952 29034
rect 33952 28982 34004 29034
rect 34004 28982 34006 29034
rect 33950 28980 34006 28982
rect 34054 29034 34110 29036
rect 34054 28982 34056 29034
rect 34056 28982 34108 29034
rect 34108 28982 34110 29034
rect 34054 28980 34110 28982
rect 33846 27466 33902 27468
rect 33846 27414 33848 27466
rect 33848 27414 33900 27466
rect 33900 27414 33902 27466
rect 33846 27412 33902 27414
rect 33950 27466 34006 27468
rect 33950 27414 33952 27466
rect 33952 27414 34004 27466
rect 34004 27414 34006 27466
rect 33950 27412 34006 27414
rect 34054 27466 34110 27468
rect 34054 27414 34056 27466
rect 34056 27414 34108 27466
rect 34108 27414 34110 27466
rect 34054 27412 34110 27414
rect 33068 26460 33124 26516
rect 35308 35420 35364 35476
rect 34412 35308 34468 35364
rect 34412 30268 34468 30324
rect 35756 27244 35812 27300
rect 36092 33964 36148 34020
rect 34188 26012 34244 26068
rect 35308 26908 35364 26964
rect 33846 25898 33902 25900
rect 33846 25846 33848 25898
rect 33848 25846 33900 25898
rect 33900 25846 33902 25898
rect 33846 25844 33902 25846
rect 33950 25898 34006 25900
rect 33950 25846 33952 25898
rect 33952 25846 34004 25898
rect 34004 25846 34006 25898
rect 33950 25844 34006 25846
rect 34054 25898 34110 25900
rect 34054 25846 34056 25898
rect 34056 25846 34108 25898
rect 34108 25846 34110 25898
rect 34054 25844 34110 25846
rect 35308 24780 35364 24836
rect 33846 24330 33902 24332
rect 33846 24278 33848 24330
rect 33848 24278 33900 24330
rect 33900 24278 33902 24330
rect 33846 24276 33902 24278
rect 33950 24330 34006 24332
rect 33950 24278 33952 24330
rect 33952 24278 34004 24330
rect 34004 24278 34006 24330
rect 33950 24276 34006 24278
rect 34054 24330 34110 24332
rect 34054 24278 34056 24330
rect 34056 24278 34108 24330
rect 34108 24278 34110 24330
rect 34054 24276 34110 24278
rect 35308 23772 35364 23828
rect 33846 22762 33902 22764
rect 33846 22710 33848 22762
rect 33848 22710 33900 22762
rect 33900 22710 33902 22762
rect 33846 22708 33902 22710
rect 33950 22762 34006 22764
rect 33950 22710 33952 22762
rect 33952 22710 34004 22762
rect 34004 22710 34006 22762
rect 33950 22708 34006 22710
rect 34054 22762 34110 22764
rect 34054 22710 34056 22762
rect 34056 22710 34108 22762
rect 34108 22710 34110 22762
rect 34054 22708 34110 22710
rect 35308 22428 35364 22484
rect 32060 21308 32116 21364
rect 31612 20860 31668 20916
rect 30716 20802 30772 20804
rect 30716 20750 30718 20802
rect 30718 20750 30770 20802
rect 30770 20750 30772 20802
rect 30716 20748 30772 20750
rect 31724 20690 31780 20692
rect 31724 20638 31726 20690
rect 31726 20638 31778 20690
rect 31778 20638 31780 20690
rect 31724 20636 31780 20638
rect 31164 20524 31220 20580
rect 31836 20524 31892 20580
rect 33846 21194 33902 21196
rect 33846 21142 33848 21194
rect 33848 21142 33900 21194
rect 33900 21142 33902 21194
rect 33846 21140 33902 21142
rect 33950 21194 34006 21196
rect 33950 21142 33952 21194
rect 33952 21142 34004 21194
rect 34004 21142 34006 21194
rect 33950 21140 34006 21142
rect 34054 21194 34110 21196
rect 34054 21142 34056 21194
rect 34056 21142 34108 21194
rect 34108 21142 34110 21194
rect 34054 21140 34110 21142
rect 32284 20914 32340 20916
rect 32284 20862 32286 20914
rect 32286 20862 32338 20914
rect 32338 20862 32340 20914
rect 32284 20860 32340 20862
rect 32956 20690 33012 20692
rect 32956 20638 32958 20690
rect 32958 20638 33010 20690
rect 33010 20638 33012 20690
rect 32956 20636 33012 20638
rect 33292 20690 33348 20692
rect 33292 20638 33294 20690
rect 33294 20638 33346 20690
rect 33346 20638 33348 20690
rect 33292 20636 33348 20638
rect 36316 24556 36372 24612
rect 37548 35644 37604 35700
rect 38508 36090 38564 36092
rect 38508 36038 38510 36090
rect 38510 36038 38562 36090
rect 38562 36038 38564 36090
rect 38508 36036 38564 36038
rect 38612 36090 38668 36092
rect 38612 36038 38614 36090
rect 38614 36038 38666 36090
rect 38666 36038 38668 36090
rect 38612 36036 38668 36038
rect 38716 36090 38772 36092
rect 38716 36038 38718 36090
rect 38718 36038 38770 36090
rect 38770 36038 38772 36090
rect 38716 36036 38772 36038
rect 37884 35308 37940 35364
rect 38220 34972 38276 35028
rect 37660 34802 37716 34804
rect 37660 34750 37662 34802
rect 37662 34750 37714 34802
rect 37714 34750 37716 34802
rect 37660 34748 37716 34750
rect 38508 34522 38564 34524
rect 38508 34470 38510 34522
rect 38510 34470 38562 34522
rect 38562 34470 38564 34522
rect 38508 34468 38564 34470
rect 38612 34522 38668 34524
rect 38612 34470 38614 34522
rect 38614 34470 38666 34522
rect 38666 34470 38668 34522
rect 38612 34468 38668 34470
rect 38716 34522 38772 34524
rect 38716 34470 38718 34522
rect 38718 34470 38770 34522
rect 38770 34470 38772 34522
rect 38716 34468 38772 34470
rect 38444 34300 38500 34356
rect 37548 34018 37604 34020
rect 37548 33966 37550 34018
rect 37550 33966 37602 34018
rect 37602 33966 37604 34018
rect 37548 33964 37604 33966
rect 37996 33964 38052 34020
rect 38220 33628 38276 33684
rect 37660 33122 37716 33124
rect 37660 33070 37662 33122
rect 37662 33070 37714 33122
rect 37714 33070 37716 33122
rect 37660 33068 37716 33070
rect 38220 33122 38276 33124
rect 38220 33070 38222 33122
rect 38222 33070 38274 33122
rect 38274 33070 38276 33122
rect 38220 33068 38276 33070
rect 38508 32954 38564 32956
rect 38508 32902 38510 32954
rect 38510 32902 38562 32954
rect 38562 32902 38564 32954
rect 38508 32900 38564 32902
rect 38612 32954 38668 32956
rect 38612 32902 38614 32954
rect 38614 32902 38666 32954
rect 38666 32902 38668 32954
rect 38612 32900 38668 32902
rect 38716 32954 38772 32956
rect 38716 32902 38718 32954
rect 38718 32902 38770 32954
rect 38770 32902 38772 32954
rect 38716 32900 38772 32902
rect 37548 32562 37604 32564
rect 37548 32510 37550 32562
rect 37550 32510 37602 32562
rect 37602 32510 37604 32562
rect 37548 32508 37604 32510
rect 37996 32562 38052 32564
rect 37996 32510 37998 32562
rect 37998 32510 38050 32562
rect 38050 32510 38052 32562
rect 37996 32508 38052 32510
rect 38220 32284 38276 32340
rect 37212 31666 37268 31668
rect 37212 31614 37214 31666
rect 37214 31614 37266 31666
rect 37266 31614 37268 31666
rect 37212 31612 37268 31614
rect 37548 31666 37604 31668
rect 37548 31614 37550 31666
rect 37550 31614 37602 31666
rect 37602 31614 37604 31666
rect 37548 31612 37604 31614
rect 37884 31164 37940 31220
rect 37884 30994 37940 30996
rect 37884 30942 37886 30994
rect 37886 30942 37938 30994
rect 37938 30942 37940 30994
rect 37884 30940 37940 30942
rect 37100 30380 37156 30436
rect 38508 31386 38564 31388
rect 38508 31334 38510 31386
rect 38510 31334 38562 31386
rect 38562 31334 38564 31386
rect 38508 31332 38564 31334
rect 38612 31386 38668 31388
rect 38612 31334 38614 31386
rect 38614 31334 38666 31386
rect 38666 31334 38668 31386
rect 38612 31332 38668 31334
rect 38716 31386 38772 31388
rect 38716 31334 38718 31386
rect 38718 31334 38770 31386
rect 38770 31334 38772 31386
rect 38716 31332 38772 31334
rect 38444 30940 38500 30996
rect 38220 30268 38276 30324
rect 37884 30098 37940 30100
rect 37884 30046 37886 30098
rect 37886 30046 37938 30098
rect 37938 30046 37940 30098
rect 37884 30044 37940 30046
rect 38220 29708 38276 29764
rect 38508 29818 38564 29820
rect 38508 29766 38510 29818
rect 38510 29766 38562 29818
rect 38562 29766 38564 29818
rect 38508 29764 38564 29766
rect 38612 29818 38668 29820
rect 38612 29766 38614 29818
rect 38614 29766 38666 29818
rect 38666 29766 38668 29818
rect 38612 29764 38668 29766
rect 38716 29818 38772 29820
rect 38716 29766 38718 29818
rect 38718 29766 38770 29818
rect 38770 29766 38772 29818
rect 38716 29764 38772 29766
rect 37884 29426 37940 29428
rect 37884 29374 37886 29426
rect 37886 29374 37938 29426
rect 37938 29374 37940 29426
rect 37884 29372 37940 29374
rect 38220 28924 38276 28980
rect 37548 27746 37604 27748
rect 37548 27694 37550 27746
rect 37550 27694 37602 27746
rect 37602 27694 37604 27746
rect 37548 27692 37604 27694
rect 37212 27132 37268 27188
rect 37548 27020 37604 27076
rect 38220 28418 38276 28420
rect 38220 28366 38222 28418
rect 38222 28366 38274 28418
rect 38274 28366 38276 28418
rect 38220 28364 38276 28366
rect 38508 28250 38564 28252
rect 38508 28198 38510 28250
rect 38510 28198 38562 28250
rect 38562 28198 38564 28250
rect 38508 28196 38564 28198
rect 38612 28250 38668 28252
rect 38612 28198 38614 28250
rect 38614 28198 38666 28250
rect 38666 28198 38668 28250
rect 38612 28196 38668 28198
rect 38716 28250 38772 28252
rect 38716 28198 38718 28250
rect 38718 28198 38770 28250
rect 38770 28198 38772 28250
rect 38716 28196 38772 28198
rect 37996 27692 38052 27748
rect 38220 27580 38276 27636
rect 37884 26962 37940 26964
rect 37884 26910 37886 26962
rect 37886 26910 37938 26962
rect 37938 26910 37940 26962
rect 37884 26908 37940 26910
rect 37660 25340 37716 25396
rect 38508 26682 38564 26684
rect 38508 26630 38510 26682
rect 38510 26630 38562 26682
rect 38562 26630 38564 26682
rect 38508 26628 38564 26630
rect 38612 26682 38668 26684
rect 38612 26630 38614 26682
rect 38614 26630 38666 26682
rect 38666 26630 38668 26682
rect 38612 26628 38668 26630
rect 38716 26682 38772 26684
rect 38716 26630 38718 26682
rect 38718 26630 38770 26682
rect 38770 26630 38772 26682
rect 38716 26628 38772 26630
rect 38108 26236 38164 26292
rect 38220 25564 38276 25620
rect 37884 24722 37940 24724
rect 37884 24670 37886 24722
rect 37886 24670 37938 24722
rect 37938 24670 37940 24722
rect 37884 24668 37940 24670
rect 37772 24108 37828 24164
rect 37884 23826 37940 23828
rect 37884 23774 37886 23826
rect 37886 23774 37938 23826
rect 37938 23774 37940 23826
rect 37884 23772 37940 23774
rect 36876 23212 36932 23268
rect 37884 22540 37940 22596
rect 38220 25282 38276 25284
rect 38220 25230 38222 25282
rect 38222 25230 38274 25282
rect 38274 25230 38276 25282
rect 38220 25228 38276 25230
rect 38508 25114 38564 25116
rect 38508 25062 38510 25114
rect 38510 25062 38562 25114
rect 38562 25062 38564 25114
rect 38508 25060 38564 25062
rect 38612 25114 38668 25116
rect 38612 25062 38614 25114
rect 38614 25062 38666 25114
rect 38666 25062 38668 25114
rect 38612 25060 38668 25062
rect 38716 25114 38772 25116
rect 38716 25062 38718 25114
rect 38718 25062 38770 25114
rect 38770 25062 38772 25114
rect 38716 25060 38772 25062
rect 38220 24220 38276 24276
rect 38220 23714 38276 23716
rect 38220 23662 38222 23714
rect 38222 23662 38274 23714
rect 38274 23662 38276 23714
rect 38220 23660 38276 23662
rect 38508 23546 38564 23548
rect 38508 23494 38510 23546
rect 38510 23494 38562 23546
rect 38562 23494 38564 23546
rect 38508 23492 38564 23494
rect 38612 23546 38668 23548
rect 38612 23494 38614 23546
rect 38614 23494 38666 23546
rect 38666 23494 38668 23546
rect 38612 23492 38668 23494
rect 38716 23546 38772 23548
rect 38716 23494 38718 23546
rect 38718 23494 38770 23546
rect 38770 23494 38772 23546
rect 38716 23492 38772 23494
rect 38220 22876 38276 22932
rect 38220 22258 38276 22260
rect 38220 22206 38222 22258
rect 38222 22206 38274 22258
rect 38274 22206 38276 22258
rect 38220 22204 38276 22206
rect 37996 21868 38052 21924
rect 38508 21978 38564 21980
rect 38508 21926 38510 21978
rect 38510 21926 38562 21978
rect 38562 21926 38564 21978
rect 38508 21924 38564 21926
rect 38612 21978 38668 21980
rect 38612 21926 38614 21978
rect 38614 21926 38666 21978
rect 38666 21926 38668 21978
rect 38612 21924 38668 21926
rect 38716 21978 38772 21980
rect 38716 21926 38718 21978
rect 38718 21926 38770 21978
rect 38770 21926 38772 21978
rect 38716 21924 38772 21926
rect 37772 21756 37828 21812
rect 37884 21698 37940 21700
rect 37884 21646 37886 21698
rect 37886 21646 37938 21698
rect 37938 21646 37940 21698
rect 37884 21644 37940 21646
rect 37548 21532 37604 21588
rect 37212 20972 37268 21028
rect 38220 20860 38276 20916
rect 37884 20802 37940 20804
rect 37884 20750 37886 20802
rect 37886 20750 37938 20802
rect 37938 20750 37940 20802
rect 37884 20748 37940 20750
rect 36092 20636 36148 20692
rect 29036 19964 29092 20020
rect 38508 20410 38564 20412
rect 38508 20358 38510 20410
rect 38510 20358 38562 20410
rect 38562 20358 38564 20410
rect 38508 20356 38564 20358
rect 38612 20410 38668 20412
rect 38612 20358 38614 20410
rect 38614 20358 38666 20410
rect 38666 20358 38668 20410
rect 38612 20356 38668 20358
rect 38716 20410 38772 20412
rect 38716 20358 38718 20410
rect 38718 20358 38770 20410
rect 38770 20358 38772 20410
rect 38716 20356 38772 20358
rect 38444 20188 38500 20244
rect 36540 20076 36596 20132
rect 33846 19626 33902 19628
rect 33846 19574 33848 19626
rect 33848 19574 33900 19626
rect 33900 19574 33902 19626
rect 33846 19572 33902 19574
rect 33950 19626 34006 19628
rect 33950 19574 33952 19626
rect 33952 19574 34004 19626
rect 34004 19574 34006 19626
rect 33950 19572 34006 19574
rect 34054 19626 34110 19628
rect 34054 19574 34056 19626
rect 34056 19574 34108 19626
rect 34108 19574 34110 19626
rect 34054 19572 34110 19574
rect 32956 19404 33012 19460
rect 29596 19180 29652 19236
rect 29148 19122 29204 19124
rect 29148 19070 29150 19122
rect 29150 19070 29202 19122
rect 29202 19070 29204 19122
rect 29148 19068 29204 19070
rect 29484 19010 29540 19012
rect 29484 18958 29486 19010
rect 29486 18958 29538 19010
rect 29538 18958 29540 19010
rect 29484 18956 29540 18958
rect 29184 18842 29240 18844
rect 29184 18790 29186 18842
rect 29186 18790 29238 18842
rect 29238 18790 29240 18842
rect 29184 18788 29240 18790
rect 29288 18842 29344 18844
rect 29288 18790 29290 18842
rect 29290 18790 29342 18842
rect 29342 18790 29344 18842
rect 29288 18788 29344 18790
rect 29392 18842 29448 18844
rect 29392 18790 29394 18842
rect 29394 18790 29446 18842
rect 29446 18790 29448 18842
rect 29392 18788 29448 18790
rect 29596 18450 29652 18452
rect 29596 18398 29598 18450
rect 29598 18398 29650 18450
rect 29650 18398 29652 18450
rect 29596 18396 29652 18398
rect 30156 19068 30212 19124
rect 30940 19122 30996 19124
rect 30940 19070 30942 19122
rect 30942 19070 30994 19122
rect 30994 19070 30996 19122
rect 30940 19068 30996 19070
rect 29820 18226 29876 18228
rect 29820 18174 29822 18226
rect 29822 18174 29874 18226
rect 29874 18174 29876 18226
rect 29820 18172 29876 18174
rect 28924 17164 28980 17220
rect 29184 17274 29240 17276
rect 29184 17222 29186 17274
rect 29186 17222 29238 17274
rect 29238 17222 29240 17274
rect 29184 17220 29240 17222
rect 29288 17274 29344 17276
rect 29288 17222 29290 17274
rect 29290 17222 29342 17274
rect 29342 17222 29344 17274
rect 29288 17220 29344 17222
rect 29392 17274 29448 17276
rect 29392 17222 29394 17274
rect 29394 17222 29446 17274
rect 29446 17222 29448 17274
rect 29392 17220 29448 17222
rect 28364 15820 28420 15876
rect 26572 15372 26628 15428
rect 26012 13356 26068 13412
rect 28812 15538 28868 15540
rect 28812 15486 28814 15538
rect 28814 15486 28866 15538
rect 28866 15486 28868 15538
rect 28812 15484 28868 15486
rect 26572 14476 26628 14532
rect 27580 15148 27636 15204
rect 27356 14476 27412 14532
rect 28028 14476 28084 14532
rect 27244 13916 27300 13972
rect 26572 13746 26628 13748
rect 26572 13694 26574 13746
rect 26574 13694 26626 13746
rect 26626 13694 26628 13746
rect 26572 13692 26628 13694
rect 27580 13746 27636 13748
rect 27580 13694 27582 13746
rect 27582 13694 27634 13746
rect 27634 13694 27636 13746
rect 27580 13692 27636 13694
rect 26684 13468 26740 13524
rect 26572 13244 26628 13300
rect 25788 12850 25844 12852
rect 25788 12798 25790 12850
rect 25790 12798 25842 12850
rect 25842 12798 25844 12850
rect 25788 12796 25844 12798
rect 25228 11676 25284 11732
rect 25788 12402 25844 12404
rect 25788 12350 25790 12402
rect 25790 12350 25842 12402
rect 25842 12350 25844 12402
rect 25788 12348 25844 12350
rect 25452 12178 25508 12180
rect 25452 12126 25454 12178
rect 25454 12126 25506 12178
rect 25506 12126 25508 12178
rect 25452 12124 25508 12126
rect 25900 11900 25956 11956
rect 24892 11340 24948 11396
rect 24556 11282 24612 11284
rect 24556 11230 24558 11282
rect 24558 11230 24610 11282
rect 24610 11230 24612 11282
rect 24556 11228 24612 11230
rect 24668 10610 24724 10612
rect 24668 10558 24670 10610
rect 24670 10558 24722 10610
rect 24722 10558 24724 10610
rect 24668 10556 24724 10558
rect 23548 9212 23604 9268
rect 23324 9154 23380 9156
rect 23324 9102 23326 9154
rect 23326 9102 23378 9154
rect 23378 9102 23380 9154
rect 23324 9100 23380 9102
rect 23548 9042 23604 9044
rect 23548 8990 23550 9042
rect 23550 8990 23602 9042
rect 23602 8990 23604 9042
rect 23548 8988 23604 8990
rect 23884 8988 23940 9044
rect 22876 8764 22932 8820
rect 22876 8428 22932 8484
rect 23100 8146 23156 8148
rect 23100 8094 23102 8146
rect 23102 8094 23154 8146
rect 23154 8094 23156 8146
rect 23100 8092 23156 8094
rect 22876 8034 22932 8036
rect 22876 7982 22878 8034
rect 22878 7982 22930 8034
rect 22930 7982 22932 8034
rect 22876 7980 22932 7982
rect 22988 7474 23044 7476
rect 22988 7422 22990 7474
rect 22990 7422 23042 7474
rect 23042 7422 23044 7474
rect 22988 7420 23044 7422
rect 23660 8204 23716 8260
rect 24108 8764 24164 8820
rect 24522 10218 24578 10220
rect 24522 10166 24524 10218
rect 24524 10166 24576 10218
rect 24576 10166 24578 10218
rect 24522 10164 24578 10166
rect 24626 10218 24682 10220
rect 24626 10166 24628 10218
rect 24628 10166 24680 10218
rect 24680 10166 24682 10218
rect 24626 10164 24682 10166
rect 24730 10218 24786 10220
rect 24730 10166 24732 10218
rect 24732 10166 24784 10218
rect 24784 10166 24786 10218
rect 24730 10164 24786 10166
rect 24892 9714 24948 9716
rect 24892 9662 24894 9714
rect 24894 9662 24946 9714
rect 24946 9662 24948 9714
rect 24892 9660 24948 9662
rect 25564 11394 25620 11396
rect 25564 11342 25566 11394
rect 25566 11342 25618 11394
rect 25618 11342 25620 11394
rect 25564 11340 25620 11342
rect 24332 8988 24388 9044
rect 23996 7868 24052 7924
rect 24220 8258 24276 8260
rect 24220 8206 24222 8258
rect 24222 8206 24274 8258
rect 24274 8206 24276 8258
rect 24220 8204 24276 8206
rect 24522 8650 24578 8652
rect 24522 8598 24524 8650
rect 24524 8598 24576 8650
rect 24576 8598 24578 8650
rect 24522 8596 24578 8598
rect 24626 8650 24682 8652
rect 24626 8598 24628 8650
rect 24628 8598 24680 8650
rect 24680 8598 24682 8650
rect 24626 8596 24682 8598
rect 24730 8650 24786 8652
rect 24730 8598 24732 8650
rect 24732 8598 24784 8650
rect 24784 8598 24786 8650
rect 24730 8596 24786 8598
rect 24668 8316 24724 8372
rect 24780 8258 24836 8260
rect 24780 8206 24782 8258
rect 24782 8206 24834 8258
rect 24834 8206 24836 8258
rect 24780 8204 24836 8206
rect 24668 8092 24724 8148
rect 24556 8034 24612 8036
rect 24556 7982 24558 8034
rect 24558 7982 24610 8034
rect 24610 7982 24612 8034
rect 24556 7980 24612 7982
rect 24522 7082 24578 7084
rect 24522 7030 24524 7082
rect 24524 7030 24576 7082
rect 24576 7030 24578 7082
rect 24522 7028 24578 7030
rect 24626 7082 24682 7084
rect 24626 7030 24628 7082
rect 24628 7030 24680 7082
rect 24680 7030 24682 7082
rect 24626 7028 24682 7030
rect 24730 7082 24786 7084
rect 24730 7030 24732 7082
rect 24732 7030 24784 7082
rect 24784 7030 24786 7082
rect 24730 7028 24786 7030
rect 24522 5514 24578 5516
rect 24522 5462 24524 5514
rect 24524 5462 24576 5514
rect 24576 5462 24578 5514
rect 24522 5460 24578 5462
rect 24626 5514 24682 5516
rect 24626 5462 24628 5514
rect 24628 5462 24680 5514
rect 24680 5462 24682 5514
rect 24626 5460 24682 5462
rect 24730 5514 24786 5516
rect 24730 5462 24732 5514
rect 24732 5462 24784 5514
rect 24784 5462 24786 5514
rect 24730 5460 24786 5462
rect 25004 8764 25060 8820
rect 25004 7868 25060 7924
rect 25228 9660 25284 9716
rect 25228 8764 25284 8820
rect 25340 8428 25396 8484
rect 25452 9548 25508 9604
rect 25116 6636 25172 6692
rect 25788 9660 25844 9716
rect 25900 8316 25956 8372
rect 25788 8258 25844 8260
rect 25788 8206 25790 8258
rect 25790 8206 25842 8258
rect 25842 8206 25844 8258
rect 25788 8204 25844 8206
rect 25676 6524 25732 6580
rect 25564 4956 25620 5012
rect 24892 4844 24948 4900
rect 26236 12124 26292 12180
rect 26124 11564 26180 11620
rect 26236 11506 26292 11508
rect 26236 11454 26238 11506
rect 26238 11454 26290 11506
rect 26290 11454 26292 11506
rect 26236 11452 26292 11454
rect 26124 9548 26180 9604
rect 27692 12908 27748 12964
rect 26796 12348 26852 12404
rect 26684 11564 26740 11620
rect 27020 11564 27076 11620
rect 26572 8204 26628 8260
rect 26684 10332 26740 10388
rect 26124 7980 26180 8036
rect 24892 4508 24948 4564
rect 24522 3946 24578 3948
rect 24522 3894 24524 3946
rect 24524 3894 24576 3946
rect 24576 3894 24578 3946
rect 24522 3892 24578 3894
rect 24626 3946 24682 3948
rect 24626 3894 24628 3946
rect 24628 3894 24680 3946
rect 24680 3894 24682 3946
rect 24626 3892 24682 3894
rect 24730 3946 24786 3948
rect 24730 3894 24732 3946
rect 24732 3894 24784 3946
rect 24784 3894 24786 3946
rect 24730 3892 24786 3894
rect 24220 3500 24276 3556
rect 23772 1820 23828 1876
rect 25228 3500 25284 3556
rect 25004 3388 25060 3444
rect 24556 1820 24612 1876
rect 27244 11170 27300 11172
rect 27244 11118 27246 11170
rect 27246 11118 27298 11170
rect 27298 11118 27300 11170
rect 27244 11116 27300 11118
rect 27244 10556 27300 10612
rect 27804 12738 27860 12740
rect 27804 12686 27806 12738
rect 27806 12686 27858 12738
rect 27858 12686 27860 12738
rect 27804 12684 27860 12686
rect 28588 14476 28644 14532
rect 28140 14364 28196 14420
rect 28252 14028 28308 14084
rect 29484 16882 29540 16884
rect 29484 16830 29486 16882
rect 29486 16830 29538 16882
rect 29538 16830 29540 16882
rect 29484 16828 29540 16830
rect 29148 16716 29204 16772
rect 29708 16770 29764 16772
rect 29708 16718 29710 16770
rect 29710 16718 29762 16770
rect 29762 16718 29764 16770
rect 29708 16716 29764 16718
rect 29184 15706 29240 15708
rect 29184 15654 29186 15706
rect 29186 15654 29238 15706
rect 29238 15654 29240 15706
rect 29184 15652 29240 15654
rect 29288 15706 29344 15708
rect 29288 15654 29290 15706
rect 29290 15654 29342 15706
rect 29342 15654 29344 15706
rect 29288 15652 29344 15654
rect 29392 15706 29448 15708
rect 29392 15654 29394 15706
rect 29394 15654 29446 15706
rect 29446 15654 29448 15706
rect 29392 15652 29448 15654
rect 29148 15148 29204 15204
rect 29372 14530 29428 14532
rect 29372 14478 29374 14530
rect 29374 14478 29426 14530
rect 29426 14478 29428 14530
rect 29372 14476 29428 14478
rect 28812 14028 28868 14084
rect 29184 14138 29240 14140
rect 29184 14086 29186 14138
rect 29186 14086 29238 14138
rect 29238 14086 29240 14138
rect 29184 14084 29240 14086
rect 29288 14138 29344 14140
rect 29288 14086 29290 14138
rect 29290 14086 29342 14138
rect 29342 14086 29344 14138
rect 29288 14084 29344 14086
rect 29392 14138 29448 14140
rect 29392 14086 29394 14138
rect 29394 14086 29446 14138
rect 29446 14086 29448 14138
rect 29392 14084 29448 14086
rect 29036 13468 29092 13524
rect 30044 13580 30100 13636
rect 28140 12796 28196 12852
rect 29184 12570 29240 12572
rect 29184 12518 29186 12570
rect 29186 12518 29238 12570
rect 29238 12518 29240 12570
rect 29184 12516 29240 12518
rect 29288 12570 29344 12572
rect 29288 12518 29290 12570
rect 29290 12518 29342 12570
rect 29342 12518 29344 12570
rect 29288 12516 29344 12518
rect 29392 12570 29448 12572
rect 29392 12518 29394 12570
rect 29394 12518 29446 12570
rect 29446 12518 29448 12570
rect 29392 12516 29448 12518
rect 29036 12290 29092 12292
rect 29036 12238 29038 12290
rect 29038 12238 29090 12290
rect 29090 12238 29092 12290
rect 29036 12236 29092 12238
rect 27580 11676 27636 11732
rect 27804 11618 27860 11620
rect 27804 11566 27806 11618
rect 27806 11566 27858 11618
rect 27858 11566 27860 11618
rect 27804 11564 27860 11566
rect 28140 11282 28196 11284
rect 28140 11230 28142 11282
rect 28142 11230 28194 11282
rect 28194 11230 28196 11282
rect 28140 11228 28196 11230
rect 29148 11282 29204 11284
rect 29148 11230 29150 11282
rect 29150 11230 29202 11282
rect 29202 11230 29204 11282
rect 29148 11228 29204 11230
rect 30380 13020 30436 13076
rect 27804 11116 27860 11172
rect 27132 10108 27188 10164
rect 27244 9602 27300 9604
rect 27244 9550 27246 9602
rect 27246 9550 27298 9602
rect 27298 9550 27300 9602
rect 27244 9548 27300 9550
rect 27244 8316 27300 8372
rect 26796 7980 26852 8036
rect 27132 8034 27188 8036
rect 27132 7982 27134 8034
rect 27134 7982 27186 8034
rect 27186 7982 27188 8034
rect 27132 7980 27188 7982
rect 25900 3442 25956 3444
rect 25900 3390 25902 3442
rect 25902 3390 25954 3442
rect 25954 3390 25956 3442
rect 25900 3388 25956 3390
rect 26460 3388 26516 3444
rect 25564 924 25620 980
rect 26572 924 26628 980
rect 27468 9212 27524 9268
rect 29184 11002 29240 11004
rect 29184 10950 29186 11002
rect 29186 10950 29238 11002
rect 29238 10950 29240 11002
rect 29184 10948 29240 10950
rect 29288 11002 29344 11004
rect 29288 10950 29290 11002
rect 29290 10950 29342 11002
rect 29342 10950 29344 11002
rect 29288 10948 29344 10950
rect 29392 11002 29448 11004
rect 29392 10950 29394 11002
rect 29394 10950 29446 11002
rect 29446 10950 29448 11002
rect 29392 10948 29448 10950
rect 29148 10556 29204 10612
rect 27804 9660 27860 9716
rect 29184 9434 29240 9436
rect 29184 9382 29186 9434
rect 29186 9382 29238 9434
rect 29238 9382 29240 9434
rect 29184 9380 29240 9382
rect 29288 9434 29344 9436
rect 29288 9382 29290 9434
rect 29290 9382 29342 9434
rect 29342 9382 29344 9434
rect 29288 9380 29344 9382
rect 29392 9434 29448 9436
rect 29392 9382 29394 9434
rect 29394 9382 29446 9434
rect 29446 9382 29448 9434
rect 29392 9380 29448 9382
rect 27580 6748 27636 6804
rect 27468 4844 27524 4900
rect 29184 7866 29240 7868
rect 29184 7814 29186 7866
rect 29186 7814 29238 7866
rect 29238 7814 29240 7866
rect 29184 7812 29240 7814
rect 29288 7866 29344 7868
rect 29288 7814 29290 7866
rect 29290 7814 29342 7866
rect 29342 7814 29344 7866
rect 29288 7812 29344 7814
rect 29392 7866 29448 7868
rect 29392 7814 29394 7866
rect 29394 7814 29446 7866
rect 29446 7814 29448 7866
rect 29392 7812 29448 7814
rect 29184 6298 29240 6300
rect 29184 6246 29186 6298
rect 29186 6246 29238 6298
rect 29238 6246 29240 6298
rect 29184 6244 29240 6246
rect 29288 6298 29344 6300
rect 29288 6246 29290 6298
rect 29290 6246 29342 6298
rect 29342 6246 29344 6298
rect 29288 6244 29344 6246
rect 29392 6298 29448 6300
rect 29392 6246 29394 6298
rect 29394 6246 29446 6298
rect 29446 6246 29448 6298
rect 29392 6244 29448 6246
rect 29184 4730 29240 4732
rect 29184 4678 29186 4730
rect 29186 4678 29238 4730
rect 29238 4678 29240 4730
rect 29184 4676 29240 4678
rect 29288 4730 29344 4732
rect 29288 4678 29290 4730
rect 29290 4678 29342 4730
rect 29342 4678 29344 4730
rect 29288 4676 29344 4678
rect 29392 4730 29448 4732
rect 29392 4678 29394 4730
rect 29394 4678 29446 4730
rect 29446 4678 29448 4730
rect 29392 4676 29448 4678
rect 30044 11116 30100 11172
rect 31276 19010 31332 19012
rect 31276 18958 31278 19010
rect 31278 18958 31330 19010
rect 31330 18958 31332 19010
rect 31276 18956 31332 18958
rect 31052 18450 31108 18452
rect 31052 18398 31054 18450
rect 31054 18398 31106 18450
rect 31106 18398 31108 18450
rect 31052 18396 31108 18398
rect 31388 18338 31444 18340
rect 31388 18286 31390 18338
rect 31390 18286 31442 18338
rect 31442 18286 31444 18338
rect 31388 18284 31444 18286
rect 31612 18226 31668 18228
rect 31612 18174 31614 18226
rect 31614 18174 31666 18226
rect 31666 18174 31668 18226
rect 31612 18172 31668 18174
rect 30828 16716 30884 16772
rect 31276 17388 31332 17444
rect 30828 16156 30884 16212
rect 31500 16770 31556 16772
rect 31500 16718 31502 16770
rect 31502 16718 31554 16770
rect 31554 16718 31556 16770
rect 31500 16716 31556 16718
rect 30716 9772 30772 9828
rect 31276 11116 31332 11172
rect 31164 9714 31220 9716
rect 31164 9662 31166 9714
rect 31166 9662 31218 9714
rect 31218 9662 31220 9714
rect 31164 9660 31220 9662
rect 30604 9212 30660 9268
rect 29932 6636 29988 6692
rect 30604 4956 30660 5012
rect 32396 18396 32452 18452
rect 32508 13580 32564 13636
rect 32620 12684 32676 12740
rect 32284 7532 32340 7588
rect 32396 6524 32452 6580
rect 36092 18620 36148 18676
rect 33846 18058 33902 18060
rect 33846 18006 33848 18058
rect 33848 18006 33900 18058
rect 33900 18006 33902 18058
rect 33846 18004 33902 18006
rect 33950 18058 34006 18060
rect 33950 18006 33952 18058
rect 33952 18006 34004 18058
rect 34004 18006 34006 18058
rect 33950 18004 34006 18006
rect 34054 18058 34110 18060
rect 34054 18006 34056 18058
rect 34056 18006 34108 18058
rect 34108 18006 34110 18058
rect 34054 18004 34110 18006
rect 34860 18060 34916 18116
rect 33846 16490 33902 16492
rect 33846 16438 33848 16490
rect 33848 16438 33900 16490
rect 33900 16438 33902 16490
rect 33846 16436 33902 16438
rect 33950 16490 34006 16492
rect 33950 16438 33952 16490
rect 33952 16438 34004 16490
rect 34004 16438 34006 16490
rect 33950 16436 34006 16438
rect 34054 16490 34110 16492
rect 34054 16438 34056 16490
rect 34056 16438 34108 16490
rect 34108 16438 34110 16490
rect 34054 16436 34110 16438
rect 33516 15820 33572 15876
rect 33846 14922 33902 14924
rect 33846 14870 33848 14922
rect 33848 14870 33900 14922
rect 33900 14870 33902 14922
rect 33846 14868 33902 14870
rect 33950 14922 34006 14924
rect 33950 14870 33952 14922
rect 33952 14870 34004 14922
rect 34004 14870 34006 14922
rect 33950 14868 34006 14870
rect 34054 14922 34110 14924
rect 34054 14870 34056 14922
rect 34056 14870 34108 14922
rect 34108 14870 34110 14922
rect 34054 14868 34110 14870
rect 33846 13354 33902 13356
rect 33846 13302 33848 13354
rect 33848 13302 33900 13354
rect 33900 13302 33902 13354
rect 33846 13300 33902 13302
rect 33950 13354 34006 13356
rect 33950 13302 33952 13354
rect 33952 13302 34004 13354
rect 34004 13302 34006 13354
rect 33950 13300 34006 13302
rect 34054 13354 34110 13356
rect 34054 13302 34056 13354
rect 34056 13302 34108 13354
rect 34108 13302 34110 13354
rect 34054 13300 34110 13302
rect 34524 12684 34580 12740
rect 33846 11786 33902 11788
rect 33846 11734 33848 11786
rect 33848 11734 33900 11786
rect 33900 11734 33902 11786
rect 33846 11732 33902 11734
rect 33950 11786 34006 11788
rect 33950 11734 33952 11786
rect 33952 11734 34004 11786
rect 34004 11734 34006 11786
rect 33950 11732 34006 11734
rect 34054 11786 34110 11788
rect 34054 11734 34056 11786
rect 34056 11734 34108 11786
rect 34108 11734 34110 11786
rect 34054 11732 34110 11734
rect 33516 10668 33572 10724
rect 33846 10218 33902 10220
rect 32956 6076 33012 6132
rect 33068 10108 33124 10164
rect 33846 10166 33848 10218
rect 33848 10166 33900 10218
rect 33900 10166 33902 10218
rect 33846 10164 33902 10166
rect 33950 10218 34006 10220
rect 33950 10166 33952 10218
rect 33952 10166 34004 10218
rect 34004 10166 34006 10218
rect 33950 10164 34006 10166
rect 34054 10218 34110 10220
rect 34054 10166 34056 10218
rect 34056 10166 34108 10218
rect 34108 10166 34110 10218
rect 34054 10164 34110 10166
rect 27244 3442 27300 3444
rect 27244 3390 27246 3442
rect 27246 3390 27298 3442
rect 27298 3390 27300 3442
rect 27244 3388 27300 3390
rect 28252 3388 28308 3444
rect 27580 924 27636 980
rect 29036 3442 29092 3444
rect 29036 3390 29038 3442
rect 29038 3390 29090 3442
rect 29090 3390 29092 3442
rect 29036 3388 29092 3390
rect 29184 3162 29240 3164
rect 29184 3110 29186 3162
rect 29186 3110 29238 3162
rect 29238 3110 29240 3162
rect 29184 3108 29240 3110
rect 29288 3162 29344 3164
rect 29288 3110 29290 3162
rect 29290 3110 29342 3162
rect 29342 3110 29344 3162
rect 29288 3108 29344 3110
rect 29392 3162 29448 3164
rect 29392 3110 29394 3162
rect 29394 3110 29446 3162
rect 29446 3110 29448 3162
rect 29392 3108 29448 3110
rect 28364 924 28420 980
rect 30940 3388 30996 3444
rect 32172 3442 32228 3444
rect 32172 3390 32174 3442
rect 32174 3390 32226 3442
rect 32226 3390 32228 3442
rect 32172 3388 32228 3390
rect 31836 3276 31892 3332
rect 32844 3276 32900 3332
rect 32956 3388 33012 3444
rect 33846 8650 33902 8652
rect 33846 8598 33848 8650
rect 33848 8598 33900 8650
rect 33900 8598 33902 8650
rect 33846 8596 33902 8598
rect 33950 8650 34006 8652
rect 33950 8598 33952 8650
rect 33952 8598 34004 8650
rect 34004 8598 34006 8650
rect 33950 8596 34006 8598
rect 34054 8650 34110 8652
rect 34054 8598 34056 8650
rect 34056 8598 34108 8650
rect 34108 8598 34110 8650
rect 34054 8596 34110 8598
rect 34524 8316 34580 8372
rect 34524 7980 34580 8036
rect 33846 7082 33902 7084
rect 33846 7030 33848 7082
rect 33848 7030 33900 7082
rect 33900 7030 33902 7082
rect 33846 7028 33902 7030
rect 33950 7082 34006 7084
rect 33950 7030 33952 7082
rect 33952 7030 34004 7082
rect 34004 7030 34006 7082
rect 33950 7028 34006 7030
rect 34054 7082 34110 7084
rect 34054 7030 34056 7082
rect 34056 7030 34108 7082
rect 34108 7030 34110 7082
rect 34054 7028 34110 7030
rect 33628 6748 33684 6804
rect 33404 5852 33460 5908
rect 33404 4508 33460 4564
rect 33846 5514 33902 5516
rect 33846 5462 33848 5514
rect 33848 5462 33900 5514
rect 33900 5462 33902 5514
rect 33846 5460 33902 5462
rect 33950 5514 34006 5516
rect 33950 5462 33952 5514
rect 33952 5462 34004 5514
rect 34004 5462 34006 5514
rect 33950 5460 34006 5462
rect 34054 5514 34110 5516
rect 34054 5462 34056 5514
rect 34056 5462 34108 5514
rect 34108 5462 34110 5514
rect 34054 5460 34110 5462
rect 33852 4562 33908 4564
rect 33852 4510 33854 4562
rect 33854 4510 33906 4562
rect 33906 4510 33908 4562
rect 33852 4508 33908 4510
rect 34412 4508 34468 4564
rect 33846 3946 33902 3948
rect 33846 3894 33848 3946
rect 33848 3894 33900 3946
rect 33900 3894 33902 3946
rect 33846 3892 33902 3894
rect 33950 3946 34006 3948
rect 33950 3894 33952 3946
rect 33952 3894 34004 3946
rect 34004 3894 34006 3946
rect 33950 3892 34006 3894
rect 34054 3946 34110 3948
rect 34054 3894 34056 3946
rect 34056 3894 34108 3946
rect 34108 3894 34110 3946
rect 34054 3892 34110 3894
rect 32508 1932 32564 1988
rect 34188 3442 34244 3444
rect 34188 3390 34190 3442
rect 34190 3390 34242 3442
rect 34242 3390 34244 3442
rect 34188 3388 34244 3390
rect 33516 1932 33572 1988
rect 36092 4508 36148 4564
rect 36316 17948 36372 18004
rect 36428 8258 36484 8260
rect 36428 8206 36430 8258
rect 36430 8206 36482 8258
rect 36482 8206 36484 8258
rect 36428 8204 36484 8206
rect 37884 20018 37940 20020
rect 37884 19966 37886 20018
rect 37886 19966 37938 20018
rect 37938 19966 37940 20018
rect 37884 19964 37940 19966
rect 38220 19516 38276 19572
rect 37884 19122 37940 19124
rect 37884 19070 37886 19122
rect 37886 19070 37938 19122
rect 37938 19070 37940 19122
rect 37884 19068 37940 19070
rect 38220 19010 38276 19012
rect 38220 18958 38222 19010
rect 38222 18958 38274 19010
rect 38274 18958 38276 19010
rect 38220 18956 38276 18958
rect 38508 18842 38564 18844
rect 38508 18790 38510 18842
rect 38510 18790 38562 18842
rect 38562 18790 38564 18842
rect 38508 18788 38564 18790
rect 38612 18842 38668 18844
rect 38612 18790 38614 18842
rect 38614 18790 38666 18842
rect 38666 18790 38668 18842
rect 38612 18788 38668 18790
rect 38716 18842 38772 18844
rect 38716 18790 38718 18842
rect 38718 18790 38770 18842
rect 38770 18790 38772 18842
rect 38716 18788 38772 18790
rect 37884 18450 37940 18452
rect 37884 18398 37886 18450
rect 37886 18398 37938 18450
rect 37938 18398 37940 18450
rect 37884 18396 37940 18398
rect 38220 18172 38276 18228
rect 37212 17666 37268 17668
rect 37212 17614 37214 17666
rect 37214 17614 37266 17666
rect 37266 17614 37268 17666
rect 37212 17612 37268 17614
rect 38220 17554 38276 17556
rect 38220 17502 38222 17554
rect 38222 17502 38274 17554
rect 38274 17502 38276 17554
rect 38220 17500 38276 17502
rect 38508 17274 38564 17276
rect 38508 17222 38510 17274
rect 38510 17222 38562 17274
rect 38562 17222 38564 17274
rect 38508 17220 38564 17222
rect 38612 17274 38668 17276
rect 38612 17222 38614 17274
rect 38614 17222 38666 17274
rect 38666 17222 38668 17274
rect 38612 17220 38668 17222
rect 38716 17274 38772 17276
rect 38716 17222 38718 17274
rect 38718 17222 38770 17274
rect 38770 17222 38772 17274
rect 38716 17220 38772 17222
rect 37884 17052 37940 17108
rect 37548 16828 37604 16884
rect 37884 16156 37940 16212
rect 38220 16156 38276 16212
rect 37884 15986 37940 15988
rect 37884 15934 37886 15986
rect 37886 15934 37938 15986
rect 37938 15934 37940 15986
rect 37884 15932 37940 15934
rect 38508 15706 38564 15708
rect 38508 15654 38510 15706
rect 38510 15654 38562 15706
rect 38562 15654 38564 15706
rect 38508 15652 38564 15654
rect 38612 15706 38668 15708
rect 38612 15654 38614 15706
rect 38614 15654 38666 15706
rect 38666 15654 38668 15706
rect 38612 15652 38668 15654
rect 38716 15706 38772 15708
rect 38716 15654 38718 15706
rect 38718 15654 38770 15706
rect 38770 15654 38772 15706
rect 38716 15652 38772 15654
rect 38444 15484 38500 15540
rect 37884 15426 37940 15428
rect 37884 15374 37886 15426
rect 37886 15374 37938 15426
rect 37938 15374 37940 15426
rect 37884 15372 37940 15374
rect 38220 14812 38276 14868
rect 37884 14418 37940 14420
rect 37884 14366 37886 14418
rect 37886 14366 37938 14418
rect 37938 14366 37940 14418
rect 37884 14364 37940 14366
rect 38220 14306 38276 14308
rect 38220 14254 38222 14306
rect 38222 14254 38274 14306
rect 38274 14254 38276 14306
rect 38220 14252 38276 14254
rect 38508 14138 38564 14140
rect 38508 14086 38510 14138
rect 38510 14086 38562 14138
rect 38562 14086 38564 14138
rect 38508 14084 38564 14086
rect 38612 14138 38668 14140
rect 38612 14086 38614 14138
rect 38614 14086 38666 14138
rect 38666 14086 38668 14138
rect 38612 14084 38668 14086
rect 38716 14138 38772 14140
rect 38716 14086 38718 14138
rect 38718 14086 38770 14138
rect 38770 14086 38772 14138
rect 38716 14084 38772 14086
rect 37660 13916 37716 13972
rect 37212 12236 37268 12292
rect 38108 13580 38164 13636
rect 37772 12908 37828 12964
rect 37884 13468 37940 13524
rect 37996 13020 38052 13076
rect 37548 12124 37604 12180
rect 37884 10722 37940 10724
rect 37884 10670 37886 10722
rect 37886 10670 37938 10722
rect 37938 10670 37940 10722
rect 37884 10668 37940 10670
rect 37884 9826 37940 9828
rect 37884 9774 37886 9826
rect 37886 9774 37938 9826
rect 37938 9774 37940 9826
rect 37884 9772 37940 9774
rect 36540 6636 36596 6692
rect 36764 9212 36820 9268
rect 38220 13468 38276 13524
rect 38220 12850 38276 12852
rect 38220 12798 38222 12850
rect 38222 12798 38274 12850
rect 38274 12798 38276 12850
rect 38220 12796 38276 12798
rect 38508 12570 38564 12572
rect 38508 12518 38510 12570
rect 38510 12518 38562 12570
rect 38562 12518 38564 12570
rect 38508 12516 38564 12518
rect 38612 12570 38668 12572
rect 38612 12518 38614 12570
rect 38614 12518 38666 12570
rect 38666 12518 38668 12570
rect 38612 12516 38668 12518
rect 38716 12570 38772 12572
rect 38716 12518 38718 12570
rect 38718 12518 38770 12570
rect 38770 12518 38772 12570
rect 38716 12516 38772 12518
rect 38220 11452 38276 11508
rect 38508 11002 38564 11004
rect 38508 10950 38510 11002
rect 38510 10950 38562 11002
rect 38562 10950 38564 11002
rect 38508 10948 38564 10950
rect 38612 11002 38668 11004
rect 38612 10950 38614 11002
rect 38614 10950 38666 11002
rect 38666 10950 38668 11002
rect 38612 10948 38668 10950
rect 38716 11002 38772 11004
rect 38716 10950 38718 11002
rect 38718 10950 38770 11002
rect 38770 10950 38772 11002
rect 38716 10948 38772 10950
rect 38444 10780 38500 10836
rect 38220 10108 38276 10164
rect 38220 9602 38276 9604
rect 38220 9550 38222 9602
rect 38222 9550 38274 9602
rect 38274 9550 38276 9602
rect 38220 9548 38276 9550
rect 38508 9434 38564 9436
rect 38508 9382 38510 9434
rect 38510 9382 38562 9434
rect 38562 9382 38564 9434
rect 38508 9380 38564 9382
rect 38612 9434 38668 9436
rect 38612 9382 38614 9434
rect 38614 9382 38666 9434
rect 38666 9382 38668 9434
rect 38612 9380 38668 9382
rect 38716 9434 38772 9436
rect 38716 9382 38718 9434
rect 38718 9382 38770 9434
rect 38770 9382 38772 9434
rect 38716 9380 38772 9382
rect 38220 8764 38276 8820
rect 37884 8316 37940 8372
rect 37212 8258 37268 8260
rect 37212 8206 37214 8258
rect 37214 8206 37266 8258
rect 37266 8206 37268 8258
rect 37212 8204 37268 8206
rect 38220 8146 38276 8148
rect 38220 8094 38222 8146
rect 38222 8094 38274 8146
rect 38274 8094 38276 8146
rect 38220 8092 38276 8094
rect 38508 7866 38564 7868
rect 38508 7814 38510 7866
rect 38510 7814 38562 7866
rect 38562 7814 38564 7866
rect 38508 7812 38564 7814
rect 38612 7866 38668 7868
rect 38612 7814 38614 7866
rect 38614 7814 38666 7866
rect 38666 7814 38668 7866
rect 38612 7812 38668 7814
rect 38716 7866 38772 7868
rect 38716 7814 38718 7866
rect 38718 7814 38770 7866
rect 38770 7814 38772 7866
rect 38716 7812 38772 7814
rect 37884 7586 37940 7588
rect 37884 7534 37886 7586
rect 37886 7534 37938 7586
rect 37938 7534 37940 7586
rect 37884 7532 37940 7534
rect 37548 7420 37604 7476
rect 38220 6748 38276 6804
rect 37548 6690 37604 6692
rect 37548 6638 37550 6690
rect 37550 6638 37602 6690
rect 37602 6638 37604 6690
rect 37548 6636 37604 6638
rect 37996 6690 38052 6692
rect 37996 6638 37998 6690
rect 37998 6638 38050 6690
rect 38050 6638 38052 6690
rect 37996 6636 38052 6638
rect 38220 6188 38276 6244
rect 38508 6298 38564 6300
rect 38508 6246 38510 6298
rect 38510 6246 38562 6298
rect 38562 6246 38564 6298
rect 38508 6244 38564 6246
rect 38612 6298 38668 6300
rect 38612 6246 38614 6298
rect 38614 6246 38666 6298
rect 38666 6246 38668 6298
rect 38612 6244 38668 6246
rect 38716 6298 38772 6300
rect 38716 6246 38718 6298
rect 38718 6246 38770 6298
rect 38770 6246 38772 6298
rect 38716 6244 38772 6246
rect 37660 6130 37716 6132
rect 37660 6078 37662 6130
rect 37662 6078 37714 6130
rect 37714 6078 37716 6130
rect 37660 6076 37716 6078
rect 38220 5404 38276 5460
rect 36764 5180 36820 5236
rect 37548 5234 37604 5236
rect 37548 5182 37550 5234
rect 37550 5182 37602 5234
rect 37602 5182 37604 5234
rect 37548 5180 37604 5182
rect 37996 5180 38052 5236
rect 38220 4898 38276 4900
rect 38220 4846 38222 4898
rect 38222 4846 38274 4898
rect 38274 4846 38276 4898
rect 38220 4844 38276 4846
rect 38508 4730 38564 4732
rect 38508 4678 38510 4730
rect 38510 4678 38562 4730
rect 38562 4678 38564 4730
rect 38508 4676 38564 4678
rect 38612 4730 38668 4732
rect 38612 4678 38614 4730
rect 38614 4678 38666 4730
rect 38666 4678 38668 4730
rect 38612 4676 38668 4678
rect 38716 4730 38772 4732
rect 38716 4678 38718 4730
rect 38718 4678 38770 4730
rect 38770 4678 38772 4730
rect 38716 4676 38772 4678
rect 37660 4562 37716 4564
rect 37660 4510 37662 4562
rect 37662 4510 37714 4562
rect 37714 4510 37716 4562
rect 37660 4508 37716 4510
rect 38220 4060 38276 4116
rect 36316 3612 36372 3668
rect 37548 3666 37604 3668
rect 37548 3614 37550 3666
rect 37550 3614 37602 3666
rect 37602 3614 37604 3666
rect 37548 3612 37604 3614
rect 37996 3612 38052 3668
rect 38220 3442 38276 3444
rect 38220 3390 38222 3442
rect 38222 3390 38274 3442
rect 38274 3390 38276 3442
rect 38220 3388 38276 3390
rect 38508 3162 38564 3164
rect 38508 3110 38510 3162
rect 38510 3110 38562 3162
rect 38562 3110 38564 3162
rect 38508 3108 38564 3110
rect 38612 3162 38668 3164
rect 38612 3110 38614 3162
rect 38614 3110 38666 3162
rect 38666 3110 38668 3162
rect 38612 3108 38668 3110
rect 38716 3162 38772 3164
rect 38716 3110 38718 3162
rect 38718 3110 38770 3162
rect 38770 3110 38772 3162
rect 38716 3108 38772 3110
<< metal3 >>
rect 24882 36876 24892 36932
rect 24948 36876 25900 36932
rect 25956 36876 25966 36932
rect 26226 36876 26236 36932
rect 26292 36876 27244 36932
rect 27300 36876 27310 36932
rect 31602 36876 31612 36932
rect 31668 36876 32844 36932
rect 32900 36876 32910 36932
rect 36306 36876 36316 36932
rect 36372 36876 37324 36932
rect 37380 36876 37390 36932
rect 5864 36820 5874 36876
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 6138 36820 6148 36876
rect 15188 36820 15198 36876
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15462 36820 15472 36876
rect 24512 36820 24522 36876
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24786 36820 24796 36876
rect 33836 36820 33846 36876
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 34110 36820 34120 36876
rect 24210 36652 24220 36708
rect 24276 36652 25228 36708
rect 25284 36652 25294 36708
rect 26852 36428 27468 36484
rect 27524 36428 27534 36484
rect 16034 36316 16044 36372
rect 16100 36316 18620 36372
rect 18676 36316 18686 36372
rect 20738 36316 20748 36372
rect 20804 36316 22092 36372
rect 22148 36316 22158 36372
rect 23538 36316 23548 36372
rect 23604 36316 26236 36372
rect 26292 36316 26302 36372
rect 26786 36204 26796 36260
rect 26852 36204 26908 36428
rect 27682 36316 27692 36372
rect 27748 36316 28700 36372
rect 28756 36316 28766 36372
rect 31154 36316 31164 36372
rect 31220 36316 32172 36372
rect 32228 36316 32238 36372
rect 32946 36316 32956 36372
rect 33012 36316 34188 36372
rect 34244 36316 34254 36372
rect 34962 36316 34972 36372
rect 35028 36316 35980 36372
rect 36036 36316 36046 36372
rect 28466 36204 28476 36260
rect 28532 36204 29036 36260
rect 29092 36204 29102 36260
rect 29810 36204 29820 36260
rect 29876 36204 30380 36260
rect 30436 36204 30446 36260
rect 33740 36092 34412 36148
rect 34468 36092 34478 36148
rect 10526 36036 10536 36092
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10800 36036 10810 36092
rect 19850 36036 19860 36092
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 20124 36036 20134 36092
rect 29174 36036 29184 36092
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29448 36036 29458 36092
rect 33740 35924 33796 36092
rect 38498 36036 38508 36092
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38772 36036 38782 36092
rect 24994 35868 25004 35924
rect 25060 35868 33740 35924
rect 33796 35868 33806 35924
rect 9986 35756 9996 35812
rect 10052 35756 17388 35812
rect 17444 35756 17454 35812
rect 39200 35700 40000 35728
rect 37538 35644 37548 35700
rect 37604 35644 40000 35700
rect 39200 35616 40000 35644
rect 9762 35532 9772 35588
rect 9828 35532 10444 35588
rect 10500 35532 17724 35588
rect 17780 35532 17790 35588
rect 23986 35532 23996 35588
rect 24052 35532 33180 35588
rect 33236 35532 33852 35588
rect 33908 35532 33918 35588
rect 22418 35420 22428 35476
rect 22484 35420 35308 35476
rect 35364 35420 35374 35476
rect 27570 35308 27580 35364
rect 27636 35308 30716 35364
rect 30772 35308 30782 35364
rect 34402 35308 34412 35364
rect 34468 35308 37884 35364
rect 37940 35308 37950 35364
rect 5864 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6148 35308
rect 15188 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15472 35308
rect 24512 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24796 35308
rect 33836 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34120 35308
rect 39200 35028 40000 35056
rect 38210 34972 38220 35028
rect 38276 34972 40000 35028
rect 39200 34944 40000 34972
rect 31490 34748 31500 34804
rect 31556 34748 37660 34804
rect 37716 34748 37726 34804
rect 10526 34468 10536 34524
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10800 34468 10810 34524
rect 19850 34468 19860 34524
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 20124 34468 20134 34524
rect 29174 34468 29184 34524
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29448 34468 29458 34524
rect 38498 34468 38508 34524
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38772 34468 38782 34524
rect 39200 34356 40000 34384
rect 38434 34300 38444 34356
rect 38500 34300 40000 34356
rect 39200 34272 40000 34300
rect 36082 33964 36092 34020
rect 36148 33964 37548 34020
rect 37604 33964 37996 34020
rect 38052 33964 38062 34020
rect 23426 33852 23436 33908
rect 23492 33852 24892 33908
rect 24948 33852 24958 33908
rect 10322 33740 10332 33796
rect 10388 33740 14140 33796
rect 14196 33740 14206 33796
rect 5864 33684 5874 33740
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 6138 33684 6148 33740
rect 15188 33684 15198 33740
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15462 33684 15472 33740
rect 24512 33684 24522 33740
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24786 33684 24796 33740
rect 33836 33684 33846 33740
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 34110 33684 34120 33740
rect 39200 33684 40000 33712
rect 11666 33628 11676 33684
rect 11732 33628 13692 33684
rect 13748 33628 13758 33684
rect 26450 33628 26460 33684
rect 26516 33628 32284 33684
rect 32340 33628 32350 33684
rect 38210 33628 38220 33684
rect 38276 33628 40000 33684
rect 39200 33600 40000 33628
rect 25778 33516 25788 33572
rect 25844 33516 27356 33572
rect 27412 33516 27422 33572
rect 28242 33516 28252 33572
rect 28308 33516 30044 33572
rect 30100 33516 30110 33572
rect 21746 33068 21756 33124
rect 21812 33068 22652 33124
rect 22708 33068 22718 33124
rect 23650 33068 23660 33124
rect 23716 33068 25452 33124
rect 25508 33068 25518 33124
rect 32162 33068 32172 33124
rect 32228 33068 37660 33124
rect 37716 33068 37726 33124
rect 38210 33068 38220 33124
rect 38276 33068 38948 33124
rect 0 33012 800 33040
rect 38892 33012 38948 33068
rect 39200 33012 40000 33040
rect 0 32956 1708 33012
rect 1764 32956 2492 33012
rect 2548 32956 2558 33012
rect 38892 32956 40000 33012
rect 0 32928 800 32956
rect 10526 32900 10536 32956
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10800 32900 10810 32956
rect 19850 32900 19860 32956
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 20124 32900 20134 32956
rect 29174 32900 29184 32956
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29448 32900 29458 32956
rect 38498 32900 38508 32956
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38772 32900 38782 32956
rect 39200 32928 40000 32956
rect 26338 32508 26348 32564
rect 26404 32508 37548 32564
rect 37604 32508 37996 32564
rect 38052 32508 38062 32564
rect 0 32340 800 32368
rect 39200 32340 40000 32368
rect 0 32284 1708 32340
rect 1764 32284 1774 32340
rect 38210 32284 38220 32340
rect 38276 32284 40000 32340
rect 0 32256 800 32284
rect 39200 32256 40000 32284
rect 5864 32116 5874 32172
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 6138 32116 6148 32172
rect 15188 32116 15198 32172
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15462 32116 15472 32172
rect 24512 32116 24522 32172
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24786 32116 24796 32172
rect 33836 32116 33846 32172
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 34110 32116 34120 32172
rect 17938 31836 17948 31892
rect 18004 31836 18732 31892
rect 18788 31836 18798 31892
rect 0 31668 800 31696
rect 39200 31668 40000 31696
rect 0 31612 2380 31668
rect 2436 31612 2446 31668
rect 30370 31612 30380 31668
rect 30436 31612 37212 31668
rect 37268 31612 37278 31668
rect 37538 31612 37548 31668
rect 37604 31612 40000 31668
rect 0 31584 800 31612
rect 39200 31584 40000 31612
rect 1698 31500 1708 31556
rect 1764 31500 1774 31556
rect 2706 31500 2716 31556
rect 2772 31500 3276 31556
rect 3332 31500 9324 31556
rect 9380 31500 9390 31556
rect 0 30996 800 31024
rect 1708 30996 1764 31500
rect 10526 31332 10536 31388
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10800 31332 10810 31388
rect 19850 31332 19860 31388
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 20124 31332 20134 31388
rect 29174 31332 29184 31388
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29448 31332 29458 31388
rect 38498 31332 38508 31388
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38772 31332 38782 31388
rect 32946 31164 32956 31220
rect 33012 31164 37884 31220
rect 37940 31164 37950 31220
rect 39200 30996 40000 31024
rect 0 30940 1764 30996
rect 28802 30940 28812 30996
rect 28868 30940 37884 30996
rect 37940 30940 37950 30996
rect 38434 30940 38444 30996
rect 38500 30940 40000 30996
rect 0 30912 800 30940
rect 39200 30912 40000 30940
rect 1922 30828 1932 30884
rect 1988 30828 2492 30884
rect 2548 30828 6860 30884
rect 6916 30828 6926 30884
rect 5864 30548 5874 30604
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 6138 30548 6148 30604
rect 15188 30548 15198 30604
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15462 30548 15472 30604
rect 24512 30548 24522 30604
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24786 30548 24796 30604
rect 33836 30548 33846 30604
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 34110 30548 34120 30604
rect 24322 30380 24332 30436
rect 24388 30380 37100 30436
rect 37156 30380 37166 30436
rect 0 30324 800 30352
rect 39200 30324 40000 30352
rect 0 30268 1708 30324
rect 1764 30268 1774 30324
rect 29922 30268 29932 30324
rect 29988 30268 34412 30324
rect 34468 30268 34478 30324
rect 38210 30268 38220 30324
rect 38276 30268 40000 30324
rect 0 30240 800 30268
rect 39200 30240 40000 30268
rect 7858 30156 7868 30212
rect 7924 30156 11564 30212
rect 11620 30156 11630 30212
rect 14354 30156 14364 30212
rect 14420 30156 15596 30212
rect 15652 30156 15662 30212
rect 3602 30044 3612 30100
rect 3668 30044 10108 30100
rect 10164 30044 10174 30100
rect 12226 30044 12236 30100
rect 12292 30044 14812 30100
rect 14868 30044 14878 30100
rect 32386 30044 32396 30100
rect 32452 30044 37884 30100
rect 37940 30044 37950 30100
rect 1698 29932 1708 29988
rect 1764 29932 1774 29988
rect 18386 29932 18396 29988
rect 18452 29932 19292 29988
rect 19348 29932 19358 29988
rect 1708 29764 1764 29932
rect 10526 29764 10536 29820
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10800 29764 10810 29820
rect 19850 29764 19860 29820
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 20124 29764 20134 29820
rect 29174 29764 29184 29820
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29448 29764 29458 29820
rect 38498 29764 38508 29820
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38772 29764 38782 29820
rect 924 29708 1764 29764
rect 26114 29708 26124 29764
rect 26180 29708 26796 29764
rect 26852 29708 26862 29764
rect 38210 29708 38220 29764
rect 38276 29708 38286 29764
rect 0 29652 800 29680
rect 924 29652 980 29708
rect 38220 29652 38276 29708
rect 39200 29652 40000 29680
rect 0 29596 980 29652
rect 19618 29596 19628 29652
rect 19684 29596 21980 29652
rect 22036 29596 22046 29652
rect 38220 29596 40000 29652
rect 0 29568 800 29596
rect 39200 29568 40000 29596
rect 6626 29484 6636 29540
rect 6692 29484 16940 29540
rect 16996 29484 17006 29540
rect 17948 29484 19516 29540
rect 19572 29484 19964 29540
rect 20020 29484 20030 29540
rect 17948 29428 18004 29484
rect 6738 29372 6748 29428
rect 6804 29372 15820 29428
rect 15876 29372 16716 29428
rect 16772 29372 17388 29428
rect 17444 29372 17948 29428
rect 18004 29372 18014 29428
rect 18498 29372 18508 29428
rect 18564 29372 19292 29428
rect 19348 29372 19358 29428
rect 22418 29372 22428 29428
rect 22484 29372 26908 29428
rect 30258 29372 30268 29428
rect 30324 29372 37884 29428
rect 37940 29372 37950 29428
rect 26852 29316 26908 29372
rect 2034 29260 2044 29316
rect 2100 29260 2492 29316
rect 2548 29260 4060 29316
rect 4116 29260 4126 29316
rect 4274 29260 4284 29316
rect 4340 29260 15372 29316
rect 15428 29260 16268 29316
rect 16324 29260 16548 29316
rect 20290 29260 20300 29316
rect 20356 29260 21868 29316
rect 21924 29260 22764 29316
rect 22820 29260 26572 29316
rect 26628 29260 26638 29316
rect 26852 29260 27468 29316
rect 27524 29260 27534 29316
rect 16492 29204 16548 29260
rect 13682 29148 13692 29204
rect 13748 29148 15036 29204
rect 15092 29148 16156 29204
rect 16212 29148 16222 29204
rect 16482 29148 16492 29204
rect 16548 29148 17948 29204
rect 18004 29148 18396 29204
rect 18452 29148 18462 29204
rect 21186 29148 21196 29204
rect 21252 29148 22204 29204
rect 22260 29148 22988 29204
rect 23044 29148 23884 29204
rect 23940 29148 23950 29204
rect 25442 29148 25452 29204
rect 25508 29148 26796 29204
rect 26852 29148 27356 29204
rect 27412 29148 27692 29204
rect 27748 29148 27758 29204
rect 0 28980 800 29008
rect 5864 28980 5874 29036
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 6138 28980 6148 29036
rect 15188 28980 15198 29036
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15462 28980 15472 29036
rect 24512 28980 24522 29036
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24786 28980 24796 29036
rect 33836 28980 33846 29036
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 34110 28980 34120 29036
rect 39200 28980 40000 29008
rect 0 28924 1708 28980
rect 1764 28924 1774 28980
rect 38210 28924 38220 28980
rect 38276 28924 40000 28980
rect 0 28896 800 28924
rect 39200 28896 40000 28924
rect 15092 28812 15820 28868
rect 15876 28812 16604 28868
rect 16660 28812 16670 28868
rect 15092 28756 15148 28812
rect 12674 28700 12684 28756
rect 12740 28700 13916 28756
rect 13972 28700 15148 28756
rect 13122 28588 13132 28644
rect 13188 28588 13580 28644
rect 13636 28588 13646 28644
rect 13794 28588 13804 28644
rect 13860 28588 14252 28644
rect 14308 28588 14318 28644
rect 17266 28588 17276 28644
rect 17332 28588 19012 28644
rect 2034 28476 2044 28532
rect 2100 28476 12348 28532
rect 12404 28476 12414 28532
rect 18956 28420 19012 28588
rect 23314 28476 23324 28532
rect 23380 28476 24780 28532
rect 24836 28476 24846 28532
rect 25890 28476 25900 28532
rect 25956 28476 31388 28532
rect 31444 28476 31454 28532
rect 1698 28364 1708 28420
rect 1764 28364 1774 28420
rect 11554 28364 11564 28420
rect 11620 28364 14700 28420
rect 14756 28364 14766 28420
rect 18946 28364 18956 28420
rect 19012 28364 19022 28420
rect 38210 28364 38220 28420
rect 38276 28364 38948 28420
rect 0 28308 800 28336
rect 1708 28308 1764 28364
rect 0 28252 1764 28308
rect 38892 28308 38948 28364
rect 39200 28308 40000 28336
rect 38892 28252 40000 28308
rect 0 28224 800 28252
rect 10526 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10810 28252
rect 19850 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20134 28252
rect 29174 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29458 28252
rect 38498 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38782 28252
rect 39200 28224 40000 28252
rect 14802 28028 14812 28084
rect 14868 28028 15708 28084
rect 15764 28028 16156 28084
rect 16212 28028 16222 28084
rect 23174 28028 23212 28084
rect 23268 28028 23278 28084
rect 8418 27916 8428 27972
rect 8484 27916 15596 27972
rect 15652 27916 15662 27972
rect 17490 27916 17500 27972
rect 17556 27916 17948 27972
rect 18004 27916 18014 27972
rect 20514 27916 20524 27972
rect 20580 27916 20972 27972
rect 21028 27916 21980 27972
rect 22036 27916 25452 27972
rect 25508 27916 25518 27972
rect 2034 27804 2044 27860
rect 2100 27804 9436 27860
rect 9492 27804 9502 27860
rect 22642 27804 22652 27860
rect 22708 27804 23884 27860
rect 23940 27804 23950 27860
rect 24098 27804 24108 27860
rect 24164 27804 25340 27860
rect 25396 27804 26460 27860
rect 26516 27804 26526 27860
rect 26674 27804 26684 27860
rect 26740 27804 27804 27860
rect 27860 27804 27870 27860
rect 16818 27692 16828 27748
rect 16884 27692 17500 27748
rect 17556 27692 18172 27748
rect 18228 27692 20188 27748
rect 20244 27692 20254 27748
rect 30482 27692 30492 27748
rect 30548 27692 37548 27748
rect 37604 27692 37996 27748
rect 38052 27692 38062 27748
rect 0 27636 800 27664
rect 39200 27636 40000 27664
rect 0 27580 1708 27636
rect 1764 27580 1774 27636
rect 11666 27580 11676 27636
rect 11732 27580 13580 27636
rect 13636 27580 15932 27636
rect 15988 27580 17388 27636
rect 17444 27580 17454 27636
rect 38210 27580 38220 27636
rect 38276 27580 40000 27636
rect 0 27552 800 27580
rect 39200 27552 40000 27580
rect 17826 27468 17836 27524
rect 17892 27468 18060 27524
rect 18116 27468 18126 27524
rect 5864 27412 5874 27468
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 6138 27412 6148 27468
rect 15188 27412 15198 27468
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15462 27412 15472 27468
rect 24512 27412 24522 27468
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24786 27412 24796 27468
rect 33836 27412 33846 27468
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 34110 27412 34120 27468
rect 10098 27356 10108 27412
rect 10164 27356 13580 27412
rect 13636 27356 13646 27412
rect 10434 27244 10444 27300
rect 10500 27244 15036 27300
rect 15092 27244 15102 27300
rect 19730 27244 19740 27300
rect 19796 27244 35756 27300
rect 35812 27244 35822 27300
rect 29922 27132 29932 27188
rect 29988 27132 37212 27188
rect 37268 27132 37278 27188
rect 4162 27020 4172 27076
rect 4228 27020 15372 27076
rect 15428 27020 15438 27076
rect 17826 27020 17836 27076
rect 17892 27020 18508 27076
rect 18564 27020 18574 27076
rect 22306 27020 22316 27076
rect 22372 27020 22876 27076
rect 22932 27020 22942 27076
rect 24098 27020 24108 27076
rect 24164 27020 24668 27076
rect 24724 27020 24734 27076
rect 25330 27020 25340 27076
rect 25396 27020 26460 27076
rect 26516 27020 26526 27076
rect 37538 27020 37548 27076
rect 37604 27020 39060 27076
rect 0 26964 800 26992
rect 39004 26964 39060 27020
rect 39200 26964 40000 26992
rect 0 26908 2380 26964
rect 2436 26908 2446 26964
rect 2706 26908 2716 26964
rect 2772 26908 6748 26964
rect 6804 26908 6814 26964
rect 17350 26908 17388 26964
rect 17444 26908 17454 26964
rect 17602 26908 17612 26964
rect 17668 26908 18396 26964
rect 18452 26908 18462 26964
rect 35298 26908 35308 26964
rect 35364 26908 37884 26964
rect 37940 26908 37950 26964
rect 39004 26908 40000 26964
rect 0 26880 800 26908
rect 39200 26880 40000 26908
rect 10210 26796 10220 26852
rect 10276 26796 10892 26852
rect 10948 26796 10958 26852
rect 16146 26796 16156 26852
rect 16212 26796 17948 26852
rect 18004 26796 20412 26852
rect 20468 26796 20478 26852
rect 29698 26796 29708 26852
rect 29764 26796 30380 26852
rect 30436 26796 30446 26852
rect 10526 26628 10536 26684
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10800 26628 10810 26684
rect 19850 26628 19860 26684
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 20124 26628 20134 26684
rect 29174 26628 29184 26684
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29448 26628 29458 26684
rect 38498 26628 38508 26684
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38772 26628 38782 26684
rect 16258 26572 16268 26628
rect 16324 26572 17948 26628
rect 18004 26572 18014 26628
rect 7074 26460 7084 26516
rect 7140 26460 14476 26516
rect 14532 26460 14542 26516
rect 15698 26460 15708 26516
rect 15764 26460 16604 26516
rect 16660 26460 16670 26516
rect 24210 26460 24220 26516
rect 24276 26460 33068 26516
rect 33124 26460 33134 26516
rect 10668 26348 15148 26404
rect 15586 26348 15596 26404
rect 15652 26348 17164 26404
rect 17220 26348 17500 26404
rect 17556 26348 17566 26404
rect 19170 26348 19180 26404
rect 19236 26348 20076 26404
rect 20132 26348 20142 26404
rect 21970 26348 21980 26404
rect 22036 26348 23660 26404
rect 23716 26348 24892 26404
rect 24948 26348 24958 26404
rect 0 26292 800 26320
rect 10668 26292 10724 26348
rect 15092 26292 15148 26348
rect 39200 26292 40000 26320
rect 0 26236 1820 26292
rect 1876 26236 1886 26292
rect 9650 26236 9660 26292
rect 9716 26236 10668 26292
rect 10724 26236 10734 26292
rect 14130 26236 14140 26292
rect 14196 26236 14700 26292
rect 14756 26236 14766 26292
rect 15092 26236 19740 26292
rect 19796 26236 19806 26292
rect 21298 26236 21308 26292
rect 21364 26236 23772 26292
rect 23828 26236 23838 26292
rect 38098 26236 38108 26292
rect 38164 26236 40000 26292
rect 0 26208 800 26236
rect 19740 26180 19796 26236
rect 39200 26208 40000 26236
rect 3042 26124 3052 26180
rect 3108 26124 8428 26180
rect 11554 26124 11564 26180
rect 11620 26124 13804 26180
rect 13860 26124 15708 26180
rect 15764 26124 15774 26180
rect 19740 26124 21196 26180
rect 21252 26124 21262 26180
rect 8372 26068 8428 26124
rect 8372 26012 15820 26068
rect 15876 26012 15886 26068
rect 16258 26012 16268 26068
rect 16324 26012 16940 26068
rect 16996 26012 19516 26068
rect 19572 26012 19582 26068
rect 20290 26012 20300 26068
rect 20356 26012 21420 26068
rect 21476 26012 21486 26068
rect 27010 26012 27020 26068
rect 27076 26012 34188 26068
rect 34244 26012 34254 26068
rect 5864 25844 5874 25900
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 6138 25844 6148 25900
rect 15188 25844 15198 25900
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15462 25844 15472 25900
rect 24512 25844 24522 25900
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24786 25844 24796 25900
rect 33836 25844 33846 25900
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 34110 25844 34120 25900
rect 14690 25788 14700 25844
rect 14756 25788 15036 25844
rect 15092 25788 15102 25844
rect 16380 25788 19852 25844
rect 19908 25788 21420 25844
rect 21476 25788 21486 25844
rect 16380 25732 16436 25788
rect 9762 25676 9772 25732
rect 9828 25676 16436 25732
rect 16594 25676 16604 25732
rect 16660 25676 18956 25732
rect 19012 25676 22764 25732
rect 22820 25676 22830 25732
rect 23314 25676 23324 25732
rect 23380 25676 24108 25732
rect 24164 25676 24174 25732
rect 0 25620 800 25648
rect 39200 25620 40000 25648
rect 0 25564 1708 25620
rect 1764 25564 1774 25620
rect 2034 25564 2044 25620
rect 2100 25564 13020 25620
rect 13076 25564 13086 25620
rect 14018 25564 14028 25620
rect 14084 25564 14476 25620
rect 14532 25564 14924 25620
rect 14980 25564 14990 25620
rect 17938 25564 17948 25620
rect 18004 25564 18844 25620
rect 18900 25564 18910 25620
rect 27570 25564 27580 25620
rect 27636 25564 27646 25620
rect 38210 25564 38220 25620
rect 38276 25564 40000 25620
rect 0 25536 800 25564
rect 27580 25508 27636 25564
rect 39200 25536 40000 25564
rect 11554 25452 11564 25508
rect 11620 25452 12684 25508
rect 12740 25452 14980 25508
rect 15138 25452 15148 25508
rect 15204 25452 16604 25508
rect 16660 25452 16670 25508
rect 16930 25452 16940 25508
rect 16996 25452 17388 25508
rect 17444 25452 17454 25508
rect 20066 25452 20076 25508
rect 20132 25452 24444 25508
rect 24500 25452 26796 25508
rect 26852 25452 27636 25508
rect 14924 25396 14980 25452
rect 12786 25340 12796 25396
rect 12852 25340 13356 25396
rect 13412 25340 13422 25396
rect 14924 25340 17612 25396
rect 17668 25340 17678 25396
rect 20178 25340 20188 25396
rect 20244 25340 21308 25396
rect 21364 25340 21374 25396
rect 28018 25340 28028 25396
rect 28084 25340 37660 25396
rect 37716 25340 37726 25396
rect 2258 25228 2268 25284
rect 2324 25228 11452 25284
rect 11508 25228 11518 25284
rect 14354 25228 14364 25284
rect 14420 25228 15148 25284
rect 15204 25228 15214 25284
rect 15810 25228 15820 25284
rect 15876 25228 16380 25284
rect 16436 25228 16716 25284
rect 16772 25228 20076 25284
rect 20132 25228 20142 25284
rect 38210 25228 38220 25284
rect 38276 25228 38286 25284
rect 2818 25116 2828 25172
rect 2884 25116 5068 25172
rect 5124 25116 5134 25172
rect 6514 25116 6524 25172
rect 6580 25116 6972 25172
rect 7028 25116 7038 25172
rect 12450 25116 12460 25172
rect 12516 25116 17724 25172
rect 17780 25116 17948 25172
rect 18004 25116 18014 25172
rect 22418 25116 22428 25172
rect 22484 25116 22876 25172
rect 22932 25116 22942 25172
rect 10526 25060 10536 25116
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10800 25060 10810 25116
rect 19850 25060 19860 25116
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 20124 25060 20134 25116
rect 29174 25060 29184 25116
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29448 25060 29458 25116
rect 1698 25004 1708 25060
rect 1764 25004 1774 25060
rect 15092 25004 15932 25060
rect 15988 25004 16492 25060
rect 16548 25004 16558 25060
rect 0 24948 800 24976
rect 1708 24948 1764 25004
rect 0 24892 1764 24948
rect 0 24864 800 24892
rect 2034 24780 2044 24836
rect 2100 24780 10220 24836
rect 10276 24780 10286 24836
rect 15092 24724 15148 25004
rect 38220 24948 38276 25228
rect 38498 25060 38508 25116
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38772 25060 38782 25116
rect 39200 24948 40000 24976
rect 16258 24892 16268 24948
rect 16324 24892 17388 24948
rect 17444 24892 17454 24948
rect 22418 24892 22428 24948
rect 22484 24892 23212 24948
rect 23268 24892 23278 24948
rect 26786 24892 26796 24948
rect 26852 24892 27132 24948
rect 27188 24892 27198 24948
rect 38220 24892 40000 24948
rect 39200 24864 40000 24892
rect 16034 24780 16044 24836
rect 16100 24780 16828 24836
rect 16884 24780 16894 24836
rect 24658 24780 24668 24836
rect 24724 24780 35308 24836
rect 35364 24780 35374 24836
rect 11666 24668 11676 24724
rect 11732 24668 12572 24724
rect 12628 24668 13804 24724
rect 13860 24668 13870 24724
rect 14242 24668 14252 24724
rect 14308 24668 15148 24724
rect 16044 24612 16100 24780
rect 17154 24668 17164 24724
rect 17220 24668 17612 24724
rect 17668 24668 17678 24724
rect 18918 24668 18956 24724
rect 19012 24668 19022 24724
rect 24434 24668 24444 24724
rect 24500 24668 25228 24724
rect 25284 24668 25294 24724
rect 31266 24668 31276 24724
rect 31332 24668 37884 24724
rect 37940 24668 37950 24724
rect 14354 24556 14364 24612
rect 14420 24556 16100 24612
rect 18386 24556 18396 24612
rect 18452 24556 20188 24612
rect 20244 24556 20254 24612
rect 20962 24556 20972 24612
rect 21028 24556 25788 24612
rect 25844 24556 26572 24612
rect 26628 24556 28140 24612
rect 28196 24556 28206 24612
rect 31892 24556 36316 24612
rect 36372 24556 36382 24612
rect 14018 24444 14028 24500
rect 14084 24444 14700 24500
rect 14756 24444 18284 24500
rect 18340 24444 19180 24500
rect 19236 24444 19246 24500
rect 21186 24444 21196 24500
rect 21252 24444 21980 24500
rect 22036 24444 22046 24500
rect 24322 24444 24332 24500
rect 24388 24444 25564 24500
rect 25620 24444 25630 24500
rect 31892 24388 31948 24556
rect 17378 24332 17388 24388
rect 17444 24332 17612 24388
rect 17668 24332 17678 24388
rect 22838 24332 22876 24388
rect 22932 24332 22942 24388
rect 25218 24332 25228 24388
rect 25284 24332 31948 24388
rect 0 24276 800 24304
rect 5864 24276 5874 24332
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 6138 24276 6148 24332
rect 15188 24276 15198 24332
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15462 24276 15472 24332
rect 24512 24276 24522 24332
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24786 24276 24796 24332
rect 33836 24276 33846 24332
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 34110 24276 34120 24332
rect 39200 24276 40000 24304
rect 0 24220 1708 24276
rect 1764 24220 1774 24276
rect 25666 24220 25676 24276
rect 25732 24220 26796 24276
rect 26852 24220 26862 24276
rect 38210 24220 38220 24276
rect 38276 24220 40000 24276
rect 0 24192 800 24220
rect 39200 24192 40000 24220
rect 27794 24108 27804 24164
rect 27860 24108 37772 24164
rect 37828 24108 37838 24164
rect 11778 23996 11788 24052
rect 11844 23996 12348 24052
rect 12404 23996 12414 24052
rect 18946 23996 18956 24052
rect 19012 23996 22204 24052
rect 22260 23996 23324 24052
rect 23380 23996 23390 24052
rect 10434 23884 10444 23940
rect 10500 23884 12572 23940
rect 12628 23884 12638 23940
rect 12786 23884 12796 23940
rect 12852 23884 13244 23940
rect 13300 23884 13804 23940
rect 13860 23884 13870 23940
rect 14578 23884 14588 23940
rect 14644 23884 17388 23940
rect 17444 23884 18172 23940
rect 18228 23884 18238 23940
rect 21186 23884 21196 23940
rect 21252 23884 24220 23940
rect 24276 23884 26572 23940
rect 26628 23884 26908 23940
rect 8372 23772 14364 23828
rect 14420 23772 14430 23828
rect 16482 23772 16492 23828
rect 16548 23772 17724 23828
rect 17780 23772 17790 23828
rect 21634 23772 21644 23828
rect 21700 23772 22988 23828
rect 23044 23772 23054 23828
rect 8372 23716 8428 23772
rect 1698 23660 1708 23716
rect 1764 23660 1774 23716
rect 2146 23660 2156 23716
rect 2212 23660 8428 23716
rect 18946 23660 18956 23716
rect 19012 23660 22652 23716
rect 22708 23660 23100 23716
rect 23156 23660 23166 23716
rect 0 23604 800 23632
rect 1708 23604 1764 23660
rect 26852 23604 26908 23884
rect 28466 23772 28476 23828
rect 28532 23772 29148 23828
rect 29204 23772 29214 23828
rect 35298 23772 35308 23828
rect 35364 23772 37884 23828
rect 37940 23772 37950 23828
rect 38210 23660 38220 23716
rect 38276 23660 38948 23716
rect 38892 23604 38948 23660
rect 39200 23604 40000 23632
rect 0 23548 1764 23604
rect 19254 23548 19292 23604
rect 19348 23548 19358 23604
rect 22306 23548 22316 23604
rect 22372 23548 23212 23604
rect 23268 23548 23548 23604
rect 23604 23548 23614 23604
rect 26852 23548 27916 23604
rect 27972 23548 27982 23604
rect 38892 23548 40000 23604
rect 0 23520 800 23548
rect 10526 23492 10536 23548
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10800 23492 10810 23548
rect 19850 23492 19860 23548
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 20124 23492 20134 23548
rect 29174 23492 29184 23548
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29448 23492 29458 23548
rect 38498 23492 38508 23548
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38772 23492 38782 23548
rect 39200 23520 40000 23548
rect 17826 23436 17836 23492
rect 17892 23436 17948 23492
rect 18004 23436 18014 23492
rect 2034 23324 2044 23380
rect 2100 23324 10108 23380
rect 10164 23324 10174 23380
rect 11106 23324 11116 23380
rect 11172 23324 15148 23380
rect 19618 23324 19628 23380
rect 19684 23324 25228 23380
rect 25284 23324 25294 23380
rect 27570 23324 27580 23380
rect 27636 23324 30268 23380
rect 30324 23324 30334 23380
rect 15092 23268 15148 23324
rect 5058 23212 5068 23268
rect 5124 23212 12236 23268
rect 12292 23212 12302 23268
rect 15092 23212 15596 23268
rect 15652 23212 17668 23268
rect 18162 23212 18172 23268
rect 18228 23212 19964 23268
rect 20020 23212 20300 23268
rect 20356 23212 20366 23268
rect 23762 23212 23772 23268
rect 23828 23212 30380 23268
rect 30436 23212 30446 23268
rect 30594 23212 30604 23268
rect 30660 23212 36876 23268
rect 36932 23212 36942 23268
rect 17612 23156 17668 23212
rect 13682 23100 13692 23156
rect 13748 23100 14812 23156
rect 14868 23100 14878 23156
rect 16370 23100 16380 23156
rect 16436 23100 17388 23156
rect 17444 23100 17454 23156
rect 17612 23100 18284 23156
rect 18340 23100 19404 23156
rect 19460 23100 19470 23156
rect 24434 23100 24444 23156
rect 24500 23100 28700 23156
rect 28756 23100 29036 23156
rect 29092 23100 29102 23156
rect 14812 23044 14868 23100
rect 14812 22988 18620 23044
rect 18676 22988 19180 23044
rect 19236 22988 19246 23044
rect 0 22932 800 22960
rect 39200 22932 40000 22960
rect 0 22876 1708 22932
rect 1764 22876 1774 22932
rect 18918 22876 18956 22932
rect 19012 22876 19022 22932
rect 38210 22876 38220 22932
rect 38276 22876 40000 22932
rect 0 22848 800 22876
rect 39200 22848 40000 22876
rect 29362 22764 29372 22820
rect 29428 22764 30716 22820
rect 30772 22764 31388 22820
rect 31444 22764 32508 22820
rect 32564 22764 32574 22820
rect 5864 22708 5874 22764
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 6138 22708 6148 22764
rect 15188 22708 15198 22764
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15462 22708 15472 22764
rect 24512 22708 24522 22764
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24786 22708 24796 22764
rect 33836 22708 33846 22764
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 34110 22708 34120 22764
rect 25890 22652 25900 22708
rect 25956 22652 29596 22708
rect 29652 22652 30492 22708
rect 30548 22652 30558 22708
rect 4050 22540 4060 22596
rect 4116 22540 14588 22596
rect 14644 22540 14654 22596
rect 27794 22540 27804 22596
rect 27860 22540 37884 22596
rect 37940 22540 37950 22596
rect 2706 22428 2716 22484
rect 2772 22428 14476 22484
rect 14532 22428 14542 22484
rect 24658 22428 24668 22484
rect 24724 22428 35308 22484
rect 35364 22428 35374 22484
rect 6738 22316 6748 22372
rect 6804 22316 14140 22372
rect 14196 22316 14206 22372
rect 22418 22316 22428 22372
rect 22484 22316 23212 22372
rect 23268 22316 23548 22372
rect 23604 22316 23614 22372
rect 28578 22316 28588 22372
rect 28644 22316 29820 22372
rect 29876 22316 31612 22372
rect 31668 22316 31678 22372
rect 31892 22316 32284 22372
rect 32340 22316 32350 22372
rect 0 22260 800 22288
rect 0 22204 1708 22260
rect 1764 22204 1774 22260
rect 2034 22204 2044 22260
rect 2100 22204 9212 22260
rect 9268 22204 9278 22260
rect 10322 22204 10332 22260
rect 10388 22204 12348 22260
rect 12404 22204 12414 22260
rect 14690 22204 14700 22260
rect 14756 22204 15484 22260
rect 15540 22204 15550 22260
rect 20626 22204 20636 22260
rect 20692 22204 22540 22260
rect 22596 22204 25900 22260
rect 25956 22204 25966 22260
rect 27122 22204 27132 22260
rect 27188 22204 29932 22260
rect 29988 22204 29998 22260
rect 0 22176 800 22204
rect 31892 22148 31948 22316
rect 39200 22260 40000 22288
rect 38210 22204 38220 22260
rect 38276 22204 40000 22260
rect 39200 22176 40000 22204
rect 2146 22092 2156 22148
rect 2212 22092 11228 22148
rect 11284 22092 11294 22148
rect 12114 22092 12124 22148
rect 12180 22092 12572 22148
rect 12628 22092 12638 22148
rect 13458 22092 13468 22148
rect 13524 22092 15820 22148
rect 15876 22092 15886 22148
rect 17266 22092 17276 22148
rect 17332 22092 18732 22148
rect 18788 22092 20076 22148
rect 20132 22092 20412 22148
rect 20468 22092 20478 22148
rect 26852 22092 31388 22148
rect 31444 22092 31948 22148
rect 26852 22036 26908 22092
rect 12450 21980 12460 22036
rect 12516 21980 15260 22036
rect 15316 21980 18060 22036
rect 18116 21980 18126 22036
rect 26562 21980 26572 22036
rect 26628 21980 26908 22036
rect 10526 21924 10536 21980
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10800 21924 10810 21980
rect 19850 21924 19860 21980
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 20124 21924 20134 21980
rect 29174 21924 29184 21980
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29448 21924 29458 21980
rect 38498 21924 38508 21980
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38772 21924 38782 21980
rect 12338 21868 12348 21924
rect 12404 21868 15708 21924
rect 15764 21868 16716 21924
rect 16772 21868 16782 21924
rect 32386 21868 32396 21924
rect 32452 21868 37996 21924
rect 38052 21868 38062 21924
rect 924 21756 2380 21812
rect 2436 21756 2446 21812
rect 2594 21756 2604 21812
rect 2660 21756 13244 21812
rect 13300 21756 13310 21812
rect 17714 21756 17724 21812
rect 17780 21756 25676 21812
rect 25732 21756 26460 21812
rect 26516 21756 27468 21812
rect 27524 21756 27534 21812
rect 28914 21756 28924 21812
rect 28980 21756 37772 21812
rect 37828 21756 37838 21812
rect 0 21588 800 21616
rect 924 21588 980 21756
rect 6850 21644 6860 21700
rect 6916 21644 11004 21700
rect 11060 21644 11070 21700
rect 11676 21644 13748 21700
rect 20290 21644 20300 21700
rect 20356 21644 20366 21700
rect 21298 21644 21308 21700
rect 21364 21644 23324 21700
rect 23380 21644 25508 21700
rect 26002 21644 26012 21700
rect 26068 21644 26348 21700
rect 26404 21644 26684 21700
rect 26740 21644 27804 21700
rect 27860 21644 27870 21700
rect 30146 21644 30156 21700
rect 30212 21644 37884 21700
rect 37940 21644 37950 21700
rect 11676 21588 11732 21644
rect 13692 21588 13748 21644
rect 0 21532 980 21588
rect 2034 21532 2044 21588
rect 2100 21532 11732 21588
rect 12898 21532 12908 21588
rect 12964 21532 13468 21588
rect 13524 21532 13534 21588
rect 13682 21532 13692 21588
rect 13748 21532 13758 21588
rect 15026 21532 15036 21588
rect 15092 21532 17388 21588
rect 17444 21532 17454 21588
rect 0 21504 800 21532
rect 20300 21476 20356 21644
rect 25452 21588 25508 21644
rect 39200 21588 40000 21616
rect 21634 21532 21644 21588
rect 21700 21532 22876 21588
rect 22932 21532 22942 21588
rect 24322 21532 24332 21588
rect 24388 21532 25228 21588
rect 25284 21532 25294 21588
rect 25452 21532 26572 21588
rect 26628 21532 26638 21588
rect 37538 21532 37548 21588
rect 37604 21532 40000 21588
rect 39200 21504 40000 21532
rect 6962 21420 6972 21476
rect 7028 21420 15148 21476
rect 20300 21420 27020 21476
rect 27076 21420 27086 21476
rect 15092 21364 15148 21420
rect 10322 21308 10332 21364
rect 10388 21308 12572 21364
rect 12628 21308 13244 21364
rect 13300 21308 13310 21364
rect 14466 21308 14476 21364
rect 14532 21308 14924 21364
rect 14980 21308 14990 21364
rect 15092 21308 16380 21364
rect 16436 21308 16828 21364
rect 16884 21308 18284 21364
rect 18340 21308 20972 21364
rect 21028 21308 21038 21364
rect 25554 21308 25564 21364
rect 25620 21308 32060 21364
rect 32116 21308 32126 21364
rect 25218 21196 25228 21252
rect 25284 21196 31500 21252
rect 31556 21196 31566 21252
rect 5864 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6148 21196
rect 15188 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15472 21196
rect 24512 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24796 21196
rect 33836 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34120 21196
rect 9314 21084 9324 21140
rect 9380 21084 14924 21140
rect 14980 21084 14990 21140
rect 8372 20972 17388 21028
rect 17444 20972 17454 21028
rect 29922 20972 29932 21028
rect 29988 20972 37212 21028
rect 37268 20972 37278 21028
rect 0 20916 800 20944
rect 0 20860 1708 20916
rect 1764 20860 1774 20916
rect 0 20832 800 20860
rect 8372 20692 8428 20972
rect 39200 20916 40000 20944
rect 10322 20860 10332 20916
rect 10388 20860 12572 20916
rect 12628 20860 14364 20916
rect 14420 20860 17724 20916
rect 17780 20860 17790 20916
rect 30482 20860 30492 20916
rect 30548 20860 31612 20916
rect 31668 20860 32284 20916
rect 32340 20860 32350 20916
rect 38210 20860 38220 20916
rect 38276 20860 40000 20916
rect 39200 20832 40000 20860
rect 14140 20748 15596 20804
rect 15652 20748 15662 20804
rect 29250 20748 29260 20804
rect 29316 20748 30716 20804
rect 30772 20748 30782 20804
rect 30940 20748 37884 20804
rect 37940 20748 37950 20804
rect 14140 20692 14196 20748
rect 30940 20692 30996 20748
rect 1922 20636 1932 20692
rect 1988 20636 8428 20692
rect 13794 20636 13804 20692
rect 13860 20636 14140 20692
rect 14196 20636 14206 20692
rect 14578 20636 14588 20692
rect 14644 20636 15148 20692
rect 15204 20636 15708 20692
rect 15764 20636 16604 20692
rect 16660 20636 16670 20692
rect 17378 20636 17388 20692
rect 17444 20636 18508 20692
rect 18564 20636 18574 20692
rect 21298 20636 21308 20692
rect 21364 20636 22764 20692
rect 22820 20636 22830 20692
rect 26338 20636 26348 20692
rect 26404 20636 27132 20692
rect 27188 20636 27198 20692
rect 28018 20636 28028 20692
rect 28084 20636 30996 20692
rect 31714 20636 31724 20692
rect 31780 20636 32956 20692
rect 33012 20636 33022 20692
rect 33282 20636 33292 20692
rect 33348 20636 36092 20692
rect 36148 20636 36158 20692
rect 8372 20524 14252 20580
rect 14308 20524 14318 20580
rect 15092 20524 15372 20580
rect 15428 20524 17276 20580
rect 17332 20524 17342 20580
rect 21634 20524 21644 20580
rect 21700 20524 23548 20580
rect 23604 20524 27468 20580
rect 27524 20524 31164 20580
rect 31220 20524 31836 20580
rect 31892 20524 31902 20580
rect 8372 20356 8428 20524
rect 15092 20468 15148 20524
rect 13234 20412 13244 20468
rect 13300 20412 15148 20468
rect 16258 20412 16268 20468
rect 16324 20412 16828 20468
rect 16884 20412 16894 20468
rect 10526 20356 10536 20412
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10800 20356 10810 20412
rect 19850 20356 19860 20412
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 20124 20356 20134 20412
rect 29174 20356 29184 20412
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29448 20356 29458 20412
rect 38498 20356 38508 20412
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38772 20356 38782 20412
rect 2034 20300 2044 20356
rect 2100 20300 8428 20356
rect 13682 20300 13692 20356
rect 13748 20300 14924 20356
rect 14980 20300 14990 20356
rect 0 20244 800 20272
rect 39200 20244 40000 20272
rect 0 20188 1708 20244
rect 1764 20188 1774 20244
rect 17602 20188 17612 20244
rect 17668 20188 18508 20244
rect 18564 20188 19852 20244
rect 19908 20188 21308 20244
rect 21364 20188 21374 20244
rect 22764 20188 23212 20244
rect 23268 20188 23884 20244
rect 23940 20188 23950 20244
rect 38434 20188 38444 20244
rect 38500 20188 40000 20244
rect 0 20160 800 20188
rect 22764 20132 22820 20188
rect 39200 20160 40000 20188
rect 2034 20076 2044 20132
rect 2100 20076 15148 20132
rect 16930 20076 16940 20132
rect 16996 20076 17500 20132
rect 17556 20076 17566 20132
rect 17826 20076 17836 20132
rect 17892 20076 19068 20132
rect 19124 20076 19134 20132
rect 21186 20076 21196 20132
rect 21252 20076 22820 20132
rect 22978 20076 22988 20132
rect 23044 20076 23772 20132
rect 23828 20076 23838 20132
rect 25554 20076 25564 20132
rect 25620 20076 26908 20132
rect 28578 20076 28588 20132
rect 28644 20076 36540 20132
rect 36596 20076 36606 20132
rect 15092 20020 15148 20076
rect 12002 19964 12012 20020
rect 12068 19964 12684 20020
rect 12740 19964 13244 20020
rect 13300 19964 13310 20020
rect 15092 19964 16380 20020
rect 16436 19964 16828 20020
rect 16884 19964 17948 20020
rect 18004 19964 18732 20020
rect 18788 19964 21644 20020
rect 21700 19964 21710 20020
rect 22306 19964 22316 20020
rect 22372 19964 24108 20020
rect 24164 19964 24174 20020
rect 26852 19908 26908 20076
rect 27010 19964 27020 20020
rect 27076 19964 29036 20020
rect 29092 19964 29102 20020
rect 31892 19964 37884 20020
rect 37940 19964 37950 20020
rect 31892 19908 31948 19964
rect 19282 19852 19292 19908
rect 19348 19852 20524 19908
rect 20580 19852 21980 19908
rect 22036 19852 22046 19908
rect 26852 19852 31948 19908
rect 2930 19740 2940 19796
rect 2996 19740 12572 19796
rect 12628 19740 12638 19796
rect 22530 19740 22540 19796
rect 22596 19740 23548 19796
rect 23604 19740 27020 19796
rect 27076 19740 27086 19796
rect 0 19572 800 19600
rect 5864 19572 5874 19628
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 6138 19572 6148 19628
rect 15188 19572 15198 19628
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15462 19572 15472 19628
rect 24512 19572 24522 19628
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24786 19572 24796 19628
rect 33836 19572 33846 19628
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 34110 19572 34120 19628
rect 39200 19572 40000 19600
rect 0 19516 1708 19572
rect 1764 19516 2492 19572
rect 2548 19516 2558 19572
rect 9650 19516 9660 19572
rect 9716 19516 11228 19572
rect 11284 19516 14700 19572
rect 14756 19516 14766 19572
rect 38210 19516 38220 19572
rect 38276 19516 40000 19572
rect 0 19488 800 19516
rect 39200 19488 40000 19516
rect 14466 19404 14476 19460
rect 14532 19404 15596 19460
rect 15652 19404 15662 19460
rect 22642 19404 22652 19460
rect 22708 19404 32956 19460
rect 33012 19404 33022 19460
rect 15596 19348 15652 19404
rect 10546 19292 10556 19348
rect 10612 19292 11452 19348
rect 11508 19292 11518 19348
rect 15596 19292 25900 19348
rect 25956 19292 26124 19348
rect 26180 19292 26572 19348
rect 26628 19292 26638 19348
rect 18162 19180 18172 19236
rect 18228 19180 18844 19236
rect 18900 19180 18910 19236
rect 23986 19180 23996 19236
rect 24052 19180 27580 19236
rect 27636 19180 29596 19236
rect 29652 19180 29662 19236
rect 15922 19068 15932 19124
rect 15988 19068 16604 19124
rect 16660 19068 16670 19124
rect 17826 19068 17836 19124
rect 17892 19068 19180 19124
rect 19236 19068 20524 19124
rect 20580 19068 20590 19124
rect 28130 19068 28140 19124
rect 28196 19068 29148 19124
rect 29204 19068 29214 19124
rect 30146 19068 30156 19124
rect 30212 19068 30940 19124
rect 30996 19068 31006 19124
rect 31892 19068 37884 19124
rect 37940 19068 37950 19124
rect 31892 19012 31948 19068
rect 2034 18956 2044 19012
rect 2100 18956 14364 19012
rect 14420 18956 15372 19012
rect 15428 18956 15438 19012
rect 20066 18956 20076 19012
rect 20132 18956 20748 19012
rect 20804 18956 20814 19012
rect 29474 18956 29484 19012
rect 29540 18956 30772 19012
rect 31266 18956 31276 19012
rect 31332 18956 31948 19012
rect 38210 18956 38220 19012
rect 38276 18956 38948 19012
rect 0 18900 800 18928
rect 0 18844 1708 18900
rect 1764 18844 2492 18900
rect 2548 18844 2558 18900
rect 0 18816 800 18844
rect 10526 18788 10536 18844
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10800 18788 10810 18844
rect 19850 18788 19860 18844
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 20124 18788 20134 18844
rect 29174 18788 29184 18844
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29448 18788 29458 18844
rect 13458 18732 13468 18788
rect 13524 18732 14252 18788
rect 14308 18732 14318 18788
rect 30716 18676 30772 18956
rect 38892 18900 38948 18956
rect 39200 18900 40000 18928
rect 38892 18844 40000 18900
rect 38498 18788 38508 18844
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38772 18788 38782 18844
rect 39200 18816 40000 18844
rect 14690 18620 14700 18676
rect 14756 18620 20188 18676
rect 20244 18620 20860 18676
rect 20916 18620 20926 18676
rect 30716 18620 36092 18676
rect 36148 18620 36158 18676
rect 16594 18508 16604 18564
rect 16660 18508 17276 18564
rect 17332 18508 19964 18564
rect 20020 18508 20030 18564
rect 2034 18396 2044 18452
rect 2100 18396 8428 18452
rect 13010 18396 13020 18452
rect 13076 18396 13692 18452
rect 13748 18396 13758 18452
rect 18386 18396 18396 18452
rect 18452 18396 18956 18452
rect 19012 18396 19022 18452
rect 19394 18396 19404 18452
rect 19460 18396 24108 18452
rect 24164 18396 25228 18452
rect 25284 18396 25294 18452
rect 29586 18396 29596 18452
rect 29652 18396 31052 18452
rect 31108 18396 31118 18452
rect 32386 18396 32396 18452
rect 32452 18396 37884 18452
rect 37940 18396 37950 18452
rect 8372 18340 8428 18396
rect 8372 18284 13356 18340
rect 13412 18284 13422 18340
rect 14242 18284 14252 18340
rect 14308 18284 15148 18340
rect 15362 18284 15372 18340
rect 15428 18284 18844 18340
rect 18900 18284 19516 18340
rect 19572 18284 21084 18340
rect 21140 18284 23324 18340
rect 23380 18284 23390 18340
rect 24322 18284 24332 18340
rect 24388 18284 27468 18340
rect 27524 18284 31388 18340
rect 31444 18284 31454 18340
rect 0 18228 800 18256
rect 15092 18228 15148 18284
rect 39200 18228 40000 18256
rect 0 18172 1708 18228
rect 1764 18172 1774 18228
rect 8754 18172 8764 18228
rect 8820 18172 10556 18228
rect 10612 18172 10622 18228
rect 15092 18172 16156 18228
rect 16212 18172 16222 18228
rect 29810 18172 29820 18228
rect 29876 18172 31612 18228
rect 31668 18172 31678 18228
rect 31892 18172 34916 18228
rect 38210 18172 38220 18228
rect 38276 18172 40000 18228
rect 0 18144 800 18172
rect 10070 18060 10108 18116
rect 10164 18060 10174 18116
rect 10322 18060 10332 18116
rect 10388 18060 10892 18116
rect 10948 18060 10958 18116
rect 5864 18004 5874 18060
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 6138 18004 6148 18060
rect 15188 18004 15198 18060
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15462 18004 15472 18060
rect 24512 18004 24522 18060
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24786 18004 24796 18060
rect 31892 18004 31948 18172
rect 34860 18116 34916 18172
rect 39200 18144 40000 18172
rect 34850 18060 34860 18116
rect 34916 18060 34926 18116
rect 33836 18004 33846 18060
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 34110 18004 34120 18060
rect 12114 17948 12124 18004
rect 12180 17948 12908 18004
rect 12964 17948 12974 18004
rect 25218 17948 25228 18004
rect 25284 17948 31948 18004
rect 34188 17948 36316 18004
rect 36372 17948 36382 18004
rect 10434 17836 10444 17892
rect 10500 17836 12684 17892
rect 12740 17836 12750 17892
rect 14802 17836 14812 17892
rect 14868 17836 15484 17892
rect 15540 17836 15550 17892
rect 24220 17836 26348 17892
rect 26404 17836 26414 17892
rect 2706 17724 2716 17780
rect 2772 17724 8708 17780
rect 0 17556 800 17584
rect 0 17500 1708 17556
rect 1764 17500 1774 17556
rect 2034 17500 2044 17556
rect 2100 17500 8428 17556
rect 8484 17500 8494 17556
rect 0 17472 800 17500
rect 8652 17444 8708 17724
rect 12684 17668 12740 17836
rect 24220 17780 24276 17836
rect 34188 17780 34244 17948
rect 15092 17668 15148 17780
rect 15204 17724 15214 17780
rect 16146 17724 16156 17780
rect 16212 17724 18284 17780
rect 18340 17724 19404 17780
rect 19460 17724 19470 17780
rect 23538 17724 23548 17780
rect 23604 17724 24220 17780
rect 24276 17724 24286 17780
rect 25778 17724 25788 17780
rect 25844 17724 34244 17780
rect 12684 17612 14812 17668
rect 14868 17612 15148 17668
rect 21746 17612 21756 17668
rect 21812 17612 22764 17668
rect 22820 17612 22988 17668
rect 23044 17612 23054 17668
rect 24882 17612 24892 17668
rect 24948 17612 25564 17668
rect 25620 17612 25630 17668
rect 28578 17612 28588 17668
rect 28644 17612 37212 17668
rect 37268 17612 37278 17668
rect 39200 17556 40000 17584
rect 10658 17500 10668 17556
rect 10724 17500 10892 17556
rect 10948 17500 10958 17556
rect 11666 17500 11676 17556
rect 11732 17500 12572 17556
rect 12628 17500 15708 17556
rect 15764 17500 15774 17556
rect 17014 17500 17052 17556
rect 17108 17500 17118 17556
rect 23762 17500 23772 17556
rect 23828 17500 26124 17556
rect 26180 17500 26908 17556
rect 38210 17500 38220 17556
rect 38276 17500 40000 17556
rect 26852 17444 26908 17500
rect 39200 17472 40000 17500
rect 8652 17388 15596 17444
rect 15652 17388 15662 17444
rect 18386 17388 18396 17444
rect 18452 17388 18462 17444
rect 23314 17388 23324 17444
rect 23380 17388 24668 17444
rect 24724 17388 25116 17444
rect 25172 17388 25900 17444
rect 25956 17388 25966 17444
rect 26852 17388 27132 17444
rect 27188 17388 31276 17444
rect 31332 17388 31342 17444
rect 10526 17220 10536 17276
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10800 17220 10810 17276
rect 18396 17220 18452 17388
rect 19850 17220 19860 17276
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 20124 17220 20134 17276
rect 29174 17220 29184 17276
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29448 17220 29458 17276
rect 38498 17220 38508 17276
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38772 17220 38782 17276
rect 18162 17164 18172 17220
rect 18228 17164 18452 17220
rect 25778 17164 25788 17220
rect 25844 17164 28364 17220
rect 28420 17164 28924 17220
rect 28980 17164 28990 17220
rect 10770 17052 10780 17108
rect 10836 17052 11228 17108
rect 11284 17052 11294 17108
rect 14578 17052 14588 17108
rect 14644 17052 17388 17108
rect 17444 17052 17454 17108
rect 17602 17052 17612 17108
rect 17668 17052 23660 17108
rect 23716 17052 23726 17108
rect 25666 17052 25676 17108
rect 25732 17052 37884 17108
rect 37940 17052 37950 17108
rect 17612 16996 17668 17052
rect 2034 16940 2044 16996
rect 2100 16940 15148 16996
rect 15204 16940 15214 16996
rect 16482 16940 16492 16996
rect 16548 16940 17668 16996
rect 18946 16940 18956 16996
rect 19012 16940 19964 16996
rect 20020 16940 21532 16996
rect 21588 16940 21980 16996
rect 22036 16940 22046 16996
rect 26562 16940 26572 16996
rect 26628 16940 27244 16996
rect 27300 16940 27310 16996
rect 0 16884 800 16912
rect 39200 16884 40000 16912
rect 0 16828 2380 16884
rect 2436 16828 2446 16884
rect 2604 16828 12852 16884
rect 13010 16828 13020 16884
rect 13076 16828 13580 16884
rect 13636 16828 13646 16884
rect 13804 16828 14868 16884
rect 15026 16828 15036 16884
rect 15092 16828 15932 16884
rect 15988 16828 15998 16884
rect 21858 16828 21868 16884
rect 21924 16828 22876 16884
rect 22932 16828 22942 16884
rect 23874 16828 23884 16884
rect 23940 16828 24892 16884
rect 24948 16828 27132 16884
rect 27188 16828 29484 16884
rect 29540 16828 29550 16884
rect 37538 16828 37548 16884
rect 37604 16828 40000 16884
rect 0 16800 800 16828
rect 2604 16772 2660 16828
rect 12796 16772 12852 16828
rect 13804 16772 13860 16828
rect 2146 16716 2156 16772
rect 2212 16716 2660 16772
rect 10434 16716 10444 16772
rect 10500 16716 11676 16772
rect 11732 16716 11742 16772
rect 12796 16716 13860 16772
rect 14812 16772 14868 16828
rect 39200 16800 40000 16828
rect 14812 16716 15148 16772
rect 15204 16716 15214 16772
rect 20626 16716 20636 16772
rect 20692 16716 22652 16772
rect 22708 16716 22718 16772
rect 29138 16716 29148 16772
rect 29204 16716 29708 16772
rect 29764 16716 30828 16772
rect 30884 16716 31500 16772
rect 31556 16716 31566 16772
rect 2034 16604 2044 16660
rect 2100 16604 11116 16660
rect 11172 16604 11182 16660
rect 14812 16604 16380 16660
rect 16436 16604 16446 16660
rect 17266 16604 17276 16660
rect 17332 16604 17724 16660
rect 17780 16604 17790 16660
rect 14812 16548 14868 16604
rect 10098 16492 10108 16548
rect 10164 16492 12684 16548
rect 12740 16492 14812 16548
rect 14868 16492 14878 16548
rect 17602 16492 17612 16548
rect 17668 16492 17678 16548
rect 5864 16436 5874 16492
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 6138 16436 6148 16492
rect 15188 16436 15198 16492
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15462 16436 15472 16492
rect 17612 16436 17668 16492
rect 24512 16436 24522 16492
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24786 16436 24796 16492
rect 33836 16436 33846 16492
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 34110 16436 34120 16492
rect 10658 16380 10668 16436
rect 10724 16380 10892 16436
rect 10948 16380 10958 16436
rect 17014 16380 17052 16436
rect 17108 16380 17118 16436
rect 17378 16380 17388 16436
rect 17444 16380 17668 16436
rect 8866 16268 8876 16324
rect 8932 16268 19516 16324
rect 19572 16268 19582 16324
rect 0 16212 800 16240
rect 39200 16212 40000 16240
rect 0 16156 1708 16212
rect 1764 16156 1774 16212
rect 9762 16156 9772 16212
rect 9828 16156 10332 16212
rect 10388 16156 10398 16212
rect 10546 16156 10556 16212
rect 10612 16156 12572 16212
rect 12628 16156 15484 16212
rect 15540 16156 15550 16212
rect 16604 16156 18620 16212
rect 18676 16156 18686 16212
rect 23202 16156 23212 16212
rect 23268 16156 23278 16212
rect 30818 16156 30828 16212
rect 30884 16156 37884 16212
rect 37940 16156 37950 16212
rect 38210 16156 38220 16212
rect 38276 16156 40000 16212
rect 0 16128 800 16156
rect 16604 16100 16660 16156
rect 23212 16100 23268 16156
rect 39200 16128 40000 16156
rect 12786 16044 12796 16100
rect 12852 16044 14140 16100
rect 14196 16044 14206 16100
rect 14364 16044 16660 16100
rect 16716 16044 20636 16100
rect 20692 16044 20702 16100
rect 23212 16044 23772 16100
rect 23828 16044 25004 16100
rect 25060 16044 25070 16100
rect 14364 15988 14420 16044
rect 16716 15988 16772 16044
rect 9090 15932 9100 15988
rect 9156 15932 10108 15988
rect 10164 15932 10174 15988
rect 11442 15932 11452 15988
rect 11508 15932 12012 15988
rect 12068 15932 12078 15988
rect 12338 15932 12348 15988
rect 12404 15932 13468 15988
rect 13524 15932 13534 15988
rect 13794 15932 13804 15988
rect 13860 15932 14028 15988
rect 14084 15932 14420 15988
rect 15092 15932 16772 15988
rect 16930 15932 16940 15988
rect 16996 15932 17836 15988
rect 17892 15932 17902 15988
rect 24546 15932 24556 15988
rect 24612 15932 37884 15988
rect 37940 15932 37950 15988
rect 13804 15876 13860 15932
rect 1698 15820 1708 15876
rect 1764 15820 1774 15876
rect 2258 15820 2268 15876
rect 2324 15820 10444 15876
rect 10500 15820 10510 15876
rect 12450 15820 12460 15876
rect 12516 15820 13860 15876
rect 1708 15652 1764 15820
rect 15092 15764 15148 15932
rect 16258 15820 16268 15876
rect 16324 15820 18172 15876
rect 18228 15820 18238 15876
rect 21410 15820 21420 15876
rect 21476 15820 21980 15876
rect 22036 15820 22046 15876
rect 28354 15820 28364 15876
rect 28420 15820 33516 15876
rect 33572 15820 33582 15876
rect 11330 15708 11340 15764
rect 11396 15708 11676 15764
rect 11732 15708 15148 15764
rect 15810 15708 15820 15764
rect 15876 15708 16492 15764
rect 16548 15708 16716 15764
rect 16772 15708 16782 15764
rect 10526 15652 10536 15708
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10800 15652 10810 15708
rect 19850 15652 19860 15708
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 20124 15652 20134 15708
rect 29174 15652 29184 15708
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29448 15652 29458 15708
rect 38498 15652 38508 15708
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38772 15652 38782 15708
rect 924 15596 1764 15652
rect 20514 15596 20524 15652
rect 20580 15596 25564 15652
rect 25620 15596 26236 15652
rect 26292 15596 26302 15652
rect 0 15540 800 15568
rect 924 15540 980 15596
rect 39200 15540 40000 15568
rect 0 15484 980 15540
rect 8194 15484 8204 15540
rect 8260 15484 14476 15540
rect 14532 15484 15596 15540
rect 15652 15484 16828 15540
rect 16884 15484 17948 15540
rect 18004 15484 23660 15540
rect 23716 15484 23726 15540
rect 28802 15484 28812 15540
rect 28868 15484 31948 15540
rect 38434 15484 38444 15540
rect 38500 15484 40000 15540
rect 0 15456 800 15484
rect 31892 15428 31948 15484
rect 39200 15456 40000 15484
rect 9538 15372 9548 15428
rect 9604 15372 9996 15428
rect 10052 15372 11340 15428
rect 11396 15372 11406 15428
rect 17602 15372 17612 15428
rect 17668 15372 22316 15428
rect 22372 15372 22382 15428
rect 25890 15372 25900 15428
rect 25956 15372 26572 15428
rect 26628 15372 26638 15428
rect 31892 15372 37884 15428
rect 37940 15372 37950 15428
rect 6290 15260 6300 15316
rect 6356 15260 16044 15316
rect 16100 15260 16110 15316
rect 18386 15260 18396 15316
rect 18452 15260 18844 15316
rect 18900 15260 18910 15316
rect 19170 15260 19180 15316
rect 19236 15260 21196 15316
rect 21252 15260 21262 15316
rect 21634 15260 21644 15316
rect 21700 15260 25676 15316
rect 25732 15260 25742 15316
rect 15586 15148 15596 15204
rect 15652 15148 18956 15204
rect 19012 15148 19022 15204
rect 20178 15148 20188 15204
rect 20244 15148 20972 15204
rect 21028 15148 21756 15204
rect 21812 15148 21822 15204
rect 22978 15148 22988 15204
rect 23044 15148 24892 15204
rect 24948 15148 27580 15204
rect 27636 15148 29148 15204
rect 29204 15148 29214 15204
rect 0 14868 800 14896
rect 5864 14868 5874 14924
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 6138 14868 6148 14924
rect 15188 14868 15198 14924
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15462 14868 15472 14924
rect 24512 14868 24522 14924
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24786 14868 24796 14924
rect 33836 14868 33846 14924
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 34110 14868 34120 14924
rect 39200 14868 40000 14896
rect 0 14812 1708 14868
rect 1764 14812 1774 14868
rect 10322 14812 10332 14868
rect 10388 14812 10444 14868
rect 10500 14812 10510 14868
rect 38210 14812 38220 14868
rect 38276 14812 40000 14868
rect 0 14784 800 14812
rect 39200 14784 40000 14812
rect 7634 14700 7644 14756
rect 7700 14700 18844 14756
rect 18900 14700 18910 14756
rect 6402 14588 6412 14644
rect 6468 14588 15596 14644
rect 15652 14588 15662 14644
rect 17266 14588 17276 14644
rect 17332 14588 17836 14644
rect 17892 14588 17902 14644
rect 9202 14476 9212 14532
rect 9268 14476 10220 14532
rect 10276 14476 10286 14532
rect 10658 14476 10668 14532
rect 10724 14476 13916 14532
rect 13972 14476 14924 14532
rect 14980 14476 15596 14532
rect 15652 14476 15662 14532
rect 17938 14476 17948 14532
rect 18004 14476 18508 14532
rect 18564 14476 20188 14532
rect 20244 14476 21308 14532
rect 21364 14476 21374 14532
rect 22194 14476 22204 14532
rect 22260 14476 22988 14532
rect 23044 14476 23436 14532
rect 23492 14476 23502 14532
rect 26562 14476 26572 14532
rect 26628 14476 27356 14532
rect 27412 14476 27422 14532
rect 28018 14476 28028 14532
rect 28084 14476 28588 14532
rect 28644 14476 29372 14532
rect 29428 14476 29438 14532
rect 9874 14364 9884 14420
rect 9940 14364 10332 14420
rect 10388 14364 10398 14420
rect 11890 14364 11900 14420
rect 11956 14364 12908 14420
rect 12964 14364 13692 14420
rect 13748 14364 13758 14420
rect 14578 14364 14588 14420
rect 14644 14364 17724 14420
rect 17780 14364 17790 14420
rect 18050 14364 18060 14420
rect 18116 14364 19628 14420
rect 19684 14364 20524 14420
rect 20580 14364 20590 14420
rect 21970 14364 21980 14420
rect 22036 14364 22316 14420
rect 22372 14364 23212 14420
rect 23268 14364 23278 14420
rect 24770 14364 24780 14420
rect 24836 14364 25452 14420
rect 25508 14364 25518 14420
rect 28130 14364 28140 14420
rect 28196 14364 37884 14420
rect 37940 14364 37950 14420
rect 1698 14252 1708 14308
rect 1764 14252 1774 14308
rect 3332 14252 12572 14308
rect 12628 14252 12638 14308
rect 12786 14252 12796 14308
rect 12852 14252 13580 14308
rect 13636 14252 13646 14308
rect 14242 14252 14252 14308
rect 14308 14252 15708 14308
rect 15764 14252 17500 14308
rect 17556 14252 17566 14308
rect 19170 14252 19180 14308
rect 19236 14252 19684 14308
rect 20962 14252 20972 14308
rect 21028 14252 21868 14308
rect 21924 14252 21934 14308
rect 38210 14252 38220 14308
rect 38276 14252 38948 14308
rect 0 14196 800 14224
rect 1708 14196 1764 14252
rect 0 14140 1764 14196
rect 0 14112 800 14140
rect 3332 14084 3388 14252
rect 19628 14196 19684 14252
rect 38892 14196 38948 14252
rect 39200 14196 40000 14224
rect 12450 14140 12460 14196
rect 12516 14140 13244 14196
rect 13300 14140 16044 14196
rect 16100 14140 17164 14196
rect 17220 14140 17230 14196
rect 19618 14140 19628 14196
rect 19684 14140 19694 14196
rect 38892 14140 40000 14196
rect 10526 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10810 14140
rect 19850 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20134 14140
rect 29174 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29458 14140
rect 38498 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38782 14140
rect 39200 14112 40000 14140
rect 2034 14028 2044 14084
rect 2100 14028 3388 14084
rect 16930 14028 16940 14084
rect 16996 14028 17276 14084
rect 17332 14028 17500 14084
rect 17556 14028 17566 14084
rect 26852 14028 28252 14084
rect 28308 14028 28812 14084
rect 28868 14028 28878 14084
rect 26852 13972 26908 14028
rect 10322 13916 10332 13972
rect 10388 13916 10556 13972
rect 10612 13916 10622 13972
rect 12786 13916 12796 13972
rect 12852 13916 13468 13972
rect 13524 13916 13534 13972
rect 16370 13916 16380 13972
rect 16436 13916 17052 13972
rect 17108 13916 19516 13972
rect 19572 13916 19582 13972
rect 22306 13916 22316 13972
rect 22372 13916 26908 13972
rect 27234 13916 27244 13972
rect 27300 13916 37660 13972
rect 37716 13916 37726 13972
rect 2034 13804 2044 13860
rect 2100 13804 11452 13860
rect 11508 13804 11518 13860
rect 25554 13804 25564 13860
rect 25620 13804 25630 13860
rect 6738 13692 6748 13748
rect 6804 13692 16156 13748
rect 16212 13692 17724 13748
rect 17780 13692 17790 13748
rect 25564 13636 25620 13804
rect 26562 13692 26572 13748
rect 26628 13692 27580 13748
rect 27636 13692 27646 13748
rect 9986 13580 9996 13636
rect 10052 13580 14364 13636
rect 14420 13580 15708 13636
rect 15764 13580 17500 13636
rect 17556 13580 17566 13636
rect 25564 13580 30044 13636
rect 30100 13580 30110 13636
rect 32498 13580 32508 13636
rect 32564 13580 38108 13636
rect 38164 13580 38174 13636
rect 0 13524 800 13552
rect 39200 13524 40000 13552
rect 0 13468 1708 13524
rect 1764 13468 1774 13524
rect 11106 13468 11116 13524
rect 11172 13468 11676 13524
rect 11732 13468 11742 13524
rect 15036 13468 15652 13524
rect 23090 13468 23100 13524
rect 23156 13468 25228 13524
rect 25284 13468 26684 13524
rect 26740 13468 26750 13524
rect 29026 13468 29036 13524
rect 29092 13468 37884 13524
rect 37940 13468 37950 13524
rect 38210 13468 38220 13524
rect 38276 13468 40000 13524
rect 0 13440 800 13468
rect 10770 13356 10780 13412
rect 10836 13356 13132 13412
rect 13188 13356 13198 13412
rect 5864 13300 5874 13356
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 6138 13300 6148 13356
rect 15036 13300 15092 13468
rect 15596 13412 15652 13468
rect 39200 13440 40000 13468
rect 15596 13356 15932 13412
rect 15988 13356 15998 13412
rect 26002 13356 26012 13412
rect 26068 13356 26628 13412
rect 15188 13300 15198 13356
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15462 13300 15472 13356
rect 24512 13300 24522 13356
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24786 13300 24796 13356
rect 26572 13300 26628 13356
rect 33836 13300 33846 13356
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 34110 13300 34120 13356
rect 9212 13244 15092 13300
rect 26562 13244 26572 13300
rect 26628 13244 26638 13300
rect 9212 13188 9268 13244
rect 2706 13132 2716 13188
rect 2772 13132 9268 13188
rect 13346 13132 13356 13188
rect 13412 13132 14028 13188
rect 14084 13132 14094 13188
rect 14802 13132 14812 13188
rect 14868 13132 15260 13188
rect 15316 13132 16156 13188
rect 16212 13132 16222 13188
rect 13916 13020 15596 13076
rect 15652 13020 16044 13076
rect 16100 13020 16110 13076
rect 20412 13020 21420 13076
rect 21476 13020 21486 13076
rect 30370 13020 30380 13076
rect 30436 13020 37996 13076
rect 38052 13020 38062 13076
rect 13916 12964 13972 13020
rect 20412 12964 20468 13020
rect 2034 12908 2044 12964
rect 2100 12908 9548 12964
rect 9604 12908 9614 12964
rect 10546 12908 10556 12964
rect 10612 12908 13916 12964
rect 13972 12908 13982 12964
rect 14914 12908 14924 12964
rect 14980 12908 15372 12964
rect 15428 12908 15820 12964
rect 15876 12908 15886 12964
rect 16482 12908 16492 12964
rect 16548 12908 17052 12964
rect 17108 12908 17118 12964
rect 17714 12908 17724 12964
rect 17780 12908 20412 12964
rect 20468 12908 20478 12964
rect 20738 12908 20748 12964
rect 20804 12908 22092 12964
rect 22148 12908 24556 12964
rect 24612 12908 27692 12964
rect 27748 12908 27758 12964
rect 31892 12908 37772 12964
rect 37828 12908 37838 12964
rect 0 12852 800 12880
rect 0 12796 1708 12852
rect 1764 12796 1774 12852
rect 13122 12796 13132 12852
rect 13188 12796 15148 12852
rect 15204 12796 16268 12852
rect 16324 12796 16334 12852
rect 16818 12796 16828 12852
rect 16884 12796 17500 12852
rect 17556 12796 17948 12852
rect 18004 12796 18014 12852
rect 25778 12796 25788 12852
rect 25844 12796 28140 12852
rect 28196 12796 28206 12852
rect 0 12768 800 12796
rect 31892 12740 31948 12908
rect 39200 12852 40000 12880
rect 38210 12796 38220 12852
rect 38276 12796 40000 12852
rect 39200 12768 40000 12796
rect 12786 12684 12796 12740
rect 12852 12684 13580 12740
rect 13636 12684 13646 12740
rect 17042 12684 17052 12740
rect 17108 12684 19740 12740
rect 19796 12684 19806 12740
rect 20178 12684 20188 12740
rect 20244 12684 20972 12740
rect 21028 12684 21038 12740
rect 27794 12684 27804 12740
rect 27860 12684 31948 12740
rect 32610 12684 32620 12740
rect 32676 12684 34524 12740
rect 34580 12684 34590 12740
rect 10526 12516 10536 12572
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10800 12516 10810 12572
rect 19850 12516 19860 12572
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 20124 12516 20134 12572
rect 29174 12516 29184 12572
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29448 12516 29458 12572
rect 38498 12516 38508 12572
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38772 12516 38782 12572
rect 12012 12460 14252 12516
rect 14308 12460 14318 12516
rect 12012 12404 12068 12460
rect 9874 12348 9884 12404
rect 9940 12348 12068 12404
rect 12226 12348 12236 12404
rect 12292 12348 13356 12404
rect 13412 12348 13422 12404
rect 17490 12348 17500 12404
rect 17556 12348 17724 12404
rect 17780 12348 17790 12404
rect 25778 12348 25788 12404
rect 25844 12348 26796 12404
rect 26852 12348 26862 12404
rect 10546 12236 10556 12292
rect 10612 12236 11340 12292
rect 11396 12236 11406 12292
rect 11666 12236 11676 12292
rect 11732 12236 13804 12292
rect 13860 12236 13870 12292
rect 29026 12236 29036 12292
rect 29092 12236 37212 12292
rect 37268 12236 37278 12292
rect 0 12180 800 12208
rect 39200 12180 40000 12208
rect 0 12124 2380 12180
rect 2436 12124 2446 12180
rect 13458 12124 13468 12180
rect 13524 12124 14028 12180
rect 14084 12124 14094 12180
rect 20066 12124 20076 12180
rect 20132 12124 23100 12180
rect 23156 12124 23166 12180
rect 24994 12124 25004 12180
rect 25060 12124 25452 12180
rect 25508 12124 26236 12180
rect 26292 12124 26302 12180
rect 37538 12124 37548 12180
rect 37604 12124 40000 12180
rect 0 12096 800 12124
rect 39200 12096 40000 12124
rect 10546 12012 10556 12068
rect 10612 12012 12012 12068
rect 12068 12012 15260 12068
rect 15316 12012 15820 12068
rect 15876 12012 15886 12068
rect 11666 11900 11676 11956
rect 11732 11900 12684 11956
rect 12740 11900 12750 11956
rect 13794 11900 13804 11956
rect 13860 11900 15708 11956
rect 15764 11900 15774 11956
rect 24322 11900 24332 11956
rect 24388 11900 25900 11956
rect 25956 11900 25966 11956
rect 11004 11788 12572 11844
rect 12628 11788 12638 11844
rect 5864 11732 5874 11788
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 6138 11732 6148 11788
rect 11004 11732 11060 11788
rect 15188 11732 15198 11788
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15462 11732 15472 11788
rect 24512 11732 24522 11788
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24786 11732 24796 11788
rect 33836 11732 33846 11788
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 34110 11732 34120 11788
rect 10994 11676 11004 11732
rect 11060 11676 11070 11732
rect 12450 11676 12460 11732
rect 12516 11676 12526 11732
rect 23202 11676 23212 11732
rect 23268 11676 24220 11732
rect 24276 11676 24286 11732
rect 25218 11676 25228 11732
rect 25284 11676 27580 11732
rect 27636 11676 27646 11732
rect 12460 11620 12516 11676
rect 3332 11564 12516 11620
rect 19394 11564 19404 11620
rect 19460 11564 23324 11620
rect 23380 11564 26124 11620
rect 26180 11564 26684 11620
rect 26740 11564 26750 11620
rect 27010 11564 27020 11620
rect 27076 11564 27804 11620
rect 27860 11564 27870 11620
rect 0 11508 800 11536
rect 3332 11508 3388 11564
rect 39200 11508 40000 11536
rect 0 11452 1708 11508
rect 1764 11452 1774 11508
rect 2034 11452 2044 11508
rect 2100 11452 3388 11508
rect 10322 11452 10332 11508
rect 10388 11452 14924 11508
rect 14980 11452 14990 11508
rect 16034 11452 16044 11508
rect 16100 11452 17276 11508
rect 17332 11452 17342 11508
rect 24210 11452 24220 11508
rect 24276 11452 26236 11508
rect 26292 11452 26302 11508
rect 38210 11452 38220 11508
rect 38276 11452 40000 11508
rect 0 11424 800 11452
rect 39200 11424 40000 11452
rect 12338 11340 12348 11396
rect 12404 11340 13692 11396
rect 13748 11340 13758 11396
rect 16706 11340 16716 11396
rect 16772 11340 17724 11396
rect 17780 11340 17790 11396
rect 20402 11340 20412 11396
rect 20468 11340 22092 11396
rect 22148 11340 22158 11396
rect 24882 11340 24892 11396
rect 24948 11340 25564 11396
rect 25620 11340 25630 11396
rect 16370 11228 16380 11284
rect 16436 11228 17612 11284
rect 17668 11228 17678 11284
rect 18386 11228 18396 11284
rect 18452 11228 21420 11284
rect 21476 11228 21486 11284
rect 21746 11228 21756 11284
rect 21812 11228 24556 11284
rect 24612 11228 24622 11284
rect 28130 11228 28140 11284
rect 28196 11228 29148 11284
rect 29204 11228 29214 11284
rect 1698 11116 1708 11172
rect 1764 11116 1774 11172
rect 8754 11116 8764 11172
rect 8820 11116 15036 11172
rect 15092 11116 15484 11172
rect 15540 11116 15550 11172
rect 16930 11116 16940 11172
rect 16996 11116 18956 11172
rect 19012 11116 19022 11172
rect 27234 11116 27244 11172
rect 27300 11116 27804 11172
rect 27860 11116 27870 11172
rect 30034 11116 30044 11172
rect 30100 11116 31276 11172
rect 31332 11116 31342 11172
rect 1708 10948 1764 11116
rect 16258 11004 16268 11060
rect 16324 11004 17276 11060
rect 17332 11004 19068 11060
rect 19124 11004 19134 11060
rect 10526 10948 10536 11004
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10800 10948 10810 11004
rect 19850 10948 19860 11004
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 20124 10948 20134 11004
rect 29174 10948 29184 11004
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29448 10948 29458 11004
rect 38498 10948 38508 11004
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38772 10948 38782 11004
rect 924 10892 1764 10948
rect 0 10836 800 10864
rect 924 10836 980 10892
rect 39200 10836 40000 10864
rect 0 10780 980 10836
rect 15474 10780 15484 10836
rect 15540 10780 16156 10836
rect 16212 10780 19404 10836
rect 19460 10780 19740 10836
rect 19796 10780 19806 10836
rect 38434 10780 38444 10836
rect 38500 10780 40000 10836
rect 0 10752 800 10780
rect 39200 10752 40000 10780
rect 2034 10668 2044 10724
rect 2100 10668 11004 10724
rect 11060 10668 11070 10724
rect 16706 10668 16716 10724
rect 16772 10668 18732 10724
rect 18788 10668 18798 10724
rect 20626 10668 20636 10724
rect 20692 10668 21756 10724
rect 21812 10668 21822 10724
rect 33506 10668 33516 10724
rect 33572 10668 37884 10724
rect 37940 10668 37950 10724
rect 24658 10556 24668 10612
rect 24724 10556 27244 10612
rect 27300 10556 29148 10612
rect 29204 10556 29214 10612
rect 23986 10332 23996 10388
rect 24052 10332 26684 10388
rect 26740 10332 26750 10388
rect 20738 10220 20748 10276
rect 20804 10220 21756 10276
rect 21812 10220 22540 10276
rect 22596 10220 22606 10276
rect 0 10164 800 10192
rect 5864 10164 5874 10220
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 6138 10164 6148 10220
rect 15188 10164 15198 10220
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15462 10164 15472 10220
rect 24512 10164 24522 10220
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24786 10164 24796 10220
rect 33836 10164 33846 10220
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 34110 10164 34120 10220
rect 39200 10164 40000 10192
rect 0 10108 1708 10164
rect 1764 10108 1774 10164
rect 18946 10108 18956 10164
rect 19012 10108 21308 10164
rect 21364 10108 21374 10164
rect 21858 10108 21868 10164
rect 21924 10108 23212 10164
rect 23268 10108 23278 10164
rect 27122 10108 27132 10164
rect 27188 10108 33068 10164
rect 33124 10108 33134 10164
rect 38210 10108 38220 10164
rect 38276 10108 40000 10164
rect 0 10080 800 10108
rect 39200 10080 40000 10108
rect 2034 9772 2044 9828
rect 2100 9772 10108 9828
rect 10164 9772 10174 9828
rect 30706 9772 30716 9828
rect 30772 9772 37884 9828
rect 37940 9772 37950 9828
rect 20514 9660 20524 9716
rect 20580 9660 22316 9716
rect 22372 9660 22382 9716
rect 23426 9660 23436 9716
rect 23492 9660 24892 9716
rect 24948 9660 25228 9716
rect 25284 9660 25294 9716
rect 25778 9660 25788 9716
rect 25844 9660 27804 9716
rect 27860 9660 31164 9716
rect 31220 9660 31230 9716
rect 1698 9548 1708 9604
rect 1764 9548 1774 9604
rect 25442 9548 25452 9604
rect 25508 9548 26124 9604
rect 26180 9548 27244 9604
rect 27300 9548 27310 9604
rect 38210 9548 38220 9604
rect 38276 9548 38948 9604
rect 0 9492 800 9520
rect 1708 9492 1764 9548
rect 0 9436 1764 9492
rect 38892 9492 38948 9548
rect 39200 9492 40000 9520
rect 38892 9436 40000 9492
rect 0 9408 800 9436
rect 10526 9380 10536 9436
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10800 9380 10810 9436
rect 19850 9380 19860 9436
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 20124 9380 20134 9436
rect 29174 9380 29184 9436
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29448 9380 29458 9436
rect 38498 9380 38508 9436
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38772 9380 38782 9436
rect 39200 9408 40000 9436
rect 23538 9212 23548 9268
rect 23604 9212 24892 9268
rect 24948 9212 24958 9268
rect 26852 9212 27468 9268
rect 27524 9212 27534 9268
rect 30594 9212 30604 9268
rect 30660 9212 36764 9268
rect 36820 9212 36830 9268
rect 2034 9100 2044 9156
rect 2100 9100 10332 9156
rect 10388 9100 10398 9156
rect 18722 9100 18732 9156
rect 18788 9100 19516 9156
rect 19572 9100 19740 9156
rect 19796 9100 19806 9156
rect 22306 9100 22316 9156
rect 22372 9100 23324 9156
rect 23380 9100 23390 9156
rect 26852 9044 26908 9212
rect 23538 8988 23548 9044
rect 23604 8988 23884 9044
rect 23940 8988 23950 9044
rect 24322 8988 24332 9044
rect 24388 8988 26908 9044
rect 0 8820 800 8848
rect 25228 8820 25284 8988
rect 39200 8820 40000 8848
rect 0 8764 1708 8820
rect 1764 8764 1774 8820
rect 22418 8764 22428 8820
rect 22484 8764 22876 8820
rect 22932 8764 24108 8820
rect 24164 8764 25004 8820
rect 25060 8764 25070 8820
rect 25218 8764 25228 8820
rect 25284 8764 25294 8820
rect 38210 8764 38220 8820
rect 38276 8764 40000 8820
rect 0 8736 800 8764
rect 39200 8736 40000 8764
rect 5864 8596 5874 8652
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 6138 8596 6148 8652
rect 15188 8596 15198 8652
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15462 8596 15472 8652
rect 24512 8596 24522 8652
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24786 8596 24796 8652
rect 33836 8596 33846 8652
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 34110 8596 34120 8652
rect 12338 8428 12348 8484
rect 12404 8428 13468 8484
rect 13524 8428 13534 8484
rect 22866 8428 22876 8484
rect 22932 8428 25340 8484
rect 25396 8428 25406 8484
rect 2594 8316 2604 8372
rect 2660 8316 3164 8372
rect 3220 8316 11228 8372
rect 11284 8316 11294 8372
rect 24658 8316 24668 8372
rect 24724 8316 25900 8372
rect 25956 8316 27244 8372
rect 27300 8316 27310 8372
rect 34514 8316 34524 8372
rect 34580 8316 37884 8372
rect 37940 8316 37950 8372
rect 23650 8204 23660 8260
rect 23716 8204 24220 8260
rect 24276 8204 24286 8260
rect 24770 8204 24780 8260
rect 24836 8204 25788 8260
rect 25844 8204 25854 8260
rect 26562 8204 26572 8260
rect 26628 8204 36428 8260
rect 36484 8204 37212 8260
rect 37268 8204 37278 8260
rect 0 8148 800 8176
rect 39200 8148 40000 8176
rect 0 8092 1708 8148
rect 1764 8092 1774 8148
rect 23090 8092 23100 8148
rect 23156 8092 24668 8148
rect 24724 8092 24734 8148
rect 38210 8092 38220 8148
rect 38276 8092 40000 8148
rect 0 8064 800 8092
rect 39200 8064 40000 8092
rect 22082 7980 22092 8036
rect 22148 7980 22876 8036
rect 22932 7980 22942 8036
rect 24546 7980 24556 8036
rect 24612 7980 26124 8036
rect 26180 7980 26190 8036
rect 26786 7980 26796 8036
rect 26852 7980 27132 8036
rect 27188 7980 34524 8036
rect 34580 7980 34590 8036
rect 23986 7868 23996 7924
rect 24052 7868 25004 7924
rect 25060 7868 25070 7924
rect 10526 7812 10536 7868
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10800 7812 10810 7868
rect 19850 7812 19860 7868
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 20124 7812 20134 7868
rect 29174 7812 29184 7868
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29448 7812 29458 7868
rect 38498 7812 38508 7868
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38772 7812 38782 7868
rect 2370 7644 2380 7700
rect 2436 7644 2446 7700
rect 0 7476 800 7504
rect 2380 7476 2436 7644
rect 32274 7532 32284 7588
rect 32340 7532 37884 7588
rect 37940 7532 37950 7588
rect 39200 7476 40000 7504
rect 0 7420 2436 7476
rect 18946 7420 18956 7476
rect 19012 7420 22988 7476
rect 23044 7420 23054 7476
rect 37538 7420 37548 7476
rect 37604 7420 40000 7476
rect 0 7392 800 7420
rect 39200 7392 40000 7420
rect 2370 7308 2380 7364
rect 2436 7308 13244 7364
rect 13300 7308 13310 7364
rect 5864 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6148 7084
rect 15188 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15472 7084
rect 24512 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24796 7084
rect 33836 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34120 7084
rect 39200 6804 40000 6832
rect 27570 6748 27580 6804
rect 27636 6748 33628 6804
rect 33684 6748 33694 6804
rect 38210 6748 38220 6804
rect 38276 6748 40000 6804
rect 39200 6720 40000 6748
rect 25106 6636 25116 6692
rect 25172 6636 29932 6692
rect 29988 6636 29998 6692
rect 36530 6636 36540 6692
rect 36596 6636 37548 6692
rect 37604 6636 37996 6692
rect 38052 6636 38062 6692
rect 25666 6524 25676 6580
rect 25732 6524 32396 6580
rect 32452 6524 32462 6580
rect 10526 6244 10536 6300
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10800 6244 10810 6300
rect 19850 6244 19860 6300
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 20124 6244 20134 6300
rect 29174 6244 29184 6300
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29448 6244 29458 6300
rect 38498 6244 38508 6300
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38772 6244 38782 6300
rect 38210 6188 38220 6244
rect 38276 6188 38286 6244
rect 38220 6132 38276 6188
rect 39200 6132 40000 6160
rect 32946 6076 32956 6132
rect 33012 6076 37660 6132
rect 37716 6076 37726 6132
rect 38220 6076 40000 6132
rect 39200 6048 40000 6076
rect 20850 5852 20860 5908
rect 20916 5852 33404 5908
rect 33460 5852 33470 5908
rect 5864 5460 5874 5516
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 6138 5460 6148 5516
rect 15188 5460 15198 5516
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15462 5460 15472 5516
rect 24512 5460 24522 5516
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24786 5460 24796 5516
rect 33836 5460 33846 5516
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 34110 5460 34120 5516
rect 39200 5460 40000 5488
rect 38210 5404 38220 5460
rect 38276 5404 40000 5460
rect 39200 5376 40000 5404
rect 36754 5180 36764 5236
rect 36820 5180 37548 5236
rect 37604 5180 37996 5236
rect 38052 5180 38062 5236
rect 25554 4956 25564 5012
rect 25620 4956 30604 5012
rect 30660 4956 30670 5012
rect 24882 4844 24892 4900
rect 24948 4844 27468 4900
rect 27524 4844 27534 4900
rect 38210 4844 38220 4900
rect 38276 4844 38948 4900
rect 38892 4788 38948 4844
rect 39200 4788 40000 4816
rect 38892 4732 40000 4788
rect 10526 4676 10536 4732
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10800 4676 10810 4732
rect 19850 4676 19860 4732
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 20124 4676 20134 4732
rect 29174 4676 29184 4732
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29448 4676 29458 4732
rect 38498 4676 38508 4732
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38772 4676 38782 4732
rect 39200 4704 40000 4732
rect 24854 4508 24892 4564
rect 24948 4508 24958 4564
rect 33394 4508 33404 4564
rect 33460 4508 33852 4564
rect 33908 4508 34412 4564
rect 34468 4508 34478 4564
rect 36082 4508 36092 4564
rect 36148 4508 37660 4564
rect 37716 4508 37726 4564
rect 39200 4116 40000 4144
rect 38210 4060 38220 4116
rect 38276 4060 40000 4116
rect 39200 4032 40000 4060
rect 5864 3892 5874 3948
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 6138 3892 6148 3948
rect 15188 3892 15198 3948
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15462 3892 15472 3948
rect 24512 3892 24522 3948
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24786 3892 24796 3948
rect 33836 3892 33846 3948
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 34110 3892 34120 3948
rect 36306 3612 36316 3668
rect 36372 3612 37548 3668
rect 37604 3612 37996 3668
rect 38052 3612 38062 3668
rect 14466 3500 14476 3556
rect 14532 3500 16044 3556
rect 16100 3500 16110 3556
rect 24210 3500 24220 3556
rect 24276 3500 25228 3556
rect 25284 3500 25294 3556
rect 39200 3444 40000 3472
rect 9538 3388 9548 3444
rect 9604 3388 10108 3444
rect 10164 3388 10174 3444
rect 24994 3388 25004 3444
rect 25060 3388 25900 3444
rect 25956 3388 25966 3444
rect 26450 3388 26460 3444
rect 26516 3388 27244 3444
rect 27300 3388 27310 3444
rect 28242 3388 28252 3444
rect 28308 3388 29036 3444
rect 29092 3388 29102 3444
rect 30930 3388 30940 3444
rect 30996 3388 32172 3444
rect 32228 3388 32238 3444
rect 32946 3388 32956 3444
rect 33012 3388 34188 3444
rect 34244 3388 34254 3444
rect 38210 3388 38220 3444
rect 38276 3388 40000 3444
rect 39200 3360 40000 3388
rect 31826 3276 31836 3332
rect 31892 3276 32844 3332
rect 32900 3276 32910 3332
rect 10526 3108 10536 3164
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10800 3108 10810 3164
rect 19850 3108 19860 3164
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 20124 3108 20134 3164
rect 29174 3108 29184 3164
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29448 3108 29458 3164
rect 38498 3108 38508 3164
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38772 3108 38782 3164
rect 32498 1932 32508 1988
rect 32564 1932 33516 1988
rect 33572 1932 33582 1988
rect 23762 1820 23772 1876
rect 23828 1820 24556 1876
rect 24612 1820 24622 1876
rect 25554 924 25564 980
rect 25620 924 26572 980
rect 26628 924 26638 980
rect 27570 924 27580 980
rect 27636 924 28364 980
rect 28420 924 28430 980
<< via3 >>
rect 5874 36820 5930 36876
rect 5978 36820 6034 36876
rect 6082 36820 6138 36876
rect 15198 36820 15254 36876
rect 15302 36820 15358 36876
rect 15406 36820 15462 36876
rect 24522 36820 24578 36876
rect 24626 36820 24682 36876
rect 24730 36820 24786 36876
rect 33846 36820 33902 36876
rect 33950 36820 34006 36876
rect 34054 36820 34110 36876
rect 10536 36036 10592 36092
rect 10640 36036 10696 36092
rect 10744 36036 10800 36092
rect 19860 36036 19916 36092
rect 19964 36036 20020 36092
rect 20068 36036 20124 36092
rect 29184 36036 29240 36092
rect 29288 36036 29344 36092
rect 29392 36036 29448 36092
rect 38508 36036 38564 36092
rect 38612 36036 38668 36092
rect 38716 36036 38772 36092
rect 5874 35252 5930 35308
rect 5978 35252 6034 35308
rect 6082 35252 6138 35308
rect 15198 35252 15254 35308
rect 15302 35252 15358 35308
rect 15406 35252 15462 35308
rect 24522 35252 24578 35308
rect 24626 35252 24682 35308
rect 24730 35252 24786 35308
rect 33846 35252 33902 35308
rect 33950 35252 34006 35308
rect 34054 35252 34110 35308
rect 10536 34468 10592 34524
rect 10640 34468 10696 34524
rect 10744 34468 10800 34524
rect 19860 34468 19916 34524
rect 19964 34468 20020 34524
rect 20068 34468 20124 34524
rect 29184 34468 29240 34524
rect 29288 34468 29344 34524
rect 29392 34468 29448 34524
rect 38508 34468 38564 34524
rect 38612 34468 38668 34524
rect 38716 34468 38772 34524
rect 5874 33684 5930 33740
rect 5978 33684 6034 33740
rect 6082 33684 6138 33740
rect 15198 33684 15254 33740
rect 15302 33684 15358 33740
rect 15406 33684 15462 33740
rect 24522 33684 24578 33740
rect 24626 33684 24682 33740
rect 24730 33684 24786 33740
rect 33846 33684 33902 33740
rect 33950 33684 34006 33740
rect 34054 33684 34110 33740
rect 10536 32900 10592 32956
rect 10640 32900 10696 32956
rect 10744 32900 10800 32956
rect 19860 32900 19916 32956
rect 19964 32900 20020 32956
rect 20068 32900 20124 32956
rect 29184 32900 29240 32956
rect 29288 32900 29344 32956
rect 29392 32900 29448 32956
rect 38508 32900 38564 32956
rect 38612 32900 38668 32956
rect 38716 32900 38772 32956
rect 5874 32116 5930 32172
rect 5978 32116 6034 32172
rect 6082 32116 6138 32172
rect 15198 32116 15254 32172
rect 15302 32116 15358 32172
rect 15406 32116 15462 32172
rect 24522 32116 24578 32172
rect 24626 32116 24682 32172
rect 24730 32116 24786 32172
rect 33846 32116 33902 32172
rect 33950 32116 34006 32172
rect 34054 32116 34110 32172
rect 10536 31332 10592 31388
rect 10640 31332 10696 31388
rect 10744 31332 10800 31388
rect 19860 31332 19916 31388
rect 19964 31332 20020 31388
rect 20068 31332 20124 31388
rect 29184 31332 29240 31388
rect 29288 31332 29344 31388
rect 29392 31332 29448 31388
rect 38508 31332 38564 31388
rect 38612 31332 38668 31388
rect 38716 31332 38772 31388
rect 5874 30548 5930 30604
rect 5978 30548 6034 30604
rect 6082 30548 6138 30604
rect 15198 30548 15254 30604
rect 15302 30548 15358 30604
rect 15406 30548 15462 30604
rect 24522 30548 24578 30604
rect 24626 30548 24682 30604
rect 24730 30548 24786 30604
rect 33846 30548 33902 30604
rect 33950 30548 34006 30604
rect 34054 30548 34110 30604
rect 10536 29764 10592 29820
rect 10640 29764 10696 29820
rect 10744 29764 10800 29820
rect 19860 29764 19916 29820
rect 19964 29764 20020 29820
rect 20068 29764 20124 29820
rect 29184 29764 29240 29820
rect 29288 29764 29344 29820
rect 29392 29764 29448 29820
rect 38508 29764 38564 29820
rect 38612 29764 38668 29820
rect 38716 29764 38772 29820
rect 19292 29372 19348 29428
rect 5874 28980 5930 29036
rect 5978 28980 6034 29036
rect 6082 28980 6138 29036
rect 15198 28980 15254 29036
rect 15302 28980 15358 29036
rect 15406 28980 15462 29036
rect 24522 28980 24578 29036
rect 24626 28980 24682 29036
rect 24730 28980 24786 29036
rect 33846 28980 33902 29036
rect 33950 28980 34006 29036
rect 34054 28980 34110 29036
rect 10536 28196 10592 28252
rect 10640 28196 10696 28252
rect 10744 28196 10800 28252
rect 19860 28196 19916 28252
rect 19964 28196 20020 28252
rect 20068 28196 20124 28252
rect 29184 28196 29240 28252
rect 29288 28196 29344 28252
rect 29392 28196 29448 28252
rect 38508 28196 38564 28252
rect 38612 28196 38668 28252
rect 38716 28196 38772 28252
rect 23212 28028 23268 28084
rect 17836 27468 17892 27524
rect 5874 27412 5930 27468
rect 5978 27412 6034 27468
rect 6082 27412 6138 27468
rect 15198 27412 15254 27468
rect 15302 27412 15358 27468
rect 15406 27412 15462 27468
rect 24522 27412 24578 27468
rect 24626 27412 24682 27468
rect 24730 27412 24786 27468
rect 33846 27412 33902 27468
rect 33950 27412 34006 27468
rect 34054 27412 34110 27468
rect 22876 27020 22932 27076
rect 17388 26908 17444 26964
rect 10536 26628 10592 26684
rect 10640 26628 10696 26684
rect 10744 26628 10800 26684
rect 19860 26628 19916 26684
rect 19964 26628 20020 26684
rect 20068 26628 20124 26684
rect 29184 26628 29240 26684
rect 29288 26628 29344 26684
rect 29392 26628 29448 26684
rect 38508 26628 38564 26684
rect 38612 26628 38668 26684
rect 38716 26628 38772 26684
rect 5874 25844 5930 25900
rect 5978 25844 6034 25900
rect 6082 25844 6138 25900
rect 15198 25844 15254 25900
rect 15302 25844 15358 25900
rect 15406 25844 15462 25900
rect 24522 25844 24578 25900
rect 24626 25844 24682 25900
rect 24730 25844 24786 25900
rect 33846 25844 33902 25900
rect 33950 25844 34006 25900
rect 34054 25844 34110 25900
rect 10536 25060 10592 25116
rect 10640 25060 10696 25116
rect 10744 25060 10800 25116
rect 19860 25060 19916 25116
rect 19964 25060 20020 25116
rect 20068 25060 20124 25116
rect 29184 25060 29240 25116
rect 29288 25060 29344 25116
rect 29392 25060 29448 25116
rect 38508 25060 38564 25116
rect 38612 25060 38668 25116
rect 38716 25060 38772 25116
rect 23212 24892 23268 24948
rect 18956 24668 19012 24724
rect 17388 24332 17444 24388
rect 22876 24332 22932 24388
rect 5874 24276 5930 24332
rect 5978 24276 6034 24332
rect 6082 24276 6138 24332
rect 15198 24276 15254 24332
rect 15302 24276 15358 24332
rect 15406 24276 15462 24332
rect 24522 24276 24578 24332
rect 24626 24276 24682 24332
rect 24730 24276 24786 24332
rect 33846 24276 33902 24332
rect 33950 24276 34006 24332
rect 34054 24276 34110 24332
rect 18956 23996 19012 24052
rect 19292 23548 19348 23604
rect 10536 23492 10592 23548
rect 10640 23492 10696 23548
rect 10744 23492 10800 23548
rect 19860 23492 19916 23548
rect 19964 23492 20020 23548
rect 20068 23492 20124 23548
rect 29184 23492 29240 23548
rect 29288 23492 29344 23548
rect 29392 23492 29448 23548
rect 38508 23492 38564 23548
rect 38612 23492 38668 23548
rect 38716 23492 38772 23548
rect 17836 23436 17892 23492
rect 18956 22876 19012 22932
rect 5874 22708 5930 22764
rect 5978 22708 6034 22764
rect 6082 22708 6138 22764
rect 15198 22708 15254 22764
rect 15302 22708 15358 22764
rect 15406 22708 15462 22764
rect 24522 22708 24578 22764
rect 24626 22708 24682 22764
rect 24730 22708 24786 22764
rect 33846 22708 33902 22764
rect 33950 22708 34006 22764
rect 34054 22708 34110 22764
rect 10536 21924 10592 21980
rect 10640 21924 10696 21980
rect 10744 21924 10800 21980
rect 19860 21924 19916 21980
rect 19964 21924 20020 21980
rect 20068 21924 20124 21980
rect 29184 21924 29240 21980
rect 29288 21924 29344 21980
rect 29392 21924 29448 21980
rect 38508 21924 38564 21980
rect 38612 21924 38668 21980
rect 38716 21924 38772 21980
rect 5874 21140 5930 21196
rect 5978 21140 6034 21196
rect 6082 21140 6138 21196
rect 15198 21140 15254 21196
rect 15302 21140 15358 21196
rect 15406 21140 15462 21196
rect 24522 21140 24578 21196
rect 24626 21140 24682 21196
rect 24730 21140 24786 21196
rect 33846 21140 33902 21196
rect 33950 21140 34006 21196
rect 34054 21140 34110 21196
rect 10536 20356 10592 20412
rect 10640 20356 10696 20412
rect 10744 20356 10800 20412
rect 19860 20356 19916 20412
rect 19964 20356 20020 20412
rect 20068 20356 20124 20412
rect 29184 20356 29240 20412
rect 29288 20356 29344 20412
rect 29392 20356 29448 20412
rect 38508 20356 38564 20412
rect 38612 20356 38668 20412
rect 38716 20356 38772 20412
rect 5874 19572 5930 19628
rect 5978 19572 6034 19628
rect 6082 19572 6138 19628
rect 15198 19572 15254 19628
rect 15302 19572 15358 19628
rect 15406 19572 15462 19628
rect 24522 19572 24578 19628
rect 24626 19572 24682 19628
rect 24730 19572 24786 19628
rect 33846 19572 33902 19628
rect 33950 19572 34006 19628
rect 34054 19572 34110 19628
rect 10536 18788 10592 18844
rect 10640 18788 10696 18844
rect 10744 18788 10800 18844
rect 19860 18788 19916 18844
rect 19964 18788 20020 18844
rect 20068 18788 20124 18844
rect 29184 18788 29240 18844
rect 29288 18788 29344 18844
rect 29392 18788 29448 18844
rect 38508 18788 38564 18844
rect 38612 18788 38668 18844
rect 38716 18788 38772 18844
rect 10108 18060 10164 18116
rect 5874 18004 5930 18060
rect 5978 18004 6034 18060
rect 6082 18004 6138 18060
rect 15198 18004 15254 18060
rect 15302 18004 15358 18060
rect 15406 18004 15462 18060
rect 24522 18004 24578 18060
rect 24626 18004 24682 18060
rect 24730 18004 24786 18060
rect 33846 18004 33902 18060
rect 33950 18004 34006 18060
rect 34054 18004 34110 18060
rect 10892 17500 10948 17556
rect 17052 17500 17108 17556
rect 10536 17220 10592 17276
rect 10640 17220 10696 17276
rect 10744 17220 10800 17276
rect 19860 17220 19916 17276
rect 19964 17220 20020 17276
rect 20068 17220 20124 17276
rect 29184 17220 29240 17276
rect 29288 17220 29344 17276
rect 29392 17220 29448 17276
rect 38508 17220 38564 17276
rect 38612 17220 38668 17276
rect 38716 17220 38772 17276
rect 10108 16492 10164 16548
rect 5874 16436 5930 16492
rect 5978 16436 6034 16492
rect 6082 16436 6138 16492
rect 15198 16436 15254 16492
rect 15302 16436 15358 16492
rect 15406 16436 15462 16492
rect 24522 16436 24578 16492
rect 24626 16436 24682 16492
rect 24730 16436 24786 16492
rect 33846 16436 33902 16492
rect 33950 16436 34006 16492
rect 34054 16436 34110 16492
rect 10892 16380 10948 16436
rect 17052 16380 17108 16436
rect 10536 15652 10592 15708
rect 10640 15652 10696 15708
rect 10744 15652 10800 15708
rect 19860 15652 19916 15708
rect 19964 15652 20020 15708
rect 20068 15652 20124 15708
rect 29184 15652 29240 15708
rect 29288 15652 29344 15708
rect 29392 15652 29448 15708
rect 38508 15652 38564 15708
rect 38612 15652 38668 15708
rect 38716 15652 38772 15708
rect 15596 15148 15652 15204
rect 5874 14868 5930 14924
rect 5978 14868 6034 14924
rect 6082 14868 6138 14924
rect 15198 14868 15254 14924
rect 15302 14868 15358 14924
rect 15406 14868 15462 14924
rect 24522 14868 24578 14924
rect 24626 14868 24682 14924
rect 24730 14868 24786 14924
rect 33846 14868 33902 14924
rect 33950 14868 34006 14924
rect 34054 14868 34110 14924
rect 10332 14812 10388 14868
rect 15596 14588 15652 14644
rect 10536 14084 10592 14140
rect 10640 14084 10696 14140
rect 10744 14084 10800 14140
rect 19860 14084 19916 14140
rect 19964 14084 20020 14140
rect 20068 14084 20124 14140
rect 29184 14084 29240 14140
rect 29288 14084 29344 14140
rect 29392 14084 29448 14140
rect 38508 14084 38564 14140
rect 38612 14084 38668 14140
rect 38716 14084 38772 14140
rect 10332 13916 10388 13972
rect 5874 13300 5930 13356
rect 5978 13300 6034 13356
rect 6082 13300 6138 13356
rect 15198 13300 15254 13356
rect 15302 13300 15358 13356
rect 15406 13300 15462 13356
rect 24522 13300 24578 13356
rect 24626 13300 24682 13356
rect 24730 13300 24786 13356
rect 33846 13300 33902 13356
rect 33950 13300 34006 13356
rect 34054 13300 34110 13356
rect 10536 12516 10592 12572
rect 10640 12516 10696 12572
rect 10744 12516 10800 12572
rect 19860 12516 19916 12572
rect 19964 12516 20020 12572
rect 20068 12516 20124 12572
rect 29184 12516 29240 12572
rect 29288 12516 29344 12572
rect 29392 12516 29448 12572
rect 38508 12516 38564 12572
rect 38612 12516 38668 12572
rect 38716 12516 38772 12572
rect 5874 11732 5930 11788
rect 5978 11732 6034 11788
rect 6082 11732 6138 11788
rect 15198 11732 15254 11788
rect 15302 11732 15358 11788
rect 15406 11732 15462 11788
rect 24522 11732 24578 11788
rect 24626 11732 24682 11788
rect 24730 11732 24786 11788
rect 33846 11732 33902 11788
rect 33950 11732 34006 11788
rect 34054 11732 34110 11788
rect 10536 10948 10592 11004
rect 10640 10948 10696 11004
rect 10744 10948 10800 11004
rect 19860 10948 19916 11004
rect 19964 10948 20020 11004
rect 20068 10948 20124 11004
rect 29184 10948 29240 11004
rect 29288 10948 29344 11004
rect 29392 10948 29448 11004
rect 38508 10948 38564 11004
rect 38612 10948 38668 11004
rect 38716 10948 38772 11004
rect 5874 10164 5930 10220
rect 5978 10164 6034 10220
rect 6082 10164 6138 10220
rect 15198 10164 15254 10220
rect 15302 10164 15358 10220
rect 15406 10164 15462 10220
rect 24522 10164 24578 10220
rect 24626 10164 24682 10220
rect 24730 10164 24786 10220
rect 33846 10164 33902 10220
rect 33950 10164 34006 10220
rect 34054 10164 34110 10220
rect 10536 9380 10592 9436
rect 10640 9380 10696 9436
rect 10744 9380 10800 9436
rect 19860 9380 19916 9436
rect 19964 9380 20020 9436
rect 20068 9380 20124 9436
rect 29184 9380 29240 9436
rect 29288 9380 29344 9436
rect 29392 9380 29448 9436
rect 38508 9380 38564 9436
rect 38612 9380 38668 9436
rect 38716 9380 38772 9436
rect 24892 9212 24948 9268
rect 5874 8596 5930 8652
rect 5978 8596 6034 8652
rect 6082 8596 6138 8652
rect 15198 8596 15254 8652
rect 15302 8596 15358 8652
rect 15406 8596 15462 8652
rect 24522 8596 24578 8652
rect 24626 8596 24682 8652
rect 24730 8596 24786 8652
rect 33846 8596 33902 8652
rect 33950 8596 34006 8652
rect 34054 8596 34110 8652
rect 10536 7812 10592 7868
rect 10640 7812 10696 7868
rect 10744 7812 10800 7868
rect 19860 7812 19916 7868
rect 19964 7812 20020 7868
rect 20068 7812 20124 7868
rect 29184 7812 29240 7868
rect 29288 7812 29344 7868
rect 29392 7812 29448 7868
rect 38508 7812 38564 7868
rect 38612 7812 38668 7868
rect 38716 7812 38772 7868
rect 5874 7028 5930 7084
rect 5978 7028 6034 7084
rect 6082 7028 6138 7084
rect 15198 7028 15254 7084
rect 15302 7028 15358 7084
rect 15406 7028 15462 7084
rect 24522 7028 24578 7084
rect 24626 7028 24682 7084
rect 24730 7028 24786 7084
rect 33846 7028 33902 7084
rect 33950 7028 34006 7084
rect 34054 7028 34110 7084
rect 10536 6244 10592 6300
rect 10640 6244 10696 6300
rect 10744 6244 10800 6300
rect 19860 6244 19916 6300
rect 19964 6244 20020 6300
rect 20068 6244 20124 6300
rect 29184 6244 29240 6300
rect 29288 6244 29344 6300
rect 29392 6244 29448 6300
rect 38508 6244 38564 6300
rect 38612 6244 38668 6300
rect 38716 6244 38772 6300
rect 5874 5460 5930 5516
rect 5978 5460 6034 5516
rect 6082 5460 6138 5516
rect 15198 5460 15254 5516
rect 15302 5460 15358 5516
rect 15406 5460 15462 5516
rect 24522 5460 24578 5516
rect 24626 5460 24682 5516
rect 24730 5460 24786 5516
rect 33846 5460 33902 5516
rect 33950 5460 34006 5516
rect 34054 5460 34110 5516
rect 10536 4676 10592 4732
rect 10640 4676 10696 4732
rect 10744 4676 10800 4732
rect 19860 4676 19916 4732
rect 19964 4676 20020 4732
rect 20068 4676 20124 4732
rect 29184 4676 29240 4732
rect 29288 4676 29344 4732
rect 29392 4676 29448 4732
rect 38508 4676 38564 4732
rect 38612 4676 38668 4732
rect 38716 4676 38772 4732
rect 24892 4508 24948 4564
rect 5874 3892 5930 3948
rect 5978 3892 6034 3948
rect 6082 3892 6138 3948
rect 15198 3892 15254 3948
rect 15302 3892 15358 3948
rect 15406 3892 15462 3948
rect 24522 3892 24578 3948
rect 24626 3892 24682 3948
rect 24730 3892 24786 3948
rect 33846 3892 33902 3948
rect 33950 3892 34006 3948
rect 34054 3892 34110 3948
rect 10536 3108 10592 3164
rect 10640 3108 10696 3164
rect 10744 3108 10800 3164
rect 19860 3108 19916 3164
rect 19964 3108 20020 3164
rect 20068 3108 20124 3164
rect 29184 3108 29240 3164
rect 29288 3108 29344 3164
rect 29392 3108 29448 3164
rect 38508 3108 38564 3164
rect 38612 3108 38668 3164
rect 38716 3108 38772 3164
<< metal4 >>
rect 5846 36876 6166 36908
rect 5846 36820 5874 36876
rect 5930 36820 5978 36876
rect 6034 36820 6082 36876
rect 6138 36820 6166 36876
rect 5846 35308 6166 36820
rect 5846 35252 5874 35308
rect 5930 35252 5978 35308
rect 6034 35252 6082 35308
rect 6138 35252 6166 35308
rect 5846 33740 6166 35252
rect 5846 33684 5874 33740
rect 5930 33684 5978 33740
rect 6034 33684 6082 33740
rect 6138 33684 6166 33740
rect 5846 32172 6166 33684
rect 5846 32116 5874 32172
rect 5930 32116 5978 32172
rect 6034 32116 6082 32172
rect 6138 32116 6166 32172
rect 5846 30604 6166 32116
rect 5846 30548 5874 30604
rect 5930 30548 5978 30604
rect 6034 30548 6082 30604
rect 6138 30548 6166 30604
rect 5846 29036 6166 30548
rect 5846 28980 5874 29036
rect 5930 28980 5978 29036
rect 6034 28980 6082 29036
rect 6138 28980 6166 29036
rect 5846 27468 6166 28980
rect 5846 27412 5874 27468
rect 5930 27412 5978 27468
rect 6034 27412 6082 27468
rect 6138 27412 6166 27468
rect 5846 25900 6166 27412
rect 5846 25844 5874 25900
rect 5930 25844 5978 25900
rect 6034 25844 6082 25900
rect 6138 25844 6166 25900
rect 5846 24332 6166 25844
rect 5846 24276 5874 24332
rect 5930 24276 5978 24332
rect 6034 24276 6082 24332
rect 6138 24276 6166 24332
rect 5846 22764 6166 24276
rect 5846 22708 5874 22764
rect 5930 22708 5978 22764
rect 6034 22708 6082 22764
rect 6138 22708 6166 22764
rect 5846 21196 6166 22708
rect 5846 21140 5874 21196
rect 5930 21140 5978 21196
rect 6034 21140 6082 21196
rect 6138 21140 6166 21196
rect 5846 19628 6166 21140
rect 5846 19572 5874 19628
rect 5930 19572 5978 19628
rect 6034 19572 6082 19628
rect 6138 19572 6166 19628
rect 5846 18060 6166 19572
rect 10508 36092 10828 36908
rect 10508 36036 10536 36092
rect 10592 36036 10640 36092
rect 10696 36036 10744 36092
rect 10800 36036 10828 36092
rect 10508 34524 10828 36036
rect 10508 34468 10536 34524
rect 10592 34468 10640 34524
rect 10696 34468 10744 34524
rect 10800 34468 10828 34524
rect 10508 32956 10828 34468
rect 10508 32900 10536 32956
rect 10592 32900 10640 32956
rect 10696 32900 10744 32956
rect 10800 32900 10828 32956
rect 10508 31388 10828 32900
rect 10508 31332 10536 31388
rect 10592 31332 10640 31388
rect 10696 31332 10744 31388
rect 10800 31332 10828 31388
rect 10508 29820 10828 31332
rect 10508 29764 10536 29820
rect 10592 29764 10640 29820
rect 10696 29764 10744 29820
rect 10800 29764 10828 29820
rect 10508 28252 10828 29764
rect 10508 28196 10536 28252
rect 10592 28196 10640 28252
rect 10696 28196 10744 28252
rect 10800 28196 10828 28252
rect 10508 26684 10828 28196
rect 10508 26628 10536 26684
rect 10592 26628 10640 26684
rect 10696 26628 10744 26684
rect 10800 26628 10828 26684
rect 10508 25116 10828 26628
rect 10508 25060 10536 25116
rect 10592 25060 10640 25116
rect 10696 25060 10744 25116
rect 10800 25060 10828 25116
rect 10508 23548 10828 25060
rect 10508 23492 10536 23548
rect 10592 23492 10640 23548
rect 10696 23492 10744 23548
rect 10800 23492 10828 23548
rect 10508 21980 10828 23492
rect 10508 21924 10536 21980
rect 10592 21924 10640 21980
rect 10696 21924 10744 21980
rect 10800 21924 10828 21980
rect 10508 20412 10828 21924
rect 10508 20356 10536 20412
rect 10592 20356 10640 20412
rect 10696 20356 10744 20412
rect 10800 20356 10828 20412
rect 10508 18844 10828 20356
rect 10508 18788 10536 18844
rect 10592 18788 10640 18844
rect 10696 18788 10744 18844
rect 10800 18788 10828 18844
rect 5846 18004 5874 18060
rect 5930 18004 5978 18060
rect 6034 18004 6082 18060
rect 6138 18004 6166 18060
rect 5846 16492 6166 18004
rect 5846 16436 5874 16492
rect 5930 16436 5978 16492
rect 6034 16436 6082 16492
rect 6138 16436 6166 16492
rect 10108 18116 10164 18126
rect 10108 16548 10164 18060
rect 10108 16482 10164 16492
rect 10508 17276 10828 18788
rect 15170 36876 15490 36908
rect 15170 36820 15198 36876
rect 15254 36820 15302 36876
rect 15358 36820 15406 36876
rect 15462 36820 15490 36876
rect 15170 35308 15490 36820
rect 15170 35252 15198 35308
rect 15254 35252 15302 35308
rect 15358 35252 15406 35308
rect 15462 35252 15490 35308
rect 15170 33740 15490 35252
rect 15170 33684 15198 33740
rect 15254 33684 15302 33740
rect 15358 33684 15406 33740
rect 15462 33684 15490 33740
rect 15170 32172 15490 33684
rect 15170 32116 15198 32172
rect 15254 32116 15302 32172
rect 15358 32116 15406 32172
rect 15462 32116 15490 32172
rect 15170 30604 15490 32116
rect 15170 30548 15198 30604
rect 15254 30548 15302 30604
rect 15358 30548 15406 30604
rect 15462 30548 15490 30604
rect 15170 29036 15490 30548
rect 19832 36092 20152 36908
rect 19832 36036 19860 36092
rect 19916 36036 19964 36092
rect 20020 36036 20068 36092
rect 20124 36036 20152 36092
rect 19832 34524 20152 36036
rect 19832 34468 19860 34524
rect 19916 34468 19964 34524
rect 20020 34468 20068 34524
rect 20124 34468 20152 34524
rect 19832 32956 20152 34468
rect 19832 32900 19860 32956
rect 19916 32900 19964 32956
rect 20020 32900 20068 32956
rect 20124 32900 20152 32956
rect 19832 31388 20152 32900
rect 19832 31332 19860 31388
rect 19916 31332 19964 31388
rect 20020 31332 20068 31388
rect 20124 31332 20152 31388
rect 19832 29820 20152 31332
rect 19832 29764 19860 29820
rect 19916 29764 19964 29820
rect 20020 29764 20068 29820
rect 20124 29764 20152 29820
rect 15170 28980 15198 29036
rect 15254 28980 15302 29036
rect 15358 28980 15406 29036
rect 15462 28980 15490 29036
rect 15170 27468 15490 28980
rect 19292 29428 19348 29438
rect 15170 27412 15198 27468
rect 15254 27412 15302 27468
rect 15358 27412 15406 27468
rect 15462 27412 15490 27468
rect 15170 25900 15490 27412
rect 17836 27524 17892 27534
rect 15170 25844 15198 25900
rect 15254 25844 15302 25900
rect 15358 25844 15406 25900
rect 15462 25844 15490 25900
rect 15170 24332 15490 25844
rect 15170 24276 15198 24332
rect 15254 24276 15302 24332
rect 15358 24276 15406 24332
rect 15462 24276 15490 24332
rect 17388 26964 17444 26974
rect 17388 24388 17444 26908
rect 17388 24322 17444 24332
rect 15170 22764 15490 24276
rect 17836 23492 17892 27468
rect 17836 23426 17892 23436
rect 18956 24724 19012 24734
rect 18956 24052 19012 24668
rect 18956 22932 19012 23996
rect 19292 23604 19348 29372
rect 19292 23538 19348 23548
rect 19832 28252 20152 29764
rect 19832 28196 19860 28252
rect 19916 28196 19964 28252
rect 20020 28196 20068 28252
rect 20124 28196 20152 28252
rect 19832 26684 20152 28196
rect 24494 36876 24814 36908
rect 24494 36820 24522 36876
rect 24578 36820 24626 36876
rect 24682 36820 24730 36876
rect 24786 36820 24814 36876
rect 24494 35308 24814 36820
rect 24494 35252 24522 35308
rect 24578 35252 24626 35308
rect 24682 35252 24730 35308
rect 24786 35252 24814 35308
rect 24494 33740 24814 35252
rect 24494 33684 24522 33740
rect 24578 33684 24626 33740
rect 24682 33684 24730 33740
rect 24786 33684 24814 33740
rect 24494 32172 24814 33684
rect 24494 32116 24522 32172
rect 24578 32116 24626 32172
rect 24682 32116 24730 32172
rect 24786 32116 24814 32172
rect 24494 30604 24814 32116
rect 24494 30548 24522 30604
rect 24578 30548 24626 30604
rect 24682 30548 24730 30604
rect 24786 30548 24814 30604
rect 24494 29036 24814 30548
rect 24494 28980 24522 29036
rect 24578 28980 24626 29036
rect 24682 28980 24730 29036
rect 24786 28980 24814 29036
rect 23212 28084 23268 28094
rect 19832 26628 19860 26684
rect 19916 26628 19964 26684
rect 20020 26628 20068 26684
rect 20124 26628 20152 26684
rect 19832 25116 20152 26628
rect 19832 25060 19860 25116
rect 19916 25060 19964 25116
rect 20020 25060 20068 25116
rect 20124 25060 20152 25116
rect 19832 23548 20152 25060
rect 22876 27076 22932 27086
rect 22876 24388 22932 27020
rect 23212 24948 23268 28028
rect 23212 24882 23268 24892
rect 24494 27468 24814 28980
rect 24494 27412 24522 27468
rect 24578 27412 24626 27468
rect 24682 27412 24730 27468
rect 24786 27412 24814 27468
rect 24494 25900 24814 27412
rect 24494 25844 24522 25900
rect 24578 25844 24626 25900
rect 24682 25844 24730 25900
rect 24786 25844 24814 25900
rect 22876 24322 22932 24332
rect 24494 24332 24814 25844
rect 18956 22866 19012 22876
rect 19832 23492 19860 23548
rect 19916 23492 19964 23548
rect 20020 23492 20068 23548
rect 20124 23492 20152 23548
rect 15170 22708 15198 22764
rect 15254 22708 15302 22764
rect 15358 22708 15406 22764
rect 15462 22708 15490 22764
rect 15170 21196 15490 22708
rect 15170 21140 15198 21196
rect 15254 21140 15302 21196
rect 15358 21140 15406 21196
rect 15462 21140 15490 21196
rect 15170 19628 15490 21140
rect 15170 19572 15198 19628
rect 15254 19572 15302 19628
rect 15358 19572 15406 19628
rect 15462 19572 15490 19628
rect 15170 18060 15490 19572
rect 15170 18004 15198 18060
rect 15254 18004 15302 18060
rect 15358 18004 15406 18060
rect 15462 18004 15490 18060
rect 10508 17220 10536 17276
rect 10592 17220 10640 17276
rect 10696 17220 10744 17276
rect 10800 17220 10828 17276
rect 5846 14924 6166 16436
rect 5846 14868 5874 14924
rect 5930 14868 5978 14924
rect 6034 14868 6082 14924
rect 6138 14868 6166 14924
rect 10508 15708 10828 17220
rect 10892 17556 10948 17566
rect 10892 16436 10948 17500
rect 10892 16370 10948 16380
rect 15170 16492 15490 18004
rect 19832 21980 20152 23492
rect 19832 21924 19860 21980
rect 19916 21924 19964 21980
rect 20020 21924 20068 21980
rect 20124 21924 20152 21980
rect 19832 20412 20152 21924
rect 19832 20356 19860 20412
rect 19916 20356 19964 20412
rect 20020 20356 20068 20412
rect 20124 20356 20152 20412
rect 19832 18844 20152 20356
rect 19832 18788 19860 18844
rect 19916 18788 19964 18844
rect 20020 18788 20068 18844
rect 20124 18788 20152 18844
rect 15170 16436 15198 16492
rect 15254 16436 15302 16492
rect 15358 16436 15406 16492
rect 15462 16436 15490 16492
rect 10508 15652 10536 15708
rect 10592 15652 10640 15708
rect 10696 15652 10744 15708
rect 10800 15652 10828 15708
rect 5846 13356 6166 14868
rect 10332 14868 10388 14878
rect 10332 13972 10388 14812
rect 10332 13906 10388 13916
rect 10508 14140 10828 15652
rect 10508 14084 10536 14140
rect 10592 14084 10640 14140
rect 10696 14084 10744 14140
rect 10800 14084 10828 14140
rect 5846 13300 5874 13356
rect 5930 13300 5978 13356
rect 6034 13300 6082 13356
rect 6138 13300 6166 13356
rect 5846 11788 6166 13300
rect 5846 11732 5874 11788
rect 5930 11732 5978 11788
rect 6034 11732 6082 11788
rect 6138 11732 6166 11788
rect 5846 10220 6166 11732
rect 5846 10164 5874 10220
rect 5930 10164 5978 10220
rect 6034 10164 6082 10220
rect 6138 10164 6166 10220
rect 5846 8652 6166 10164
rect 5846 8596 5874 8652
rect 5930 8596 5978 8652
rect 6034 8596 6082 8652
rect 6138 8596 6166 8652
rect 5846 7084 6166 8596
rect 5846 7028 5874 7084
rect 5930 7028 5978 7084
rect 6034 7028 6082 7084
rect 6138 7028 6166 7084
rect 5846 5516 6166 7028
rect 5846 5460 5874 5516
rect 5930 5460 5978 5516
rect 6034 5460 6082 5516
rect 6138 5460 6166 5516
rect 5846 3948 6166 5460
rect 5846 3892 5874 3948
rect 5930 3892 5978 3948
rect 6034 3892 6082 3948
rect 6138 3892 6166 3948
rect 5846 3076 6166 3892
rect 10508 12572 10828 14084
rect 10508 12516 10536 12572
rect 10592 12516 10640 12572
rect 10696 12516 10744 12572
rect 10800 12516 10828 12572
rect 10508 11004 10828 12516
rect 10508 10948 10536 11004
rect 10592 10948 10640 11004
rect 10696 10948 10744 11004
rect 10800 10948 10828 11004
rect 10508 9436 10828 10948
rect 10508 9380 10536 9436
rect 10592 9380 10640 9436
rect 10696 9380 10744 9436
rect 10800 9380 10828 9436
rect 10508 7868 10828 9380
rect 10508 7812 10536 7868
rect 10592 7812 10640 7868
rect 10696 7812 10744 7868
rect 10800 7812 10828 7868
rect 10508 6300 10828 7812
rect 10508 6244 10536 6300
rect 10592 6244 10640 6300
rect 10696 6244 10744 6300
rect 10800 6244 10828 6300
rect 10508 4732 10828 6244
rect 10508 4676 10536 4732
rect 10592 4676 10640 4732
rect 10696 4676 10744 4732
rect 10800 4676 10828 4732
rect 10508 3164 10828 4676
rect 10508 3108 10536 3164
rect 10592 3108 10640 3164
rect 10696 3108 10744 3164
rect 10800 3108 10828 3164
rect 10508 3076 10828 3108
rect 15170 14924 15490 16436
rect 17052 17556 17108 17566
rect 17052 16436 17108 17500
rect 17052 16370 17108 16380
rect 19832 17276 20152 18788
rect 19832 17220 19860 17276
rect 19916 17220 19964 17276
rect 20020 17220 20068 17276
rect 20124 17220 20152 17276
rect 19832 15708 20152 17220
rect 19832 15652 19860 15708
rect 19916 15652 19964 15708
rect 20020 15652 20068 15708
rect 20124 15652 20152 15708
rect 15170 14868 15198 14924
rect 15254 14868 15302 14924
rect 15358 14868 15406 14924
rect 15462 14868 15490 14924
rect 15170 13356 15490 14868
rect 15596 15204 15652 15214
rect 15596 14644 15652 15148
rect 15596 14578 15652 14588
rect 15170 13300 15198 13356
rect 15254 13300 15302 13356
rect 15358 13300 15406 13356
rect 15462 13300 15490 13356
rect 15170 11788 15490 13300
rect 15170 11732 15198 11788
rect 15254 11732 15302 11788
rect 15358 11732 15406 11788
rect 15462 11732 15490 11788
rect 15170 10220 15490 11732
rect 15170 10164 15198 10220
rect 15254 10164 15302 10220
rect 15358 10164 15406 10220
rect 15462 10164 15490 10220
rect 15170 8652 15490 10164
rect 15170 8596 15198 8652
rect 15254 8596 15302 8652
rect 15358 8596 15406 8652
rect 15462 8596 15490 8652
rect 15170 7084 15490 8596
rect 15170 7028 15198 7084
rect 15254 7028 15302 7084
rect 15358 7028 15406 7084
rect 15462 7028 15490 7084
rect 15170 5516 15490 7028
rect 15170 5460 15198 5516
rect 15254 5460 15302 5516
rect 15358 5460 15406 5516
rect 15462 5460 15490 5516
rect 15170 3948 15490 5460
rect 15170 3892 15198 3948
rect 15254 3892 15302 3948
rect 15358 3892 15406 3948
rect 15462 3892 15490 3948
rect 15170 3076 15490 3892
rect 19832 14140 20152 15652
rect 19832 14084 19860 14140
rect 19916 14084 19964 14140
rect 20020 14084 20068 14140
rect 20124 14084 20152 14140
rect 19832 12572 20152 14084
rect 19832 12516 19860 12572
rect 19916 12516 19964 12572
rect 20020 12516 20068 12572
rect 20124 12516 20152 12572
rect 19832 11004 20152 12516
rect 19832 10948 19860 11004
rect 19916 10948 19964 11004
rect 20020 10948 20068 11004
rect 20124 10948 20152 11004
rect 19832 9436 20152 10948
rect 19832 9380 19860 9436
rect 19916 9380 19964 9436
rect 20020 9380 20068 9436
rect 20124 9380 20152 9436
rect 19832 7868 20152 9380
rect 19832 7812 19860 7868
rect 19916 7812 19964 7868
rect 20020 7812 20068 7868
rect 20124 7812 20152 7868
rect 19832 6300 20152 7812
rect 19832 6244 19860 6300
rect 19916 6244 19964 6300
rect 20020 6244 20068 6300
rect 20124 6244 20152 6300
rect 19832 4732 20152 6244
rect 19832 4676 19860 4732
rect 19916 4676 19964 4732
rect 20020 4676 20068 4732
rect 20124 4676 20152 4732
rect 19832 3164 20152 4676
rect 19832 3108 19860 3164
rect 19916 3108 19964 3164
rect 20020 3108 20068 3164
rect 20124 3108 20152 3164
rect 19832 3076 20152 3108
rect 24494 24276 24522 24332
rect 24578 24276 24626 24332
rect 24682 24276 24730 24332
rect 24786 24276 24814 24332
rect 24494 22764 24814 24276
rect 24494 22708 24522 22764
rect 24578 22708 24626 22764
rect 24682 22708 24730 22764
rect 24786 22708 24814 22764
rect 24494 21196 24814 22708
rect 24494 21140 24522 21196
rect 24578 21140 24626 21196
rect 24682 21140 24730 21196
rect 24786 21140 24814 21196
rect 24494 19628 24814 21140
rect 24494 19572 24522 19628
rect 24578 19572 24626 19628
rect 24682 19572 24730 19628
rect 24786 19572 24814 19628
rect 24494 18060 24814 19572
rect 24494 18004 24522 18060
rect 24578 18004 24626 18060
rect 24682 18004 24730 18060
rect 24786 18004 24814 18060
rect 24494 16492 24814 18004
rect 24494 16436 24522 16492
rect 24578 16436 24626 16492
rect 24682 16436 24730 16492
rect 24786 16436 24814 16492
rect 24494 14924 24814 16436
rect 24494 14868 24522 14924
rect 24578 14868 24626 14924
rect 24682 14868 24730 14924
rect 24786 14868 24814 14924
rect 24494 13356 24814 14868
rect 24494 13300 24522 13356
rect 24578 13300 24626 13356
rect 24682 13300 24730 13356
rect 24786 13300 24814 13356
rect 24494 11788 24814 13300
rect 24494 11732 24522 11788
rect 24578 11732 24626 11788
rect 24682 11732 24730 11788
rect 24786 11732 24814 11788
rect 24494 10220 24814 11732
rect 24494 10164 24522 10220
rect 24578 10164 24626 10220
rect 24682 10164 24730 10220
rect 24786 10164 24814 10220
rect 24494 8652 24814 10164
rect 29156 36092 29476 36908
rect 29156 36036 29184 36092
rect 29240 36036 29288 36092
rect 29344 36036 29392 36092
rect 29448 36036 29476 36092
rect 29156 34524 29476 36036
rect 29156 34468 29184 34524
rect 29240 34468 29288 34524
rect 29344 34468 29392 34524
rect 29448 34468 29476 34524
rect 29156 32956 29476 34468
rect 29156 32900 29184 32956
rect 29240 32900 29288 32956
rect 29344 32900 29392 32956
rect 29448 32900 29476 32956
rect 29156 31388 29476 32900
rect 29156 31332 29184 31388
rect 29240 31332 29288 31388
rect 29344 31332 29392 31388
rect 29448 31332 29476 31388
rect 29156 29820 29476 31332
rect 29156 29764 29184 29820
rect 29240 29764 29288 29820
rect 29344 29764 29392 29820
rect 29448 29764 29476 29820
rect 29156 28252 29476 29764
rect 29156 28196 29184 28252
rect 29240 28196 29288 28252
rect 29344 28196 29392 28252
rect 29448 28196 29476 28252
rect 29156 26684 29476 28196
rect 29156 26628 29184 26684
rect 29240 26628 29288 26684
rect 29344 26628 29392 26684
rect 29448 26628 29476 26684
rect 29156 25116 29476 26628
rect 29156 25060 29184 25116
rect 29240 25060 29288 25116
rect 29344 25060 29392 25116
rect 29448 25060 29476 25116
rect 29156 23548 29476 25060
rect 29156 23492 29184 23548
rect 29240 23492 29288 23548
rect 29344 23492 29392 23548
rect 29448 23492 29476 23548
rect 29156 21980 29476 23492
rect 29156 21924 29184 21980
rect 29240 21924 29288 21980
rect 29344 21924 29392 21980
rect 29448 21924 29476 21980
rect 29156 20412 29476 21924
rect 29156 20356 29184 20412
rect 29240 20356 29288 20412
rect 29344 20356 29392 20412
rect 29448 20356 29476 20412
rect 29156 18844 29476 20356
rect 29156 18788 29184 18844
rect 29240 18788 29288 18844
rect 29344 18788 29392 18844
rect 29448 18788 29476 18844
rect 29156 17276 29476 18788
rect 29156 17220 29184 17276
rect 29240 17220 29288 17276
rect 29344 17220 29392 17276
rect 29448 17220 29476 17276
rect 29156 15708 29476 17220
rect 29156 15652 29184 15708
rect 29240 15652 29288 15708
rect 29344 15652 29392 15708
rect 29448 15652 29476 15708
rect 29156 14140 29476 15652
rect 29156 14084 29184 14140
rect 29240 14084 29288 14140
rect 29344 14084 29392 14140
rect 29448 14084 29476 14140
rect 29156 12572 29476 14084
rect 29156 12516 29184 12572
rect 29240 12516 29288 12572
rect 29344 12516 29392 12572
rect 29448 12516 29476 12572
rect 29156 11004 29476 12516
rect 29156 10948 29184 11004
rect 29240 10948 29288 11004
rect 29344 10948 29392 11004
rect 29448 10948 29476 11004
rect 29156 9436 29476 10948
rect 29156 9380 29184 9436
rect 29240 9380 29288 9436
rect 29344 9380 29392 9436
rect 29448 9380 29476 9436
rect 24494 8596 24522 8652
rect 24578 8596 24626 8652
rect 24682 8596 24730 8652
rect 24786 8596 24814 8652
rect 24494 7084 24814 8596
rect 24494 7028 24522 7084
rect 24578 7028 24626 7084
rect 24682 7028 24730 7084
rect 24786 7028 24814 7084
rect 24494 5516 24814 7028
rect 24494 5460 24522 5516
rect 24578 5460 24626 5516
rect 24682 5460 24730 5516
rect 24786 5460 24814 5516
rect 24494 3948 24814 5460
rect 24892 9268 24948 9278
rect 24892 4564 24948 9212
rect 24892 4498 24948 4508
rect 29156 7868 29476 9380
rect 29156 7812 29184 7868
rect 29240 7812 29288 7868
rect 29344 7812 29392 7868
rect 29448 7812 29476 7868
rect 29156 6300 29476 7812
rect 29156 6244 29184 6300
rect 29240 6244 29288 6300
rect 29344 6244 29392 6300
rect 29448 6244 29476 6300
rect 29156 4732 29476 6244
rect 29156 4676 29184 4732
rect 29240 4676 29288 4732
rect 29344 4676 29392 4732
rect 29448 4676 29476 4732
rect 24494 3892 24522 3948
rect 24578 3892 24626 3948
rect 24682 3892 24730 3948
rect 24786 3892 24814 3948
rect 24494 3076 24814 3892
rect 29156 3164 29476 4676
rect 29156 3108 29184 3164
rect 29240 3108 29288 3164
rect 29344 3108 29392 3164
rect 29448 3108 29476 3164
rect 29156 3076 29476 3108
rect 33818 36876 34138 36908
rect 33818 36820 33846 36876
rect 33902 36820 33950 36876
rect 34006 36820 34054 36876
rect 34110 36820 34138 36876
rect 33818 35308 34138 36820
rect 33818 35252 33846 35308
rect 33902 35252 33950 35308
rect 34006 35252 34054 35308
rect 34110 35252 34138 35308
rect 33818 33740 34138 35252
rect 33818 33684 33846 33740
rect 33902 33684 33950 33740
rect 34006 33684 34054 33740
rect 34110 33684 34138 33740
rect 33818 32172 34138 33684
rect 33818 32116 33846 32172
rect 33902 32116 33950 32172
rect 34006 32116 34054 32172
rect 34110 32116 34138 32172
rect 33818 30604 34138 32116
rect 33818 30548 33846 30604
rect 33902 30548 33950 30604
rect 34006 30548 34054 30604
rect 34110 30548 34138 30604
rect 33818 29036 34138 30548
rect 33818 28980 33846 29036
rect 33902 28980 33950 29036
rect 34006 28980 34054 29036
rect 34110 28980 34138 29036
rect 33818 27468 34138 28980
rect 33818 27412 33846 27468
rect 33902 27412 33950 27468
rect 34006 27412 34054 27468
rect 34110 27412 34138 27468
rect 33818 25900 34138 27412
rect 33818 25844 33846 25900
rect 33902 25844 33950 25900
rect 34006 25844 34054 25900
rect 34110 25844 34138 25900
rect 33818 24332 34138 25844
rect 33818 24276 33846 24332
rect 33902 24276 33950 24332
rect 34006 24276 34054 24332
rect 34110 24276 34138 24332
rect 33818 22764 34138 24276
rect 33818 22708 33846 22764
rect 33902 22708 33950 22764
rect 34006 22708 34054 22764
rect 34110 22708 34138 22764
rect 33818 21196 34138 22708
rect 33818 21140 33846 21196
rect 33902 21140 33950 21196
rect 34006 21140 34054 21196
rect 34110 21140 34138 21196
rect 33818 19628 34138 21140
rect 33818 19572 33846 19628
rect 33902 19572 33950 19628
rect 34006 19572 34054 19628
rect 34110 19572 34138 19628
rect 33818 18060 34138 19572
rect 33818 18004 33846 18060
rect 33902 18004 33950 18060
rect 34006 18004 34054 18060
rect 34110 18004 34138 18060
rect 33818 16492 34138 18004
rect 33818 16436 33846 16492
rect 33902 16436 33950 16492
rect 34006 16436 34054 16492
rect 34110 16436 34138 16492
rect 33818 14924 34138 16436
rect 33818 14868 33846 14924
rect 33902 14868 33950 14924
rect 34006 14868 34054 14924
rect 34110 14868 34138 14924
rect 33818 13356 34138 14868
rect 33818 13300 33846 13356
rect 33902 13300 33950 13356
rect 34006 13300 34054 13356
rect 34110 13300 34138 13356
rect 33818 11788 34138 13300
rect 33818 11732 33846 11788
rect 33902 11732 33950 11788
rect 34006 11732 34054 11788
rect 34110 11732 34138 11788
rect 33818 10220 34138 11732
rect 33818 10164 33846 10220
rect 33902 10164 33950 10220
rect 34006 10164 34054 10220
rect 34110 10164 34138 10220
rect 33818 8652 34138 10164
rect 33818 8596 33846 8652
rect 33902 8596 33950 8652
rect 34006 8596 34054 8652
rect 34110 8596 34138 8652
rect 33818 7084 34138 8596
rect 33818 7028 33846 7084
rect 33902 7028 33950 7084
rect 34006 7028 34054 7084
rect 34110 7028 34138 7084
rect 33818 5516 34138 7028
rect 33818 5460 33846 5516
rect 33902 5460 33950 5516
rect 34006 5460 34054 5516
rect 34110 5460 34138 5516
rect 33818 3948 34138 5460
rect 33818 3892 33846 3948
rect 33902 3892 33950 3948
rect 34006 3892 34054 3948
rect 34110 3892 34138 3948
rect 33818 3076 34138 3892
rect 38480 36092 38800 36908
rect 38480 36036 38508 36092
rect 38564 36036 38612 36092
rect 38668 36036 38716 36092
rect 38772 36036 38800 36092
rect 38480 34524 38800 36036
rect 38480 34468 38508 34524
rect 38564 34468 38612 34524
rect 38668 34468 38716 34524
rect 38772 34468 38800 34524
rect 38480 32956 38800 34468
rect 38480 32900 38508 32956
rect 38564 32900 38612 32956
rect 38668 32900 38716 32956
rect 38772 32900 38800 32956
rect 38480 31388 38800 32900
rect 38480 31332 38508 31388
rect 38564 31332 38612 31388
rect 38668 31332 38716 31388
rect 38772 31332 38800 31388
rect 38480 29820 38800 31332
rect 38480 29764 38508 29820
rect 38564 29764 38612 29820
rect 38668 29764 38716 29820
rect 38772 29764 38800 29820
rect 38480 28252 38800 29764
rect 38480 28196 38508 28252
rect 38564 28196 38612 28252
rect 38668 28196 38716 28252
rect 38772 28196 38800 28252
rect 38480 26684 38800 28196
rect 38480 26628 38508 26684
rect 38564 26628 38612 26684
rect 38668 26628 38716 26684
rect 38772 26628 38800 26684
rect 38480 25116 38800 26628
rect 38480 25060 38508 25116
rect 38564 25060 38612 25116
rect 38668 25060 38716 25116
rect 38772 25060 38800 25116
rect 38480 23548 38800 25060
rect 38480 23492 38508 23548
rect 38564 23492 38612 23548
rect 38668 23492 38716 23548
rect 38772 23492 38800 23548
rect 38480 21980 38800 23492
rect 38480 21924 38508 21980
rect 38564 21924 38612 21980
rect 38668 21924 38716 21980
rect 38772 21924 38800 21980
rect 38480 20412 38800 21924
rect 38480 20356 38508 20412
rect 38564 20356 38612 20412
rect 38668 20356 38716 20412
rect 38772 20356 38800 20412
rect 38480 18844 38800 20356
rect 38480 18788 38508 18844
rect 38564 18788 38612 18844
rect 38668 18788 38716 18844
rect 38772 18788 38800 18844
rect 38480 17276 38800 18788
rect 38480 17220 38508 17276
rect 38564 17220 38612 17276
rect 38668 17220 38716 17276
rect 38772 17220 38800 17276
rect 38480 15708 38800 17220
rect 38480 15652 38508 15708
rect 38564 15652 38612 15708
rect 38668 15652 38716 15708
rect 38772 15652 38800 15708
rect 38480 14140 38800 15652
rect 38480 14084 38508 14140
rect 38564 14084 38612 14140
rect 38668 14084 38716 14140
rect 38772 14084 38800 14140
rect 38480 12572 38800 14084
rect 38480 12516 38508 12572
rect 38564 12516 38612 12572
rect 38668 12516 38716 12572
rect 38772 12516 38800 12572
rect 38480 11004 38800 12516
rect 38480 10948 38508 11004
rect 38564 10948 38612 11004
rect 38668 10948 38716 11004
rect 38772 10948 38800 11004
rect 38480 9436 38800 10948
rect 38480 9380 38508 9436
rect 38564 9380 38612 9436
rect 38668 9380 38716 9436
rect 38772 9380 38800 9436
rect 38480 7868 38800 9380
rect 38480 7812 38508 7868
rect 38564 7812 38612 7868
rect 38668 7812 38716 7868
rect 38772 7812 38800 7868
rect 38480 6300 38800 7812
rect 38480 6244 38508 6300
rect 38564 6244 38612 6300
rect 38668 6244 38716 6300
rect 38772 6244 38800 6300
rect 38480 4732 38800 6244
rect 38480 4676 38508 4732
rect 38564 4676 38612 4732
rect 38668 4676 38716 4732
rect 38772 4676 38800 4732
rect 38480 3164 38800 4676
rect 38480 3108 38508 3164
rect 38564 3108 38612 3164
rect 38668 3108 38716 3164
rect 38772 3108 38800 3164
rect 38480 3076 38800 3108
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _293_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23632 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _294_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _295_
timestamp 1698431365
transform 1 0 22624 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _296_
timestamp 1698431365
transform 1 0 22736 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _297_
timestamp 1698431365
transform 1 0 24080 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _298_
timestamp 1698431365
transform 1 0 25200 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _299_
timestamp 1698431365
transform -1 0 26544 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _300_
timestamp 1698431365
transform 1 0 25312 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _301_
timestamp 1698431365
transform 1 0 24304 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _302_
timestamp 1698431365
transform 1 0 25536 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _303_
timestamp 1698431365
transform -1 0 20496 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _304_
timestamp 1698431365
transform 1 0 21840 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _305_
timestamp 1698431365
transform 1 0 22848 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _306_
timestamp 1698431365
transform 1 0 24080 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _307_
timestamp 1698431365
transform 1 0 21616 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _308_
timestamp 1698431365
transform -1 0 23184 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _309_
timestamp 1698431365
transform 1 0 21728 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _310_
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _311_
timestamp 1698431365
transform 1 0 22736 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _312_
timestamp 1698431365
transform 1 0 23632 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _313_
timestamp 1698431365
transform 1 0 22736 0 1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _314_
timestamp 1698431365
transform 1 0 23968 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _315_
timestamp 1698431365
transform -1 0 21840 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _316_
timestamp 1698431365
transform 1 0 21280 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _317_
timestamp 1698431365
transform 1 0 22176 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _318_
timestamp 1698431365
transform 1 0 20720 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _319_
timestamp 1698431365
transform 1 0 21952 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _320_
timestamp 1698431365
transform 1 0 16016 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _321_
timestamp 1698431365
transform -1 0 17920 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _322_
timestamp 1698431365
transform 1 0 17136 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _323_
timestamp 1698431365
transform 1 0 17360 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _324_
timestamp 1698431365
transform 1 0 17808 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _325_
timestamp 1698431365
transform 1 0 19264 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _326_
timestamp 1698431365
transform -1 0 18592 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _327_
timestamp 1698431365
transform 1 0 17584 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _328_
timestamp 1698431365
transform -1 0 19264 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _329_
timestamp 1698431365
transform 1 0 17584 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _330_
timestamp 1698431365
transform -1 0 19488 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _331_
timestamp 1698431365
transform 1 0 17920 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _332_
timestamp 1698431365
transform 1 0 19376 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _333_
timestamp 1698431365
transform 1 0 17696 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _334_
timestamp 1698431365
transform 1 0 17360 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _335_
timestamp 1698431365
transform 1 0 17920 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _336_
timestamp 1698431365
transform -1 0 19824 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _337_
timestamp 1698431365
transform -1 0 19264 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _338_
timestamp 1698431365
transform 1 0 18256 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _339_
timestamp 1698431365
transform 1 0 19824 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _340_
timestamp 1698431365
transform 1 0 18368 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _341_
timestamp 1698431365
transform 1 0 19712 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _342_
timestamp 1698431365
transform 1 0 18368 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _343_
timestamp 1698431365
transform 1 0 19600 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _344_
timestamp 1698431365
transform 1 0 16464 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _345_
timestamp 1698431365
transform 1 0 15792 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _346_
timestamp 1698431365
transform 1 0 17920 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _347_
timestamp 1698431365
transform 1 0 18928 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _348_
timestamp 1698431365
transform 1 0 16464 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _349_
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _350_
timestamp 1698431365
transform -1 0 17920 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _351_
timestamp 1698431365
transform 1 0 17584 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _352_
timestamp 1698431365
transform -1 0 19488 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _353_
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _354_
timestamp 1698431365
transform -1 0 19152 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _355_
timestamp 1698431365
transform -1 0 17360 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _356_
timestamp 1698431365
transform 1 0 16352 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _357_
timestamp 1698431365
transform 1 0 17360 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _358_
timestamp 1698431365
transform -1 0 19376 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _359_
timestamp 1698431365
transform -1 0 17472 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _360_
timestamp 1698431365
transform 1 0 15792 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _361_
timestamp 1698431365
transform -1 0 19264 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _362_
timestamp 1698431365
transform 1 0 17024 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _363_
timestamp 1698431365
transform -1 0 18592 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _364_
timestamp 1698431365
transform 1 0 17472 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _365_
timestamp 1698431365
transform -1 0 19376 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _366_
timestamp 1698431365
transform 1 0 17136 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _367_
timestamp 1698431365
transform -1 0 19040 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _368_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20720 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _369_
timestamp 1698431365
transform -1 0 28448 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _370_
timestamp 1698431365
transform -1 0 27888 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _371_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24864 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _372_
timestamp 1698431365
transform 1 0 25984 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _373_
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _374_
timestamp 1698431365
transform 1 0 25312 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _375_
timestamp 1698431365
transform 1 0 26432 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _376_
timestamp 1698431365
transform 1 0 27104 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _377_
timestamp 1698431365
transform 1 0 27328 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _378_
timestamp 1698431365
transform 1 0 27776 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _379_
timestamp 1698431365
transform 1 0 28112 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _380_
timestamp 1698431365
transform 1 0 29456 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _381_
timestamp 1698431365
transform 1 0 30128 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _382_
timestamp 1698431365
transform 1 0 31248 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _383_
timestamp 1698431365
transform 1 0 31920 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _384_
timestamp 1698431365
transform 1 0 31920 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _385_
timestamp 1698431365
transform 1 0 31696 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _386_
timestamp 1698431365
transform -1 0 30912 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _387_
timestamp 1698431365
transform 1 0 29680 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _388_
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _389_
timestamp 1698431365
transform 1 0 29456 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _390_
timestamp 1698431365
transform 1 0 30800 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _391_
timestamp 1698431365
transform 1 0 31248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _392_
timestamp 1698431365
transform 1 0 31696 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _393_
timestamp 1698431365
transform 1 0 31136 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _394_
timestamp 1698431365
transform 1 0 32032 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _395_
timestamp 1698431365
transform 1 0 29456 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _396_
timestamp 1698431365
transform 1 0 30352 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _397_
timestamp 1698431365
transform -1 0 25984 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _398_
timestamp 1698431365
transform 1 0 24416 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _399_
timestamp 1698431365
transform 1 0 25312 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _400_
timestamp 1698431365
transform 1 0 24416 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _401_
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _402_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _403_
timestamp 1698431365
transform 1 0 26656 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _404_
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _405_
timestamp 1698431365
transform 1 0 26880 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _406_
timestamp 1698431365
transform 1 0 27776 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _407_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _408_
timestamp 1698431365
transform 1 0 28000 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _409_
timestamp 1698431365
transform 1 0 28896 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _410_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23296 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _411_
timestamp 1698431365
transform 1 0 23072 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _412_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20384 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _413_
timestamp 1698431365
transform 1 0 18704 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _414_
timestamp 1698431365
transform 1 0 24304 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _415_
timestamp 1698431365
transform 1 0 25200 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _416_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26432 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _417_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24080 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _418_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27888 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _419_
timestamp 1698431365
transform 1 0 18704 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _420_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16464 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _421_
timestamp 1698431365
transform -1 0 15344 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _422_
timestamp 1698431365
transform -1 0 26656 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _423_
timestamp 1698431365
transform 1 0 23296 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _424_
timestamp 1698431365
transform 1 0 24416 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _425_
timestamp 1698431365
transform 1 0 22512 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _426_
timestamp 1698431365
transform 1 0 23632 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _427_
timestamp 1698431365
transform -1 0 25984 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _428_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15568 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _429_
timestamp 1698431365
transform 1 0 21952 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _430__1 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _431_
timestamp 1698431365
transform 1 0 22288 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _432_
timestamp 1698431365
transform 1 0 26432 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _433_
timestamp 1698431365
transform 1 0 27552 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _434_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24640 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _435_
timestamp 1698431365
transform 1 0 19376 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _436_
timestamp 1698431365
transform 1 0 20272 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _437_
timestamp 1698431365
transform 1 0 23632 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _438_
timestamp 1698431365
transform 1 0 17248 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _439_
timestamp 1698431365
transform -1 0 18704 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _440_
timestamp 1698431365
transform 1 0 23744 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _441_
timestamp 1698431365
transform 1 0 27440 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _442_
timestamp 1698431365
transform 1 0 28112 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _443_
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _444_
timestamp 1698431365
transform 1 0 19600 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _445_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22064 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _446_
timestamp 1698431365
transform 1 0 18928 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _447_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19824 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _448_
timestamp 1698431365
transform -1 0 24640 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _449_
timestamp 1698431365
transform -1 0 24304 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _450_
timestamp 1698431365
transform 1 0 23520 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _451_
timestamp 1698431365
transform 1 0 23856 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _452_
timestamp 1698431365
transform 1 0 20048 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _453_
timestamp 1698431365
transform 1 0 20832 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _454_
timestamp 1698431365
transform 1 0 21280 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _455_
timestamp 1698431365
transform 1 0 19824 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _456_
timestamp 1698431365
transform 1 0 22624 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _457_
timestamp 1698431365
transform 1 0 23184 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _458_
timestamp 1698431365
transform 1 0 19152 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _459_
timestamp 1698431365
transform -1 0 22624 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _460_
timestamp 1698431365
transform 1 0 21952 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _461_
timestamp 1698431365
transform 1 0 20160 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _462_
timestamp 1698431365
transform 1 0 28896 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _463_
timestamp 1698431365
transform 1 0 30352 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _464_
timestamp 1698431365
transform 1 0 30800 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _465_
timestamp 1698431365
transform 1 0 20832 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _466_
timestamp 1698431365
transform 1 0 32144 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _467_
timestamp 1698431365
transform 1 0 31920 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _468_
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _469_
timestamp 1698431365
transform 1 0 31024 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _470_
timestamp 1698431365
transform 1 0 32816 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _471_
timestamp 1698431365
transform 1 0 21840 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _472_
timestamp 1698431365
transform 1 0 29120 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _473_
timestamp 1698431365
transform 1 0 29680 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _474_
timestamp 1698431365
transform 1 0 23184 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _475_
timestamp 1698431365
transform 1 0 28672 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _476_
timestamp 1698431365
transform -1 0 31248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _477_
timestamp 1698431365
transform 1 0 30128 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _478_
timestamp 1698431365
transform 1 0 23856 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _479_
timestamp 1698431365
transform 1 0 31024 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _480_
timestamp 1698431365
transform 1 0 31920 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _481_
timestamp 1698431365
transform 1 0 23296 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _482_
timestamp 1698431365
transform 1 0 31136 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _483_
timestamp 1698431365
transform 1 0 32032 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _484_
timestamp 1698431365
transform 1 0 23408 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _485_
timestamp 1698431365
transform 1 0 29344 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _486_
timestamp 1698431365
transform 1 0 30240 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _487_
timestamp 1698431365
transform 1 0 22512 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _488_
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _489_
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _490_
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _491_
timestamp 1698431365
transform 1 0 20272 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _492_
timestamp 1698431365
transform 1 0 27664 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _493_
timestamp 1698431365
transform 1 0 28560 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _494_
timestamp 1698431365
transform 1 0 19600 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _495_
timestamp 1698431365
transform 1 0 27440 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _496_
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _497_
timestamp 1698431365
transform 1 0 18928 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _498_
timestamp 1698431365
transform 1 0 26544 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _499_
timestamp 1698431365
transform 1 0 27888 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _500_
timestamp 1698431365
transform 1 0 20272 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _501_
timestamp 1698431365
transform 1 0 24080 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _502_
timestamp 1698431365
transform 1 0 24976 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _503_
timestamp 1698431365
transform 1 0 20048 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _504_
timestamp 1698431365
transform -1 0 25984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _505_
timestamp 1698431365
transform 1 0 24192 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _506_
timestamp 1698431365
transform 1 0 19712 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _507_
timestamp 1698431365
transform 1 0 14560 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _508_
timestamp 1698431365
transform -1 0 15344 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _509_
timestamp 1698431365
transform -1 0 16912 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _510_
timestamp 1698431365
transform -1 0 20272 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _511_
timestamp 1698431365
transform -1 0 17024 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _512_
timestamp 1698431365
transform 1 0 12544 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _513_
timestamp 1698431365
transform -1 0 19824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _514_
timestamp 1698431365
transform -1 0 17248 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _515_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _516_
timestamp 1698431365
transform 1 0 12320 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _517_
timestamp 1698431365
transform 1 0 13216 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _518_
timestamp 1698431365
transform -1 0 15008 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _519_
timestamp 1698431365
transform -1 0 20272 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _520_
timestamp 1698431365
transform -1 0 16128 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _521_
timestamp 1698431365
transform -1 0 14672 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _522_
timestamp 1698431365
transform -1 0 17696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _523_
timestamp 1698431365
transform 1 0 12992 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _524_
timestamp 1698431365
transform -1 0 14112 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _525_
timestamp 1698431365
transform -1 0 16912 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _526_
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _527_
timestamp 1698431365
transform -1 0 14896 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _528_
timestamp 1698431365
transform -1 0 16464 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _529_
timestamp 1698431365
transform 1 0 13104 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _530_
timestamp 1698431365
transform -1 0 14224 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _531_
timestamp 1698431365
transform -1 0 18368 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _532_
timestamp 1698431365
transform 1 0 11312 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _533_
timestamp 1698431365
transform -1 0 12544 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _534_
timestamp 1698431365
transform 1 0 11984 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _535_
timestamp 1698431365
transform -1 0 12768 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _536_
timestamp 1698431365
transform 1 0 11088 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _537_
timestamp 1698431365
transform 1 0 11760 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _538_
timestamp 1698431365
transform -1 0 17024 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _539_
timestamp 1698431365
transform 1 0 11760 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _540_
timestamp 1698431365
transform -1 0 11760 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _541_
timestamp 1698431365
transform -1 0 17584 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _542_
timestamp 1698431365
transform 1 0 11984 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _543_
timestamp 1698431365
transform -1 0 13776 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _544_
timestamp 1698431365
transform -1 0 18032 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _545_
timestamp 1698431365
transform 1 0 11984 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _546_
timestamp 1698431365
transform -1 0 13104 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _547_
timestamp 1698431365
transform -1 0 15568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _548_
timestamp 1698431365
transform 1 0 18256 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _549_
timestamp 1698431365
transform -1 0 14000 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _550_
timestamp 1698431365
transform -1 0 16576 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _551_
timestamp 1698431365
transform 1 0 11312 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _552_
timestamp 1698431365
transform 1 0 12096 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _553_
timestamp 1698431365
transform -1 0 13888 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _554_
timestamp 1698431365
transform 1 0 12432 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _555_
timestamp 1698431365
transform -1 0 16352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _556_
timestamp 1698431365
transform 1 0 11984 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _557_
timestamp 1698431365
transform -1 0 12096 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _558_
timestamp 1698431365
transform -1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _559_
timestamp 1698431365
transform 1 0 12096 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _560_
timestamp 1698431365
transform -1 0 13888 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _561_
timestamp 1698431365
transform -1 0 15792 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _562_
timestamp 1698431365
transform 1 0 11984 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _563_
timestamp 1698431365
transform -1 0 13328 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _564_
timestamp 1698431365
transform -1 0 15904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _565_
timestamp 1698431365
transform -1 0 12432 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _566_
timestamp 1698431365
transform 1 0 12208 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _567_
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _568_
timestamp 1698431365
transform -1 0 13104 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _569_
timestamp 1698431365
transform 1 0 13104 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _570_
timestamp 1698431365
transform -1 0 15904 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _571_
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _572_
timestamp 1698431365
transform -1 0 13104 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _573_
timestamp 1698431365
transform -1 0 16128 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _574_
timestamp 1698431365
transform 1 0 11424 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _575_
timestamp 1698431365
transform -1 0 14000 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _576_
timestamp 1698431365
transform -1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _577_
timestamp 1698431365
transform 1 0 12544 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _578_
timestamp 1698431365
transform -1 0 14336 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _579_
timestamp 1698431365
transform -1 0 18928 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _580_
timestamp 1698431365
transform -1 0 16800 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _581_
timestamp 1698431365
transform -1 0 16800 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _582_
timestamp 1698431365
transform -1 0 14336 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _583_
timestamp 1698431365
transform -1 0 14672 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _584_
timestamp 1698431365
transform 1 0 11200 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _585_
timestamp 1698431365
transform -1 0 18592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _586_
timestamp 1698431365
transform -1 0 14672 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _587_
timestamp 1698431365
transform -1 0 13552 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _588_
timestamp 1698431365
transform -1 0 22288 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _589_
timestamp 1698431365
transform 1 0 21168 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _590_
timestamp 1698431365
transform -1 0 22512 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _591_
timestamp 1698431365
transform -1 0 10976 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _592_
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _593_
timestamp 1698431365
transform -1 0 21840 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _594_
timestamp 1698431365
transform 1 0 9632 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _595_
timestamp 1698431365
transform 1 0 10976 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _596_
timestamp 1698431365
transform -1 0 11984 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _597_
timestamp 1698431365
transform 1 0 11088 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _598_
timestamp 1698431365
transform -1 0 12880 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _599_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11088 0 1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _600_
timestamp 1698431365
transform -1 0 11984 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _601_
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _602_
timestamp 1698431365
transform 1 0 10080 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _603_
timestamp 1698431365
transform -1 0 11088 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _604_
timestamp 1698431365
transform -1 0 9968 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _605_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _606_
timestamp 1698431365
transform 1 0 9184 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _607_
timestamp 1698431365
transform 1 0 9856 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _608_
timestamp 1698431365
transform -1 0 10752 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _609_
timestamp 1698431365
transform 1 0 9744 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _610_
timestamp 1698431365
transform -1 0 10640 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _611_
timestamp 1698431365
transform 1 0 9744 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _612_
timestamp 1698431365
transform -1 0 9744 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _613_
timestamp 1698431365
transform -1 0 11536 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _614_
timestamp 1698431365
transform 1 0 9744 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _615_
timestamp 1698431365
transform -1 0 11536 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _616_
timestamp 1698431365
transform -1 0 21168 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _617_
timestamp 1698431365
transform 1 0 9296 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _618_
timestamp 1698431365
transform -1 0 19936 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _619_
timestamp 1698431365
transform 1 0 8624 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _620_
timestamp 1698431365
transform 1 0 9856 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _621_
timestamp 1698431365
transform -1 0 11424 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _622_
timestamp 1698431365
transform 1 0 9856 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _623_
timestamp 1698431365
transform -1 0 11648 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _624_
timestamp 1698431365
transform 1 0 9632 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _625_
timestamp 1698431365
transform -1 0 8960 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _626_
timestamp 1698431365
transform -1 0 11648 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _627_
timestamp 1698431365
transform 1 0 9968 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _628_
timestamp 1698431365
transform -1 0 10864 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _629_
timestamp 1698431365
transform -1 0 11536 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _630_
timestamp 1698431365
transform 1 0 8736 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _631_
timestamp 1698431365
transform 1 0 10080 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _632_
timestamp 1698431365
transform -1 0 10080 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _633_
timestamp 1698431365
transform 1 0 9968 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _634_
timestamp 1698431365
transform -1 0 10864 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _635_
timestamp 1698431365
transform 1 0 9968 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _636_
timestamp 1698431365
transform -1 0 11536 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _637_
timestamp 1698431365
transform 1 0 10304 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _638_
timestamp 1698431365
transform 1 0 10192 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _639_
timestamp 1698431365
transform -1 0 11984 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _640_
timestamp 1698431365
transform -1 0 23856 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _641_
timestamp 1698431365
transform -1 0 23184 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _642_
timestamp 1698431365
transform 1 0 18592 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _643_
timestamp 1698431365
transform 1 0 19152 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _644_
timestamp 1698431365
transform 1 0 18592 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _645_
timestamp 1698431365
transform -1 0 19712 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _646_
timestamp 1698431365
transform -1 0 16800 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _647_
timestamp 1698431365
transform -1 0 16464 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _648_
timestamp 1698431365
transform -1 0 18256 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _649_
timestamp 1698431365
transform -1 0 16016 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _650_
timestamp 1698431365
transform 1 0 14672 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _651_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15344 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _652_
timestamp 1698431365
transform -1 0 16352 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _653_
timestamp 1698431365
transform -1 0 16240 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _654_
timestamp 1698431365
transform -1 0 15456 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _655_
timestamp 1698431365
transform -1 0 17136 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _656_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _657_
timestamp 1698431365
transform -1 0 15680 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _658_
timestamp 1698431365
transform 1 0 14896 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _659_
timestamp 1698431365
transform -1 0 15792 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _660_
timestamp 1698431365
transform 1 0 14000 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _661_
timestamp 1698431365
transform 1 0 14672 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _662_
timestamp 1698431365
transform 1 0 14336 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _663_
timestamp 1698431365
transform 1 0 14448 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _664_
timestamp 1698431365
transform 1 0 15344 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _665_
timestamp 1698431365
transform 1 0 14448 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _666_
timestamp 1698431365
transform 1 0 15344 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _667_
timestamp 1698431365
transform 1 0 14784 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _668_
timestamp 1698431365
transform 1 0 14448 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _669_
timestamp 1698431365
transform 1 0 14560 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _670_
timestamp 1698431365
transform -1 0 16464 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _671_
timestamp 1698431365
transform -1 0 15680 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _672_
timestamp 1698431365
transform -1 0 15568 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _673_
timestamp 1698431365
transform 1 0 14336 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _674_
timestamp 1698431365
transform -1 0 15120 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _675_
timestamp 1698431365
transform 1 0 20720 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _676_
timestamp 1698431365
transform 1 0 23632 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _677_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19824 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _678_
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _679_
timestamp 1698431365
transform -1 0 26992 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _680_
timestamp 1698431365
transform 1 0 24528 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _681_
timestamp 1698431365
transform 1 0 25648 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _682_
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _683_
timestamp 1698431365
transform 1 0 25760 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _684_
timestamp 1698431365
transform 1 0 26208 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _685_
timestamp 1698431365
transform 1 0 26656 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _686_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _687_
timestamp 1698431365
transform 1 0 27328 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _688_
timestamp 1698431365
transform 1 0 28448 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _689_
timestamp 1698431365
transform 1 0 25872 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _690_
timestamp 1698431365
transform 1 0 25536 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _691_
timestamp 1698431365
transform 1 0 26656 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _692_
timestamp 1698431365
transform 1 0 26208 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _693_
timestamp 1698431365
transform 1 0 27328 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _694_
timestamp 1698431365
transform 1 0 27328 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _695_
timestamp 1698431365
transform 1 0 28448 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _696_
timestamp 1698431365
transform 1 0 26432 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _697_
timestamp 1698431365
transform 1 0 26656 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _698_
timestamp 1698431365
transform 1 0 27552 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _699_
timestamp 1698431365
transform 1 0 26096 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _700_
timestamp 1698431365
transform 1 0 27216 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _701_
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _702_
timestamp 1698431365
transform 1 0 27104 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _703_
timestamp 1698431365
transform 1 0 28112 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _704_
timestamp 1698431365
transform 1 0 26992 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _705_
timestamp 1698431365
transform 1 0 28112 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _706_
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _707_
timestamp 1698431365
transform 1 0 26768 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _708_
timestamp 1698431365
transform 1 0 27888 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _709_
timestamp 1698431365
transform 1 0 25424 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _710_
timestamp 1698431365
transform 1 0 27216 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _711_
timestamp 1698431365
transform 1 0 28336 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _712_
timestamp 1698431365
transform 1 0 27440 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _713_
timestamp 1698431365
transform 1 0 28560 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _714_
timestamp 1698431365
transform 1 0 26320 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _715_
timestamp 1698431365
transform 1 0 27328 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _716_
timestamp 1698431365
transform 1 0 25760 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _717_
timestamp 1698431365
transform 1 0 26096 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _718_
timestamp 1698431365
transform 1 0 26768 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _719_
timestamp 1698431365
transform 1 0 26208 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _720_
timestamp 1698431365
transform 1 0 27104 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _721_
timestamp 1698431365
transform 1 0 26208 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _722_
timestamp 1698431365
transform 1 0 27328 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _723_
timestamp 1698431365
transform 1 0 21056 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _724_
timestamp 1698431365
transform 1 0 21728 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _725_
timestamp 1698431365
transform 1 0 22960 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _726_
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _727_
timestamp 1698431365
transform 1 0 21504 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _728_
timestamp 1698431365
transform 1 0 21616 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _729_
timestamp 1698431365
transform 1 0 23744 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _730_
timestamp 1698431365
transform 1 0 21504 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _731_
timestamp 1698431365
transform 1 0 22848 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _732_
timestamp 1698431365
transform 1 0 21728 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _733_
timestamp 1698431365
transform 1 0 23072 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _734_
timestamp 1698431365
transform -1 0 24080 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _735_
timestamp 1698431365
transform 1 0 22176 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _736_
timestamp 1698431365
transform 1 0 23296 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _737_
timestamp 1698431365
transform 1 0 22512 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _738_
timestamp 1698431365
transform 1 0 21840 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _739_
timestamp 1698431365
transform 1 0 23072 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _740_
timestamp 1698431365
transform 1 0 24192 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _741_
timestamp 1698431365
transform 1 0 23184 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _742_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _743_
timestamp 1698431365
transform 1 0 23184 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _744_
timestamp 1698431365
transform 1 0 24752 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _745_
timestamp 1698431365
transform 1 0 22960 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _746_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18816 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _747_
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _748_
timestamp 1698431365
transform 1 0 18704 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__A2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15792 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__I
timestamp 1698431365
transform -1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__323__I
timestamp 1698431365
transform 1 0 15568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__A2
timestamp 1698431365
transform 1 0 20160 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__A2
timestamp 1698431365
transform 1 0 17360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__329__A2
timestamp 1698431365
transform 1 0 16464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__A2
timestamp 1698431365
transform 1 0 17360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__I
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__I
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__A2
timestamp 1698431365
transform 1 0 16352 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__A2
timestamp 1698431365
transform 1 0 19824 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__A2
timestamp 1698431365
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__A2
timestamp 1698431365
transform 1 0 19488 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__A2
timestamp 1698431365
transform 1 0 19376 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__A2
timestamp 1698431365
transform 1 0 17360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__A2
timestamp 1698431365
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__A2
timestamp 1698431365
transform 1 0 17472 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__A2
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__A2
timestamp 1698431365
transform 1 0 15008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__A2
timestamp 1698431365
transform 1 0 16128 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__A1
timestamp 1698431365
transform 1 0 15344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__I
timestamp 1698431365
transform 1 0 20048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__I
timestamp 1698431365
transform 1 0 19824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__I
timestamp 1698431365
transform 1 0 19600 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__I
timestamp 1698431365
transform 1 0 18368 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__461__I
timestamp 1698431365
transform 1 0 19936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__I
timestamp 1698431365
transform -1 0 20832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__I
timestamp 1698431365
transform 1 0 22736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__I
timestamp 1698431365
transform 1 0 21616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__I
timestamp 1698431365
transform 1 0 21056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__I
timestamp 1698431365
transform -1 0 25312 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__I
timestamp 1698431365
transform 1 0 23632 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__I
timestamp 1698431365
transform 1 0 24192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__487__I
timestamp 1698431365
transform 1 0 22288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__491__I
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__494__I
timestamp 1698431365
transform 1 0 19376 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__I
timestamp 1698431365
transform 1 0 20048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__I
timestamp 1698431365
transform -1 0 16912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__I
timestamp 1698431365
transform 1 0 16912 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__I
timestamp 1698431365
transform 1 0 15792 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__I
timestamp 1698431365
transform 1 0 15344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__I
timestamp 1698431365
transform -1 0 17920 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__538__I
timestamp 1698431365
transform 1 0 15904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__I
timestamp 1698431365
transform -1 0 17696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__544__I
timestamp 1698431365
transform 1 0 16352 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__547__I
timestamp 1698431365
transform 1 0 14336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__549__I
timestamp 1698431365
transform 1 0 14000 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__I
timestamp 1698431365
transform 1 0 11984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__555__I
timestamp 1698431365
transform -1 0 14336 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__558__I
timestamp 1698431365
transform 1 0 16016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__561__I
timestamp 1698431365
transform 1 0 14448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__I
timestamp 1698431365
transform 1 0 14560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__565__I
timestamp 1698431365
transform 1 0 12432 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__566__I
timestamp 1698431365
transform -1 0 13328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__570__I
timestamp 1698431365
transform -1 0 14448 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__573__I
timestamp 1698431365
transform 1 0 15456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__579__I
timestamp 1698431365
transform 1 0 17248 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__617__I
timestamp 1698431365
transform 1 0 9968 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__619__I
timestamp 1698431365
transform -1 0 8624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__629__I
timestamp 1698431365
transform -1 0 11760 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__630__I
timestamp 1698431365
transform 1 0 8512 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__638__A1
timestamp 1698431365
transform -1 0 11536 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__642__A1
timestamp 1698431365
transform 1 0 18256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__644__A1
timestamp 1698431365
transform 1 0 19376 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__726__I
timestamp 1698431365
transform -1 0 21392 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__727__I
timestamp 1698431365
transform 1 0 22400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__737__I
timestamp 1698431365
transform 1 0 22848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__738__I
timestamp 1698431365
transform 1 0 20496 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform 1 0 27104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 3136 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 5488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 8064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 10416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 15904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 6944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 15232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 6384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 6944 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 4480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 5488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 2464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 2464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 34720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 15904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 21616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 22288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 20384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output23_I
timestamp 1698431365
transform 1 0 33824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output31_I
timestamp 1698431365
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output32_I
timestamp 1698431365
transform 1 0 37520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output33_I
timestamp 1698431365
transform 1 0 36400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output38_I
timestamp 1698431365
transform -1 0 37744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output41_I
timestamp 1698431365
transform 1 0 35728 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output47_I
timestamp 1698431365
transform 1 0 34160 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output52_I
timestamp 1698431365
transform 1 0 6384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output58_I
timestamp 1698431365
transform 1 0 7616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output65_I
timestamp 1698431365
transform 1 0 36848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output78_I
timestamp 1698431365
transform 1 0 38080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output82_I
timestamp 1698431365
transform 1 0 37520 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output85_I
timestamp 1698431365
transform 1 0 3584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output89_I
timestamp 1698431365
transform -1 0 2688 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output91_I
timestamp 1698431365
transform -1 0 2688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output92_I
timestamp 1698431365
transform 1 0 2912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output94_I
timestamp 1698431365
transform 1 0 3136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output95_I
timestamp 1698431365
transform -1 0 2464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output108_I
timestamp 1698431365
transform 1 0 35280 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output112_I
timestamp 1698431365
transform 1 0 2464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output122_I
timestamp 1698431365
transform 1 0 36288 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output124_I
timestamp 1698431365
transform -1 0 4256 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output129_I
timestamp 1698431365
transform -1 0 3360 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output141_I
timestamp 1698431365
transform 1 0 37520 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output142_I
timestamp 1698431365
transform 1 0 2464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output153_I
timestamp 1698431365
transform -1 0 37744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output154_I
timestamp 1698431365
transform 1 0 37520 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output163_I
timestamp 1698431365
transform 1 0 37520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output165_I
timestamp 1698431365
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output166_I
timestamp 1698431365
transform 1 0 33712 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output168_I
timestamp 1698431365
transform 1 0 37520 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output170_I
timestamp 1698431365
transform -1 0 37744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output171_I
timestamp 1698431365
transform -1 0 37744 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output177_I
timestamp 1698431365
transform 1 0 32480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output181_I
timestamp 1698431365
transform 1 0 10416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0__276_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk
timestamp 1698431365
transform -1 0 27104 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f__276_
timestamp 1698431365
transform -1 0 24864 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698431365
transform -1 0 24080 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f__276_
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout183
timestamp 1698431365
transform -1 0 20944 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout184
timestamp 1698431365
transform 1 0 18256 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_36 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_199 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698431365
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_270
timestamp 1698431365
transform 1 0 31584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_304
timestamp 1698431365
transform 1 0 35392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_308 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_316
timestamp 1698431365
transform 1 0 36736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_320
timestamp 1698431365
transform 1 0 37184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_322
timestamp 1698431365
transform 1 0 37408 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_34
timestamp 1698431365
transform 1 0 5152 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_43
timestamp 1698431365
transform 1 0 6160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_47
timestamp 1698431365
transform 1 0 6608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_49
timestamp 1698431365
transform 1 0 6832 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_52
timestamp 1698431365
transform 1 0 7168 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_58
timestamp 1698431365
transform 1 0 7840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_62
timestamp 1698431365
transform 1 0 8288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_79
timestamp 1698431365
transform 1 0 10192 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_83
timestamp 1698431365
transform 1 0 10640 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_115
timestamp 1698431365
transform 1 0 14224 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_123
timestamp 1698431365
transform 1 0 15120 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_127
timestamp 1698431365
transform 1 0 15568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_129
timestamp 1698431365
transform 1 0 15792 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_132
timestamp 1698431365
transform 1 0 16128 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_158
timestamp 1698431365
transform 1 0 19040 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_166
timestamp 1698431365
transform 1 0 19936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_172
timestamp 1698431365
transform 1 0 20608 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_176
timestamp 1698431365
transform 1 0 21056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_178
timestamp 1698431365
transform 1 0 21280 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_181
timestamp 1698431365
transform 1 0 21616 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_187
timestamp 1698431365
transform 1 0 22288 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698431365
transform 1 0 24080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698431365
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_228
timestamp 1698431365
transform 1 0 26880 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_235
timestamp 1698431365
transform 1 0 27664 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_267
timestamp 1698431365
transform 1 0 31248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_275
timestamp 1698431365
transform 1 0 32144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_292
timestamp 1698431365
transform 1 0 34048 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_298
timestamp 1698431365
transform 1 0 34720 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_314
timestamp 1698431365
transform 1 0 36512 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_322
timestamp 1698431365
transform 1 0 37408 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_321
timestamp 1698431365
transform 1 0 37296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_314
timestamp 1698431365
transform 1 0 36512 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_322
timestamp 1698431365
transform 1 0 37408 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_321
timestamp 1698431365
transform 1 0 37296 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_6
timestamp 1698431365
transform 1 0 2016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_10
timestamp 1698431365
transform 1 0 2464 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_42
timestamp 1698431365
transform 1 0 6048 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_58
timestamp 1698431365
transform 1 0 7840 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_150
timestamp 1698431365
transform 1 0 18144 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_154
timestamp 1698431365
transform 1 0 18592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_184
timestamp 1698431365
transform 1 0 21952 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_188
timestamp 1698431365
transform 1 0 22400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_190
timestamp 1698431365
transform 1 0 22624 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_195
timestamp 1698431365
transform 1 0 23184 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_200
timestamp 1698431365
transform 1 0 23744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_314
timestamp 1698431365
transform 1 0 36512 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_322
timestamp 1698431365
transform 1 0 37408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_324
timestamp 1698431365
transform 1 0 37632 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_14
timestamp 1698431365
transform 1 0 2912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_18
timestamp 1698431365
transform 1 0 3360 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_181
timestamp 1698431365
transform 1 0 21616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_183
timestamp 1698431365
transform 1 0 21840 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_196
timestamp 1698431365
transform 1 0 23296 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_198
timestamp 1698431365
transform 1 0 23520 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_221
timestamp 1698431365
transform 1 0 26096 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_229
timestamp 1698431365
transform 1 0 26992 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_232
timestamp 1698431365
transform 1 0 27328 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_240
timestamp 1698431365
transform 1 0 28224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_8
timestamp 1698431365
transform 1 0 2240 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_40
timestamp 1698431365
transform 1 0 5824 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_56
timestamp 1698431365
transform 1 0 7616 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_64
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_68
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_150
timestamp 1698431365
transform 1 0 18144 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_154
timestamp 1698431365
transform 1 0 18592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_185
timestamp 1698431365
transform 1 0 22064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_262
timestamp 1698431365
transform 1 0 30688 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_278
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_314
timestamp 1698431365
transform 1 0 36512 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_322
timestamp 1698431365
transform 1 0 37408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_324
timestamp 1698431365
transform 1 0 37632 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_8
timestamp 1698431365
transform 1 0 2240 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_24
timestamp 1698431365
transform 1 0 4032 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698431365
transform 1 0 4928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_139
timestamp 1698431365
transform 1 0 16912 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_155
timestamp 1698431365
transform 1 0 18704 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_159
timestamp 1698431365
transform 1 0 19152 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_163
timestamp 1698431365
transform 1 0 19600 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_167
timestamp 1698431365
transform 1 0 20048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_169
timestamp 1698431365
transform 1 0 20272 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_179
timestamp 1698431365
transform 1 0 21392 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_243
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_297
timestamp 1698431365
transform 1 0 34608 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_313
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_8
timestamp 1698431365
transform 1 0 2240 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_40
timestamp 1698431365
transform 1 0 5824 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_56
timestamp 1698431365
transform 1 0 7616 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_64
timestamp 1698431365
transform 1 0 8512 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_68
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_146
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_262
timestamp 1698431365
transform 1 0 30688 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_278
timestamp 1698431365
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_314
timestamp 1698431365
transform 1 0 36512 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_322
timestamp 1698431365
transform 1 0 37408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_324
timestamp 1698431365
transform 1 0 37632 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_8
timestamp 1698431365
transform 1 0 2240 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_24
timestamp 1698431365
transform 1 0 4032 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1698431365
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_69
timestamp 1698431365
transform 1 0 9072 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_77
timestamp 1698431365
transform 1 0 9968 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_91
timestamp 1698431365
transform 1 0 11536 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_99
timestamp 1698431365
transform 1 0 12432 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_103
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_113
timestamp 1698431365
transform 1 0 14000 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_121
timestamp 1698431365
transform 1 0 14896 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_124
timestamp 1698431365
transform 1 0 15232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_128
timestamp 1698431365
transform 1 0 15680 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_224
timestamp 1698431365
transform 1 0 26432 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_253
timestamp 1698431365
transform 1 0 29680 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_285
timestamp 1698431365
transform 1 0 33264 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_301
timestamp 1698431365
transform 1 0 35056 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_309
timestamp 1698431365
transform 1 0 35952 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_313
timestamp 1698431365
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_8
timestamp 1698431365
transform 1 0 2240 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_40
timestamp 1698431365
transform 1 0 5824 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_56
timestamp 1698431365
transform 1 0 7616 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_64
timestamp 1698431365
transform 1 0 8512 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_68
timestamp 1698431365
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_76
timestamp 1698431365
transform 1 0 9856 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_87
timestamp 1698431365
transform 1 0 11088 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_89
timestamp 1698431365
transform 1 0 11312 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_116
timestamp 1698431365
transform 1 0 14336 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_150
timestamp 1698431365
transform 1 0 18144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_152
timestamp 1698431365
transform 1 0 18368 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698431365
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_234
timestamp 1698431365
transform 1 0 27552 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_249
timestamp 1698431365
transform 1 0 29232 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_265
timestamp 1698431365
transform 1 0 31024 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_273
timestamp 1698431365
transform 1 0 31920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_277
timestamp 1698431365
transform 1 0 32368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_314
timestamp 1698431365
transform 1 0 36512 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_322
timestamp 1698431365
transform 1 0 37408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_324
timestamp 1698431365
transform 1 0 37632 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_14
timestamp 1698431365
transform 1 0 2912 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_30
timestamp 1698431365
transform 1 0 4704 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_69
timestamp 1698431365
transform 1 0 9072 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_87
timestamp 1698431365
transform 1 0 11088 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_91
timestamp 1698431365
transform 1 0 11536 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_117
timestamp 1698431365
transform 1 0 14448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_135
timestamp 1698431365
transform 1 0 16464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_154
timestamp 1698431365
transform 1 0 18592 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_161
timestamp 1698431365
transform 1 0 19376 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_181
timestamp 1698431365
transform 1 0 21616 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_205
timestamp 1698431365
transform 1 0 24304 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_238
timestamp 1698431365
transform 1 0 28000 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698431365
transform 1 0 28448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_8
timestamp 1698431365
transform 1 0 2240 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_40
timestamp 1698431365
transform 1 0 5824 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_56
timestamp 1698431365
transform 1 0 7616 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_64
timestamp 1698431365
transform 1 0 8512 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_68
timestamp 1698431365
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_76
timestamp 1698431365
transform 1 0 9856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_78
timestamp 1698431365
transform 1 0 10080 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_95
timestamp 1698431365
transform 1 0 11984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_103
timestamp 1698431365
transform 1 0 12880 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_107
timestamp 1698431365
transform 1 0 13328 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_123
timestamp 1698431365
transform 1 0 15120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_125
timestamp 1698431365
transform 1 0 15344 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_130
timestamp 1698431365
transform 1 0 15904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_218
timestamp 1698431365
transform 1 0 25760 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_222
timestamp 1698431365
transform 1 0 26208 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_249
timestamp 1698431365
transform 1 0 29232 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_265
timestamp 1698431365
transform 1 0 31024 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_273
timestamp 1698431365
transform 1 0 31920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698431365
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_314
timestamp 1698431365
transform 1 0 36512 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_322
timestamp 1698431365
transform 1 0 37408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_324
timestamp 1698431365
transform 1 0 37632 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_8
timestamp 1698431365
transform 1 0 2240 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_24
timestamp 1698431365
transform 1 0 4032 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_32
timestamp 1698431365
transform 1 0 4928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_53
timestamp 1698431365
transform 1 0 7280 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_61
timestamp 1698431365
transform 1 0 8176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_63
timestamp 1698431365
transform 1 0 8400 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_88
timestamp 1698431365
transform 1 0 11200 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_90
timestamp 1698431365
transform 1 0 11424 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_117
timestamp 1698431365
transform 1 0 14448 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_142
timestamp 1698431365
transform 1 0 17248 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_185
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_189
timestamp 1698431365
transform 1 0 22512 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_202
timestamp 1698431365
transform 1 0 23968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_220
timestamp 1698431365
transform 1 0 25984 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_224
timestamp 1698431365
transform 1 0 26432 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_226
timestamp 1698431365
transform 1 0 26656 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_233
timestamp 1698431365
transform 1 0 27440 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_237
timestamp 1698431365
transform 1 0 27888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_261
timestamp 1698431365
transform 1 0 30576 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_293
timestamp 1698431365
transform 1 0 34160 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_309
timestamp 1698431365
transform 1 0 35952 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_313
timestamp 1698431365
transform 1 0 36400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_8
timestamp 1698431365
transform 1 0 2240 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_40
timestamp 1698431365
transform 1 0 5824 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_56
timestamp 1698431365
transform 1 0 7616 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_64
timestamp 1698431365
transform 1 0 8512 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1698431365
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_76
timestamp 1698431365
transform 1 0 9856 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_91
timestamp 1698431365
transform 1 0 11536 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_97
timestamp 1698431365
transform 1 0 12208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_107
timestamp 1698431365
transform 1 0 13328 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_111
timestamp 1698431365
transform 1 0 13776 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_115
timestamp 1698431365
transform 1 0 14224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_117
timestamp 1698431365
transform 1 0 14448 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_126
timestamp 1698431365
transform 1 0 15456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_130
timestamp 1698431365
transform 1 0 15904 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_133
timestamp 1698431365
transform 1 0 16240 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_159
timestamp 1698431365
transform 1 0 19152 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_166
timestamp 1698431365
transform 1 0 19936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_170
timestamp 1698431365
transform 1 0 20384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_172
timestamp 1698431365
transform 1 0 20608 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_183
timestamp 1698431365
transform 1 0 21840 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_195
timestamp 1698431365
transform 1 0 23184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_214
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_247
timestamp 1698431365
transform 1 0 29008 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698431365
transform 1 0 36512 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_322
timestamp 1698431365
transform 1 0 37408 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_324
timestamp 1698431365
transform 1 0 37632 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_8
timestamp 1698431365
transform 1 0 2240 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_24
timestamp 1698431365
transform 1 0 4032 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698431365
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_53
timestamp 1698431365
transform 1 0 7280 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_61
timestamp 1698431365
transform 1 0 8176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_87
timestamp 1698431365
transform 1 0 11088 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_113
timestamp 1698431365
transform 1 0 14000 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_141
timestamp 1698431365
transform 1 0 17136 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_162
timestamp 1698431365
transform 1 0 19488 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_169
timestamp 1698431365
transform 1 0 20272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698431365
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_187
timestamp 1698431365
transform 1 0 22288 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_191
timestamp 1698431365
transform 1 0 22736 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_203
timestamp 1698431365
transform 1 0 24080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_222
timestamp 1698431365
transform 1 0 26208 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_238
timestamp 1698431365
transform 1 0 28000 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698431365
transform 1 0 28448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_265
timestamp 1698431365
transform 1 0 31024 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_280
timestamp 1698431365
transform 1 0 32704 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_8
timestamp 1698431365
transform 1 0 2240 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_40
timestamp 1698431365
transform 1 0 5824 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_56
timestamp 1698431365
transform 1 0 7616 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_64
timestamp 1698431365
transform 1 0 8512 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698431365
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_86
timestamp 1698431365
transform 1 0 10976 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_94
timestamp 1698431365
transform 1 0 11872 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_112
timestamp 1698431365
transform 1 0 13888 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_116
timestamp 1698431365
transform 1 0 14336 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698431365
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698431365
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_153
timestamp 1698431365
transform 1 0 18480 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_163
timestamp 1698431365
transform 1 0 19600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_189
timestamp 1698431365
transform 1 0 22512 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_197
timestamp 1698431365
transform 1 0 23408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_201
timestamp 1698431365
transform 1 0 23856 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_219
timestamp 1698431365
transform 1 0 25872 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_243
timestamp 1698431365
transform 1 0 28560 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_264
timestamp 1698431365
transform 1 0 30912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698431365
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_322
timestamp 1698431365
transform 1 0 37408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_324
timestamp 1698431365
transform 1 0 37632 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_14
timestamp 1698431365
transform 1 0 2912 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_30
timestamp 1698431365
transform 1 0 4704 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_53
timestamp 1698431365
transform 1 0 7280 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_61
timestamp 1698431365
transform 1 0 8176 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_68
timestamp 1698431365
transform 1 0 8960 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_92
timestamp 1698431365
transform 1 0 11648 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_94
timestamp 1698431365
transform 1 0 11872 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_115
timestamp 1698431365
transform 1 0 14224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_133
timestamp 1698431365
transform 1 0 16240 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_141
timestamp 1698431365
transform 1 0 17136 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_159
timestamp 1698431365
transform 1 0 19152 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_169
timestamp 1698431365
transform 1 0 20272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698431365
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_187
timestamp 1698431365
transform 1 0 22288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_189
timestamp 1698431365
transform 1 0 22512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_202
timestamp 1698431365
transform 1 0 23968 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_225
timestamp 1698431365
transform 1 0 26544 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_253
timestamp 1698431365
transform 1 0 29680 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_261
timestamp 1698431365
transform 1 0 30576 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_279
timestamp 1698431365
transform 1 0 32592 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_8
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_40
timestamp 1698431365
transform 1 0 5824 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_56
timestamp 1698431365
transform 1 0 7616 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_64
timestamp 1698431365
transform 1 0 8512 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_112
timestamp 1698431365
transform 1 0 13888 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_122
timestamp 1698431365
transform 1 0 15008 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_127
timestamp 1698431365
transform 1 0 15568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_129
timestamp 1698431365
transform 1 0 15792 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_134
timestamp 1698431365
transform 1 0 16352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_146
timestamp 1698431365
transform 1 0 17696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_160
timestamp 1698431365
transform 1 0 19264 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_170
timestamp 1698431365
transform 1 0 20384 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_174
timestamp 1698431365
transform 1 0 20832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_226
timestamp 1698431365
transform 1 0 26656 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_240
timestamp 1698431365
transform 1 0 28224 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_248
timestamp 1698431365
transform 1 0 29120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_250
timestamp 1698431365
transform 1 0 29344 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_275
timestamp 1698431365
transform 1 0 32144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698431365
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_322
timestamp 1698431365
transform 1 0 37408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_324
timestamp 1698431365
transform 1 0 37632 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_8
timestamp 1698431365
transform 1 0 2240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_12
timestamp 1698431365
transform 1 0 2688 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698431365
transform 1 0 4480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698431365
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_69
timestamp 1698431365
transform 1 0 9072 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_77
timestamp 1698431365
transform 1 0 9968 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_79
timestamp 1698431365
transform 1 0 10192 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_92
timestamp 1698431365
transform 1 0 11648 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_96
timestamp 1698431365
transform 1 0 12096 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_98
timestamp 1698431365
transform 1 0 12320 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_115
timestamp 1698431365
transform 1 0 14224 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_124
timestamp 1698431365
transform 1 0 15232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_144
timestamp 1698431365
transform 1 0 17472 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_169
timestamp 1698431365
transform 1 0 20272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_183
timestamp 1698431365
transform 1 0 21840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_185
timestamp 1698431365
transform 1 0 22064 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_192
timestamp 1698431365
transform 1 0 22848 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_210
timestamp 1698431365
transform 1 0 24864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_214
timestamp 1698431365
transform 1 0 25312 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_230
timestamp 1698431365
transform 1 0 27104 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_253
timestamp 1698431365
transform 1 0 29680 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_269
timestamp 1698431365
transform 1 0 31472 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_277
timestamp 1698431365
transform 1 0 32368 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_309
timestamp 1698431365
transform 1 0 35952 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_313
timestamp 1698431365
transform 1 0 36400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_8
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_12
timestamp 1698431365
transform 1 0 2688 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_44
timestamp 1698431365
transform 1 0 6272 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698431365
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698431365
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_84
timestamp 1698431365
transform 1 0 10752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_86
timestamp 1698431365
transform 1 0 10976 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_111
timestamp 1698431365
transform 1 0 13776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_119
timestamp 1698431365
transform 1 0 14672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_129
timestamp 1698431365
transform 1 0 15792 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_133
timestamp 1698431365
transform 1 0 16240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_149
timestamp 1698431365
transform 1 0 18032 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_151
timestamp 1698431365
transform 1 0 18256 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_163
timestamp 1698431365
transform 1 0 19600 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_167
timestamp 1698431365
transform 1 0 20048 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_179
timestamp 1698431365
transform 1 0 21392 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_218
timestamp 1698431365
transform 1 0 25760 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_236
timestamp 1698431365
transform 1 0 27776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_238
timestamp 1698431365
transform 1 0 28000 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_245
timestamp 1698431365
transform 1 0 28784 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_259
timestamp 1698431365
transform 1 0 30352 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_267
timestamp 1698431365
transform 1 0 31248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698431365
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698431365
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_322
timestamp 1698431365
transform 1 0 37408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_324
timestamp 1698431365
transform 1 0 37632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_8
timestamp 1698431365
transform 1 0 2240 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_24
timestamp 1698431365
transform 1 0 4032 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698431365
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698431365
transform 1 0 9072 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698431365
transform 1 0 9520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_91
timestamp 1698431365
transform 1 0 11536 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_149
timestamp 1698431365
transform 1 0 18032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_162
timestamp 1698431365
transform 1 0 19488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_170
timestamp 1698431365
transform 1 0 20384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_189
timestamp 1698431365
transform 1 0 22512 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_193
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_206
timestamp 1698431365
transform 1 0 24416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_208
timestamp 1698431365
transform 1 0 24640 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_215
timestamp 1698431365
transform 1 0 25424 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_225
timestamp 1698431365
transform 1 0 26544 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_233
timestamp 1698431365
transform 1 0 27440 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_240
timestamp 1698431365
transform 1 0 28224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_264
timestamp 1698431365
transform 1 0 30912 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_287
timestamp 1698431365
transform 1 0 33488 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_303
timestamp 1698431365
transform 1 0 35280 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_8
timestamp 1698431365
transform 1 0 2240 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_40
timestamp 1698431365
transform 1 0 5824 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_56
timestamp 1698431365
transform 1 0 7616 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_64
timestamp 1698431365
transform 1 0 8512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_74
timestamp 1698431365
transform 1 0 9632 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_91
timestamp 1698431365
transform 1 0 11536 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_111
timestamp 1698431365
transform 1 0 13776 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_119
timestamp 1698431365
transform 1 0 14672 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_128
timestamp 1698431365
transform 1 0 15680 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_132
timestamp 1698431365
transform 1 0 16128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_171
timestamp 1698431365
transform 1 0 20496 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_173
timestamp 1698431365
transform 1 0 20720 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_186
timestamp 1698431365
transform 1 0 22176 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_190
timestamp 1698431365
transform 1 0 22624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_205
timestamp 1698431365
transform 1 0 24304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_218
timestamp 1698431365
transform 1 0 25760 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_248
timestamp 1698431365
transform 1 0 29120 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_252
timestamp 1698431365
transform 1 0 29568 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_259
timestamp 1698431365
transform 1 0 30352 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_267
timestamp 1698431365
transform 1 0 31248 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_271
timestamp 1698431365
transform 1 0 31696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698431365
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_322
timestamp 1698431365
transform 1 0 37408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_324
timestamp 1698431365
transform 1 0 37632 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_14
timestamp 1698431365
transform 1 0 2912 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_30
timestamp 1698431365
transform 1 0 4704 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_85
timestamp 1698431365
transform 1 0 10864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_103
timestamp 1698431365
transform 1 0 12880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_111
timestamp 1698431365
transform 1 0 13776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_131
timestamp 1698431365
transform 1 0 16016 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_138
timestamp 1698431365
transform 1 0 16800 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_144
timestamp 1698431365
transform 1 0 17472 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_148
timestamp 1698431365
transform 1 0 17920 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_150
timestamp 1698431365
transform 1 0 18144 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_157
timestamp 1698431365
transform 1 0 18928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_165
timestamp 1698431365
transform 1 0 19824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_185
timestamp 1698431365
transform 1 0 22064 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_203
timestamp 1698431365
transform 1 0 24080 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_210
timestamp 1698431365
transform 1 0 24864 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_214
timestamp 1698431365
transform 1 0 25312 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_238
timestamp 1698431365
transform 1 0 28000 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_283
timestamp 1698431365
transform 1 0 33040 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_8
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_40
timestamp 1698431365
transform 1 0 5824 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_56
timestamp 1698431365
transform 1 0 7616 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_64
timestamp 1698431365
transform 1 0 8512 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698431365
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_76
timestamp 1698431365
transform 1 0 9856 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_83
timestamp 1698431365
transform 1 0 10640 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_91
timestamp 1698431365
transform 1 0 11536 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_95
timestamp 1698431365
transform 1 0 11984 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_102
timestamp 1698431365
transform 1 0 12768 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_130
timestamp 1698431365
transform 1 0 15904 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_152
timestamp 1698431365
transform 1 0 18368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_164
timestamp 1698431365
transform 1 0 19712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_174
timestamp 1698431365
transform 1 0 20832 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_176
timestamp 1698431365
transform 1 0 21056 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_179
timestamp 1698431365
transform 1 0 21392 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_195
timestamp 1698431365
transform 1 0 23184 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_208
timestamp 1698431365
transform 1 0 24640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_226
timestamp 1698431365
transform 1 0 26656 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_242
timestamp 1698431365
transform 1 0 28448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_252
timestamp 1698431365
transform 1 0 29568 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_256
timestamp 1698431365
transform 1 0 30016 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_269
timestamp 1698431365
transform 1 0 31472 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698431365
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_322
timestamp 1698431365
transform 1 0 37408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_324
timestamp 1698431365
transform 1 0 37632 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_8
timestamp 1698431365
transform 1 0 2240 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_24
timestamp 1698431365
transform 1 0 4032 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_69
timestamp 1698431365
transform 1 0 9072 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_86
timestamp 1698431365
transform 1 0 10976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_88
timestamp 1698431365
transform 1 0 11200 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_123
timestamp 1698431365
transform 1 0 15120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_127
timestamp 1698431365
transform 1 0 15568 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_131
timestamp 1698431365
transform 1 0 16016 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_138
timestamp 1698431365
transform 1 0 16800 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_140
timestamp 1698431365
transform 1 0 17024 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_164
timestamp 1698431365
transform 1 0 19712 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698431365
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_201
timestamp 1698431365
transform 1 0 23856 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_217
timestamp 1698431365
transform 1 0 25648 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_221
timestamp 1698431365
transform 1 0 26096 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_232
timestamp 1698431365
transform 1 0 27328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_253
timestamp 1698431365
transform 1 0 29680 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_285
timestamp 1698431365
transform 1 0 33264 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_301
timestamp 1698431365
transform 1 0 35056 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_309
timestamp 1698431365
transform 1 0 35952 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_313
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_8
timestamp 1698431365
transform 1 0 2240 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_40
timestamp 1698431365
transform 1 0 5824 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_56
timestamp 1698431365
transform 1 0 7616 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_64
timestamp 1698431365
transform 1 0 8512 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_84
timestamp 1698431365
transform 1 0 10752 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_100
timestamp 1698431365
transform 1 0 12544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_102
timestamp 1698431365
transform 1 0 12768 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_135
timestamp 1698431365
transform 1 0 16464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_148
timestamp 1698431365
transform 1 0 17920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_164
timestamp 1698431365
transform 1 0 19712 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_166
timestamp 1698431365
transform 1 0 19936 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_190
timestamp 1698431365
transform 1 0 22624 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_198
timestamp 1698431365
transform 1 0 23520 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_202
timestamp 1698431365
transform 1 0 23968 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_220
timestamp 1698431365
transform 1 0 25984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_252
timestamp 1698431365
transform 1 0 29568 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_268
timestamp 1698431365
transform 1 0 31360 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698431365
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_322
timestamp 1698431365
transform 1 0 37408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_324
timestamp 1698431365
transform 1 0 37632 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_8
timestamp 1698431365
transform 1 0 2240 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_24
timestamp 1698431365
transform 1 0 4032 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_69
timestamp 1698431365
transform 1 0 9072 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_85
timestamp 1698431365
transform 1 0 10864 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_95
timestamp 1698431365
transform 1 0 11984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_97
timestamp 1698431365
transform 1 0 12208 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_115
timestamp 1698431365
transform 1 0 14224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_127
timestamp 1698431365
transform 1 0 15568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_153
timestamp 1698431365
transform 1 0 18480 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_159
timestamp 1698431365
transform 1 0 19152 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_163
timestamp 1698431365
transform 1 0 19600 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_183
timestamp 1698431365
transform 1 0 21840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_187
timestamp 1698431365
transform 1 0 22288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_219
timestamp 1698431365
transform 1 0 25872 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_223
timestamp 1698431365
transform 1 0 26320 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_240
timestamp 1698431365
transform 1 0 28224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698431365
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_8
timestamp 1698431365
transform 1 0 2240 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_40
timestamp 1698431365
transform 1 0 5824 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_56
timestamp 1698431365
transform 1 0 7616 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_64
timestamp 1698431365
transform 1 0 8512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_96
timestamp 1698431365
transform 1 0 12096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_122
timestamp 1698431365
transform 1 0 15008 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_126
timestamp 1698431365
transform 1 0 15456 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698431365
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_172
timestamp 1698431365
transform 1 0 20608 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_205
timestamp 1698431365
transform 1 0 24304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_220
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_222
timestamp 1698431365
transform 1 0 26208 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_229
timestamp 1698431365
transform 1 0 26992 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_241
timestamp 1698431365
transform 1 0 28336 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698431365
transform 1 0 31920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698431365
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698431365
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_322
timestamp 1698431365
transform 1 0 37408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_324
timestamp 1698431365
transform 1 0 37632 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_14
timestamp 1698431365
transform 1 0 2912 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_30
timestamp 1698431365
transform 1 0 4704 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_69
timestamp 1698431365
transform 1 0 9072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_114
timestamp 1698431365
transform 1 0 14112 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_118
timestamp 1698431365
transform 1 0 14560 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_139
timestamp 1698431365
transform 1 0 16912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_158
timestamp 1698431365
transform 1 0 19040 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_166
timestamp 1698431365
transform 1 0 19936 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_170
timestamp 1698431365
transform 1 0 20384 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_198
timestamp 1698431365
transform 1 0 23520 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_206
timestamp 1698431365
transform 1 0 24416 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_223
timestamp 1698431365
transform 1 0 26320 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_225
timestamp 1698431365
transform 1 0 26544 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_232
timestamp 1698431365
transform 1 0 27328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_236
timestamp 1698431365
transform 1 0 27776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_238
timestamp 1698431365
transform 1 0 28000 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_8
timestamp 1698431365
transform 1 0 2240 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_40
timestamp 1698431365
transform 1 0 5824 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_56
timestamp 1698431365
transform 1 0 7616 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_64
timestamp 1698431365
transform 1 0 8512 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698431365
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_80
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_84
timestamp 1698431365
transform 1 0 10752 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_86
timestamp 1698431365
transform 1 0 10976 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_103
timestamp 1698431365
transform 1 0 12880 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_114
timestamp 1698431365
transform 1 0 14112 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_134
timestamp 1698431365
transform 1 0 16352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_146
timestamp 1698431365
transform 1 0 17696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_159
timestamp 1698431365
transform 1 0 19152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_173
timestamp 1698431365
transform 1 0 20720 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_181
timestamp 1698431365
transform 1 0 21616 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_193
timestamp 1698431365
transform 1 0 22960 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_248
timestamp 1698431365
transform 1 0 29120 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_314
timestamp 1698431365
transform 1 0 36512 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_322
timestamp 1698431365
transform 1 0 37408 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_8
timestamp 1698431365
transform 1 0 2240 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_24
timestamp 1698431365
transform 1 0 4032 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_32
timestamp 1698431365
transform 1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_69
timestamp 1698431365
transform 1 0 9072 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_85
timestamp 1698431365
transform 1 0 10864 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_95
timestamp 1698431365
transform 1 0 11984 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_103
timestamp 1698431365
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_117
timestamp 1698431365
transform 1 0 14448 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_133
timestamp 1698431365
transform 1 0 16240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_137
timestamp 1698431365
transform 1 0 16688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_141
timestamp 1698431365
transform 1 0 17136 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_162
timestamp 1698431365
transform 1 0 19488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_164
timestamp 1698431365
transform 1 0 19712 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_167
timestamp 1698431365
transform 1 0 20048 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_179
timestamp 1698431365
transform 1 0 21392 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_191
timestamp 1698431365
transform 1 0 22736 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_205
timestamp 1698431365
transform 1 0 24304 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_209
timestamp 1698431365
transform 1 0 24752 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_224
timestamp 1698431365
transform 1 0 26432 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_228
timestamp 1698431365
transform 1 0 26880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_230
timestamp 1698431365
transform 1 0 27104 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_237
timestamp 1698431365
transform 1 0 27888 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_8
timestamp 1698431365
transform 1 0 2240 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_12
timestamp 1698431365
transform 1 0 2688 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_44
timestamp 1698431365
transform 1 0 6272 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_60
timestamp 1698431365
transform 1 0 8064 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698431365
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_104
timestamp 1698431365
transform 1 0 12992 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_121
timestamp 1698431365
transform 1 0 14896 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_127
timestamp 1698431365
transform 1 0 15568 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698431365
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_144
timestamp 1698431365
transform 1 0 17472 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_156
timestamp 1698431365
transform 1 0 18816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_158
timestamp 1698431365
transform 1 0 19040 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_171
timestamp 1698431365
transform 1 0 20496 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_173
timestamp 1698431365
transform 1 0 20720 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_240
timestamp 1698431365
transform 1 0 28224 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_272
timestamp 1698431365
transform 1 0 31808 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_314
timestamp 1698431365
transform 1 0 36512 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_322
timestamp 1698431365
transform 1 0 37408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_324
timestamp 1698431365
transform 1 0 37632 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_8
timestamp 1698431365
transform 1 0 2240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_12
timestamp 1698431365
transform 1 0 2688 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_28
timestamp 1698431365
transform 1 0 4480 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_32
timestamp 1698431365
transform 1 0 4928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_115
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_131
timestamp 1698431365
transform 1 0 16016 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_139
timestamp 1698431365
transform 1 0 16912 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_145
timestamp 1698431365
transform 1 0 17584 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_149
timestamp 1698431365
transform 1 0 18032 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_151
timestamp 1698431365
transform 1 0 18256 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_160
timestamp 1698431365
transform 1 0 19264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_162
timestamp 1698431365
transform 1 0 19488 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_165
timestamp 1698431365
transform 1 0 19824 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_173
timestamp 1698431365
transform 1 0 20720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_190
timestamp 1698431365
transform 1 0 22624 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_194
timestamp 1698431365
transform 1 0 23072 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_207
timestamp 1698431365
transform 1 0 24528 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_211
timestamp 1698431365
transform 1 0 24976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_213
timestamp 1698431365
transform 1 0 25200 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_226
timestamp 1698431365
transform 1 0 26656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_242
timestamp 1698431365
transform 1 0 28448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_8
timestamp 1698431365
transform 1 0 2240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_12
timestamp 1698431365
transform 1 0 2688 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_44
timestamp 1698431365
transform 1 0 6272 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_60
timestamp 1698431365
transform 1 0 8064 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_68
timestamp 1698431365
transform 1 0 8960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_314
timestamp 1698431365
transform 1 0 36512 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_322
timestamp 1698431365
transform 1 0 37408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_324
timestamp 1698431365
transform 1 0 37632 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_14
timestamp 1698431365
transform 1 0 2912 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_18
timestamp 1698431365
transform 1 0 3360 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_8
timestamp 1698431365
transform 1 0 2240 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_12
timestamp 1698431365
transform 1 0 2688 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_16
timestamp 1698431365
transform 1 0 3136 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_48
timestamp 1698431365
transform 1 0 6720 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_64
timestamp 1698431365
transform 1 0 8512 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_68
timestamp 1698431365
transform 1 0 8960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_314
timestamp 1698431365
transform 1 0 36512 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_322
timestamp 1698431365
transform 1 0 37408 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_8
timestamp 1698431365
transform 1 0 2240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_12
timestamp 1698431365
transform 1 0 2688 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_28
timestamp 1698431365
transform 1 0 4480 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_32
timestamp 1698431365
transform 1 0 4928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_321
timestamp 1698431365
transform 1 0 37296 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_314
timestamp 1698431365
transform 1 0 36512 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_322
timestamp 1698431365
transform 1 0 37408 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_321
timestamp 1698431365
transform 1 0 37296 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_10
timestamp 1698431365
transform 1 0 2464 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_14
timestamp 1698431365
transform 1 0 2912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_18
timestamp 1698431365
transform 1 0 3360 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_22
timestamp 1698431365
transform 1 0 3808 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_26
timestamp 1698431365
transform 1 0 4256 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_30
timestamp 1698431365
transform 1 0 4704 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_34
timestamp 1698431365
transform 1 0 5152 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_43
timestamp 1698431365
transform 1 0 6160 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_47
timestamp 1698431365
transform 1 0 6608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_49
timestamp 1698431365
transform 1 0 6832 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_52
timestamp 1698431365
transform 1 0 7168 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_79
timestamp 1698431365
transform 1 0 10192 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_83
timestamp 1698431365
transform 1 0 10640 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_115
timestamp 1698431365
transform 1 0 14224 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_123
timestamp 1698431365
transform 1 0 15120 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_126
timestamp 1698431365
transform 1 0 15456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_132
timestamp 1698431365
transform 1 0 16128 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_228
timestamp 1698431365
transform 1 0 26880 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_235
timestamp 1698431365
transform 1 0 27664 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_267
timestamp 1698431365
transform 1 0 31248 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_275
timestamp 1698431365
transform 1 0 32144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_277
timestamp 1698431365
transform 1 0 32368 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_286
timestamp 1698431365
transform 1 0 33376 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_288
timestamp 1698431365
transform 1 0 33600 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_291
timestamp 1698431365
transform 1 0 33936 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_301
timestamp 1698431365
transform 1 0 35056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_305
timestamp 1698431365
transform 1 0 35504 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_309
timestamp 1698431365
transform 1 0 35952 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_311
timestamp 1698431365
transform 1 0 36176 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_314
timestamp 1698431365
transform 1 0 36512 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_316
timestamp 1698431365
transform 1 0 36736 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_36
timestamp 1698431365
transform 1 0 5376 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_70
timestamp 1698431365
transform 1 0 9184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_138
timestamp 1698431365
transform 1 0 16800 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_172
timestamp 1698431365
transform 1 0 20608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_199
timestamp 1698431365
transform 1 0 23632 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_203
timestamp 1698431365
transform 1 0 24080 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_236
timestamp 1698431365
transform 1 0 27776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_270
timestamp 1698431365
transform 1 0 31584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_304
timestamp 1698431365
transform 1 0 35392 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_326
timestamp 1698431365
transform 1 0 37856 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_330
timestamp 1698431365
transform 1 0 38304 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698431365
transform 1 0 2464 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input2
timestamp 1698431365
transform 1 0 5488 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input3
timestamp 1698431365
transform 1 0 7616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform 1 0 9408 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 9520 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 8288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 15232 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input8
timestamp 1698431365
transform 1 0 6272 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 14560 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 5600 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 6272 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 3808 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input13
timestamp 1698431365
transform 1 0 9520 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input14
timestamp 1698431365
transform 1 0 5488 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input15
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input16
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input17
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input18
timestamp 1698431365
transform -1 0 35392 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 15232 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform -1 0 22288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 22960 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  net99_2
timestamp 1698431365
transform -1 0 24864 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  net99_3
timestamp 1698431365
transform -1 0 26096 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  net99_4
timestamp 1698431365
transform -1 0 23184 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output23
timestamp 1698431365
transform -1 0 34720 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output24
timestamp 1698431365
transform -1 0 34048 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output25
timestamp 1698431365
transform -1 0 30240 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output26
timestamp 1698431365
transform -1 0 32704 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output27
timestamp 1698431365
transform -1 0 23632 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output28
timestamp 1698431365
transform -1 0 30912 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output29
timestamp 1698431365
transform -1 0 26432 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output30
timestamp 1698431365
transform -1 0 27776 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output31
timestamp 1698431365
transform -1 0 37856 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output32
timestamp 1698431365
transform 1 0 37744 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output33
timestamp 1698431365
transform 1 0 37072 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output34
timestamp 1698431365
transform 1 0 37744 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output35
timestamp 1698431365
transform -1 0 25088 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output36
timestamp 1698431365
transform -1 0 27104 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output37
timestamp 1698431365
transform -1 0 25760 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output38
timestamp 1698431365
transform 1 0 37744 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output39
timestamp 1698431365
transform -1 0 23632 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output40
timestamp 1698431365
transform -1 0 16912 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output41
timestamp 1698431365
transform -1 0 36512 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output42
timestamp 1698431365
transform 1 0 37744 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output43
timestamp 1698431365
transform 1 0 17696 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output44
timestamp 1698431365
transform 1 0 17024 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output45
timestamp 1698431365
transform 1 0 19712 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output46
timestamp 1698431365
transform 1 0 18368 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output47
timestamp 1698431365
transform -1 0 35056 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output48
timestamp 1698431365
transform -1 0 21616 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output49
timestamp 1698431365
transform -1 0 21616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output50
timestamp 1698431365
transform 1 0 19040 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output51
timestamp 1698431365
transform 1 0 15904 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output52
timestamp 1698431365
transform 1 0 5600 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output53
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output54
timestamp 1698431365
transform 1 0 17696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output55
timestamp 1698431365
transform 1 0 18368 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output56
timestamp 1698431365
transform -1 0 16912 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output57
timestamp 1698431365
transform 1 0 17024 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output58
timestamp 1698431365
transform 1 0 6944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output59
timestamp 1698431365
transform 1 0 15904 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output60
timestamp 1698431365
transform -1 0 32704 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output61
timestamp 1698431365
transform -1 0 27664 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output62
timestamp 1698431365
transform -1 0 30912 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output63
timestamp 1698431365
transform -1 0 30240 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output64
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output65
timestamp 1698431365
transform 1 0 37072 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output66
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output67
timestamp 1698431365
transform 1 0 37744 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output68
timestamp 1698431365
transform 1 0 37744 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output69
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output70
timestamp 1698431365
transform 1 0 37744 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output71
timestamp 1698431365
transform 1 0 37744 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output72
timestamp 1698431365
transform 1 0 37744 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output73
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output74
timestamp 1698431365
transform -1 0 31584 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output75
timestamp 1698431365
transform 1 0 37072 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output76
timestamp 1698431365
transform -1 0 33376 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output77
timestamp 1698431365
transform -1 0 27664 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output78
timestamp 1698431365
transform 1 0 37744 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output79
timestamp 1698431365
transform 1 0 37072 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output80
timestamp 1698431365
transform -1 0 29568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output81
timestamp 1698431365
transform -1 0 28896 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output82
timestamp 1698431365
transform 1 0 37744 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output83
timestamp 1698431365
transform 1 0 37744 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output84
timestamp 1698431365
transform 1 0 6944 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output85
timestamp 1698431365
transform -1 0 3808 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output86
timestamp 1698431365
transform -1 0 22960 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output87
timestamp 1698431365
transform 1 0 10080 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output88
timestamp 1698431365
transform 1 0 11424 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output89
timestamp 1698431365
transform -1 0 2240 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output90
timestamp 1698431365
transform -1 0 2240 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output91
timestamp 1698431365
transform -1 0 2240 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output92
timestamp 1698431365
transform -1 0 2240 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output93
timestamp 1698431365
transform -1 0 2240 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output94
timestamp 1698431365
transform -1 0 2912 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output95
timestamp 1698431365
transform -1 0 2240 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output96
timestamp 1698431365
transform -1 0 2240 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output97
timestamp 1698431365
transform -1 0 25760 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output98
timestamp 1698431365
transform -1 0 2240 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output99
timestamp 1698431365
transform 1 0 10752 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output100
timestamp 1698431365
transform 1 0 12096 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output101
timestamp 1698431365
transform 1 0 11424 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output102
timestamp 1698431365
transform -1 0 2912 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output103
timestamp 1698431365
transform -1 0 2240 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output104
timestamp 1698431365
transform -1 0 2240 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output105
timestamp 1698431365
transform -1 0 2240 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output106
timestamp 1698431365
transform 1 0 10752 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output107
timestamp 1698431365
transform -1 0 2240 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output108
timestamp 1698431365
transform -1 0 35392 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output109
timestamp 1698431365
transform -1 0 2240 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output110
timestamp 1698431365
transform -1 0 2240 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output111
timestamp 1698431365
transform -1 0 2240 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output112
timestamp 1698431365
transform -1 0 2240 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output113
timestamp 1698431365
transform -1 0 2240 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output114
timestamp 1698431365
transform -1 0 2240 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output115
timestamp 1698431365
transform -1 0 2240 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output116
timestamp 1698431365
transform -1 0 2240 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output117
timestamp 1698431365
transform -1 0 2240 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output118
timestamp 1698431365
transform -1 0 2240 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output119
timestamp 1698431365
transform 1 0 37744 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output120
timestamp 1698431365
transform -1 0 2240 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output121
timestamp 1698431365
transform -1 0 2240 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output122
timestamp 1698431365
transform -1 0 37184 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output123
timestamp 1698431365
transform 1 0 19040 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output124
timestamp 1698431365
transform -1 0 5152 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output125
timestamp 1698431365
transform 1 0 8288 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output126
timestamp 1698431365
transform -1 0 14560 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output127
timestamp 1698431365
transform 1 0 7616 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output128
timestamp 1698431365
transform -1 0 2912 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output129
timestamp 1698431365
transform -1 0 2912 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output130
timestamp 1698431365
transform 1 0 37744 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output131
timestamp 1698431365
transform -1 0 2240 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output132
timestamp 1698431365
transform -1 0 2240 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output133
timestamp 1698431365
transform -1 0 2240 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output134
timestamp 1698431365
transform -1 0 2912 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output135
timestamp 1698431365
transform -1 0 2240 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output136
timestamp 1698431365
transform -1 0 2912 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output137
timestamp 1698431365
transform -1 0 15232 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output138
timestamp 1698431365
transform -1 0 13888 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output139
timestamp 1698431365
transform 1 0 10080 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output140
timestamp 1698431365
transform -1 0 14560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output141
timestamp 1698431365
transform 1 0 37744 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output142
timestamp 1698431365
transform -1 0 2240 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output143
timestamp 1698431365
transform -1 0 2240 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output144
timestamp 1698431365
transform -1 0 27776 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output145
timestamp 1698431365
transform -1 0 27104 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output146
timestamp 1698431365
transform -1 0 28896 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output147
timestamp 1698431365
transform -1 0 29568 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output148
timestamp 1698431365
transform 1 0 37072 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output149
timestamp 1698431365
transform 1 0 37744 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output150
timestamp 1698431365
transform 1 0 37744 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output151
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output152
timestamp 1698431365
transform 1 0 37072 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output153
timestamp 1698431365
transform 1 0 37744 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output154
timestamp 1698431365
transform 1 0 37744 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output155
timestamp 1698431365
transform 1 0 37072 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output156
timestamp 1698431365
transform 1 0 37744 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output157
timestamp 1698431365
transform 1 0 37744 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output158
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output159
timestamp 1698431365
transform 1 0 37744 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output160
timestamp 1698431365
transform 1 0 37744 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output161
timestamp 1698431365
transform 1 0 37744 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output162
timestamp 1698431365
transform 1 0 37744 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output163
timestamp 1698431365
transform 1 0 37744 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output164
timestamp 1698431365
transform -1 0 25088 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output165
timestamp 1698431365
transform -1 0 34048 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output166
timestamp 1698431365
transform -1 0 34720 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output167
timestamp 1698431365
transform -1 0 26432 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output168
timestamp 1698431365
transform 1 0 37744 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output169
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output170
timestamp 1698431365
transform 1 0 37744 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output171
timestamp 1698431365
transform 1 0 37744 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output172
timestamp 1698431365
transform 1 0 37744 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output173
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output174
timestamp 1698431365
transform 1 0 37744 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output175
timestamp 1698431365
transform -1 0 31584 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output176
timestamp 1698431365
transform 1 0 12096 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output177
timestamp 1698431365
transform -1 0 33376 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output178
timestamp 1698431365
transform -1 0 13888 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output179
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output180
timestamp 1698431365
transform -1 0 22288 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output181
timestamp 1698431365
transform 1 0 9408 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  output182
timestamp 1698431365
transform 1 0 37744 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_43 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_44
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 38640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_45
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 38640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_46
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_47
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_48
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 38640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_49
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 38640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_50
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 38640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_51
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_52
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 38640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_53
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 38640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 38640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 38640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 38640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 38640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 38640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 38640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 38640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 38640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 38640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 38640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 38640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 38640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 38640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 38640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 38640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 38640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 38640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 38640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 38640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_86 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_87
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_88
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_89
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_95
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_96
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_97
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_98
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_99
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_100
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_101
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_102
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_103
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_104
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_105
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_106
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_107
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_108
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_109
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_110
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_111
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_112
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_113
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_114
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_115
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_116
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_117
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_118
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_119
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_120
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_121
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_122
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_123
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_124
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_125
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_126
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_127
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_128
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_129
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_130
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_131
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_132
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_133
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_134
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_135
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_136
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_137
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_138
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_139
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_140
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_141
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_142
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_143
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_144
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_145
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_146
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_147
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_148
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_149
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_150
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_151
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_152
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_153
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_154
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_155
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_156
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_157
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_158
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_159
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_160
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_161
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_162
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_163
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_164
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_165
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_166
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_167
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_168
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_169
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_170
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_171
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_172
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_173
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_174
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_175
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_176
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_177
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_178
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_179
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_180
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_181
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_182
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_183
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_184
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_185
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_186
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_187
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_188
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_189
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_190
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_191
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_192
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_193
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_194
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_195
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_196
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_197
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_198
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_199
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_200
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_201
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_202
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_203
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_204
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_205
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_206
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_207
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_208
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_209
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_210
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_211
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_212
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_213
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_214
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_215
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_216
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_217
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_218
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_219
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_220
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_221
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_222
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_223
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_224
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_225
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_226
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_227
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_228
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_229
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_230
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_231
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_232
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_233
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_234
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_235
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_236
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_237
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_238
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_239
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_240
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_241
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_242
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_243
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_244
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_245
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_246
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_247
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_248
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_249
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_250
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_251
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_252
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_253
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_254
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_255
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_256
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_257
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_258
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_259
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_260
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_261
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_262
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_263
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_264
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_265
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_266
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_267
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_268
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_269
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_270
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_271
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_272
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_273
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_274
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_275
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_276
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_277
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_278
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_279
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_280
timestamp 1698431365
transform 1 0 8960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_281
timestamp 1698431365
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_282
timestamp 1698431365
transform 1 0 16576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_283
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698431365
transform 1 0 24192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698431365
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698431365
transform 1 0 31808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 310 870
<< labels >>
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 2688 39200 2800 40000 0 FreeSans 448 90 0 0 in[0]
port 1 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 in[10]
port 2 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 in[11]
port 3 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 in[12]
port 4 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 in[13]
port 5 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 in[14]
port 6 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 in[15]
port 7 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 in[16]
port 8 nsew signal input
flabel metal2 s 14784 39200 14896 40000 0 FreeSans 448 90 0 0 in[17]
port 9 nsew signal input
flabel metal2 s 6048 39200 6160 40000 0 FreeSans 448 90 0 0 in[1]
port 10 nsew signal input
flabel metal2 s 6720 39200 6832 40000 0 FreeSans 448 90 0 0 in[2]
port 11 nsew signal input
flabel metal2 s 4032 39200 4144 40000 0 FreeSans 448 90 0 0 in[3]
port 12 nsew signal input
flabel metal2 s 9408 39200 9520 40000 0 FreeSans 448 90 0 0 in[4]
port 13 nsew signal input
flabel metal2 s 5376 39200 5488 40000 0 FreeSans 448 90 0 0 in[5]
port 14 nsew signal input
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 in[6]
port 15 nsew signal input
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 in[7]
port 16 nsew signal input
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 in[8]
port 17 nsew signal input
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 in[9]
port 18 nsew signal input
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 proj_clk[0]
port 19 nsew signal tristate
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 proj_clk[1]
port 20 nsew signal tristate
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 proj_clk[2]
port 21 nsew signal tristate
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 proj_clk[3]
port 22 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 proj_clk[4]
port 23 nsew signal tristate
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 proj_clk[5]
port 24 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 proj_clk[6]
port 25 nsew signal tristate
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 proj_clk[7]
port 26 nsew signal tristate
flabel metal2 s 36288 39200 36400 40000 0 FreeSans 448 90 0 0 proj_in[0]
port 27 nsew signal tristate
flabel metal3 s 39200 3360 40000 3472 0 FreeSans 448 0 0 0 proj_in[100]
port 28 nsew signal tristate
flabel metal3 s 39200 7392 40000 7504 0 FreeSans 448 0 0 0 proj_in[101]
port 29 nsew signal tristate
flabel metal3 s 39200 15456 40000 15568 0 FreeSans 448 0 0 0 proj_in[102]
port 30 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 proj_in[103]
port 31 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 proj_in[104]
port 32 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 proj_in[105]
port 33 nsew signal tristate
flabel metal3 s 39200 5376 40000 5488 0 FreeSans 448 0 0 0 proj_in[106]
port 34 nsew signal tristate
flabel metal2 s 22848 39200 22960 40000 0 FreeSans 448 90 0 0 proj_in[107]
port 35 nsew signal tristate
flabel metal2 s 16128 39200 16240 40000 0 FreeSans 448 90 0 0 proj_in[108]
port 36 nsew signal tristate
flabel metal2 s 34944 39200 35056 40000 0 FreeSans 448 90 0 0 proj_in[109]
port 37 nsew signal tristate
flabel metal3 s 39200 8064 40000 8176 0 FreeSans 448 0 0 0 proj_in[10]
port 38 nsew signal tristate
flabel metal2 s 18144 39200 18256 40000 0 FreeSans 448 90 0 0 proj_in[110]
port 39 nsew signal tristate
flabel metal2 s 17472 39200 17584 40000 0 FreeSans 448 90 0 0 proj_in[111]
port 40 nsew signal tristate
flabel metal2 s 20160 39200 20272 40000 0 FreeSans 448 90 0 0 proj_in[112]
port 41 nsew signal tristate
flabel metal2 s 18816 39200 18928 40000 0 FreeSans 448 90 0 0 proj_in[113]
port 42 nsew signal tristate
flabel metal2 s 34272 39200 34384 40000 0 FreeSans 448 90 0 0 proj_in[114]
port 43 nsew signal tristate
flabel metal2 s 20832 39200 20944 40000 0 FreeSans 448 90 0 0 proj_in[115]
port 44 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 proj_in[116]
port 45 nsew signal tristate
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 proj_in[117]
port 46 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 proj_in[118]
port 47 nsew signal tristate
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 proj_in[119]
port 48 nsew signal tristate
flabel metal3 s 39200 9408 40000 9520 0 FreeSans 448 0 0 0 proj_in[11]
port 49 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 proj_in[120]
port 50 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 proj_in[121]
port 51 nsew signal tristate
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 proj_in[122]
port 52 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 proj_in[123]
port 53 nsew signal tristate
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 proj_in[124]
port 54 nsew signal tristate
flabel metal2 s 16800 39200 16912 40000 0 FreeSans 448 90 0 0 proj_in[125]
port 55 nsew signal tristate
flabel metal2 s 30912 39200 31024 40000 0 FreeSans 448 90 0 0 proj_in[126]
port 56 nsew signal tristate
flabel metal2 s 26880 39200 26992 40000 0 FreeSans 448 90 0 0 proj_in[127]
port 57 nsew signal tristate
flabel metal2 s 29568 39200 29680 40000 0 FreeSans 448 90 0 0 proj_in[128]
port 58 nsew signal tristate
flabel metal2 s 28896 39200 29008 40000 0 FreeSans 448 90 0 0 proj_in[129]
port 59 nsew signal tristate
flabel metal3 s 39200 10752 40000 10864 0 FreeSans 448 0 0 0 proj_in[12]
port 60 nsew signal tristate
flabel metal3 s 39200 35616 40000 35728 0 FreeSans 448 0 0 0 proj_in[130]
port 61 nsew signal tristate
flabel metal3 s 39200 29568 40000 29680 0 FreeSans 448 0 0 0 proj_in[131]
port 62 nsew signal tristate
flabel metal3 s 39200 24864 40000 24976 0 FreeSans 448 0 0 0 proj_in[132]
port 63 nsew signal tristate
flabel metal3 s 39200 20832 40000 20944 0 FreeSans 448 0 0 0 proj_in[133]
port 64 nsew signal tristate
flabel metal3 s 39200 18816 40000 18928 0 FreeSans 448 0 0 0 proj_in[134]
port 65 nsew signal tristate
flabel metal3 s 39200 6720 40000 6832 0 FreeSans 448 0 0 0 proj_in[135]
port 66 nsew signal tristate
flabel metal3 s 39200 8736 40000 8848 0 FreeSans 448 0 0 0 proj_in[136]
port 67 nsew signal tristate
flabel metal3 s 39200 16128 40000 16240 0 FreeSans 448 0 0 0 proj_in[137]
port 68 nsew signal tristate
flabel metal3 s 39200 14112 40000 14224 0 FreeSans 448 0 0 0 proj_in[138]
port 69 nsew signal tristate
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 proj_in[139]
port 70 nsew signal tristate
flabel metal3 s 39200 12096 40000 12208 0 FreeSans 448 0 0 0 proj_in[13]
port 71 nsew signal tristate
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 proj_in[140]
port 72 nsew signal tristate
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 proj_in[141]
port 73 nsew signal tristate
flabel metal3 s 39200 34944 40000 35056 0 FreeSans 448 0 0 0 proj_in[142]
port 74 nsew signal tristate
flabel metal3 s 39200 31584 40000 31696 0 FreeSans 448 0 0 0 proj_in[143]
port 75 nsew signal tristate
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 proj_in[14]
port 76 nsew signal tristate
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 proj_in[15]
port 77 nsew signal tristate
flabel metal3 s 39200 32256 40000 32368 0 FreeSans 448 0 0 0 proj_in[16]
port 78 nsew signal tristate
flabel metal3 s 39200 26208 40000 26320 0 FreeSans 448 0 0 0 proj_in[17]
port 79 nsew signal tristate
flabel metal2 s 7392 39200 7504 40000 0 FreeSans 448 90 0 0 proj_in[18]
port 80 nsew signal tristate
flabel metal2 s 3360 39200 3472 40000 0 FreeSans 448 90 0 0 proj_in[19]
port 81 nsew signal tristate
flabel metal2 s 22176 39200 22288 40000 0 FreeSans 448 90 0 0 proj_in[1]
port 82 nsew signal tristate
flabel metal2 s 10752 39200 10864 40000 0 FreeSans 448 90 0 0 proj_in[20]
port 83 nsew signal tristate
flabel metal2 s 12096 39200 12208 40000 0 FreeSans 448 90 0 0 proj_in[21]
port 84 nsew signal tristate
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 proj_in[22]
port 85 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 proj_in[23]
port 86 nsew signal tristate
flabel metal3 s 0 29568 800 29680 0 FreeSans 448 0 0 0 proj_in[24]
port 87 nsew signal tristate
flabel metal3 s 0 32256 800 32368 0 FreeSans 448 0 0 0 proj_in[25]
port 88 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 proj_in[26]
port 89 nsew signal tristate
flabel metal3 s 0 7392 800 7504 0 FreeSans 448 0 0 0 proj_in[27]
port 90 nsew signal tristate
flabel metal3 s 0 8064 800 8176 0 FreeSans 448 0 0 0 proj_in[28]
port 91 nsew signal tristate
flabel metal3 s 0 10752 800 10864 0 FreeSans 448 0 0 0 proj_in[29]
port 92 nsew signal tristate
flabel metal2 s 24192 39200 24304 40000 0 FreeSans 448 90 0 0 proj_in[2]
port 93 nsew signal tristate
flabel metal3 s 0 14112 800 14224 0 FreeSans 448 0 0 0 proj_in[30]
port 94 nsew signal tristate
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 proj_in[31]
port 95 nsew signal tristate
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 proj_in[32]
port 96 nsew signal tristate
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 proj_in[33]
port 97 nsew signal tristate
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 proj_in[34]
port 98 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 proj_in[35]
port 99 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 proj_in[36]
port 100 nsew signal tristate
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 proj_in[37]
port 101 nsew signal tristate
flabel metal2 s 11424 39200 11536 40000 0 FreeSans 448 90 0 0 proj_in[38]
port 102 nsew signal tristate
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 proj_in[39]
port 103 nsew signal tristate
flabel metal2 s 33600 39200 33712 40000 0 FreeSans 448 90 0 0 proj_in[3]
port 104 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 proj_in[40]
port 105 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 proj_in[41]
port 106 nsew signal tristate
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 proj_in[42]
port 107 nsew signal tristate
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 proj_in[43]
port 108 nsew signal tristate
flabel metal3 s 0 11424 800 11536 0 FreeSans 448 0 0 0 proj_in[44]
port 109 nsew signal tristate
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 proj_in[45]
port 110 nsew signal tristate
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 proj_in[46]
port 111 nsew signal tristate
flabel metal3 s 0 9408 800 9520 0 FreeSans 448 0 0 0 proj_in[47]
port 112 nsew signal tristate
flabel metal3 s 0 12768 800 12880 0 FreeSans 448 0 0 0 proj_in[48]
port 113 nsew signal tristate
flabel metal3 s 0 8736 800 8848 0 FreeSans 448 0 0 0 proj_in[49]
port 114 nsew signal tristate
flabel metal3 s 39200 24192 40000 24304 0 FreeSans 448 0 0 0 proj_in[4]
port 115 nsew signal tristate
flabel metal3 s 0 10080 800 10192 0 FreeSans 448 0 0 0 proj_in[50]
port 116 nsew signal tristate
flabel metal3 s 0 13440 800 13552 0 FreeSans 448 0 0 0 proj_in[51]
port 117 nsew signal tristate
flabel metal2 s 35616 39200 35728 40000 0 FreeSans 448 90 0 0 proj_in[52]
port 118 nsew signal tristate
flabel metal2 s 19488 39200 19600 40000 0 FreeSans 448 90 0 0 proj_in[53]
port 119 nsew signal tristate
flabel metal2 s 4704 39200 4816 40000 0 FreeSans 448 90 0 0 proj_in[54]
port 120 nsew signal tristate
flabel metal2 s 8736 39200 8848 40000 0 FreeSans 448 90 0 0 proj_in[55]
port 121 nsew signal tristate
flabel metal2 s 14112 39200 14224 40000 0 FreeSans 448 90 0 0 proj_in[56]
port 122 nsew signal tristate
flabel metal2 s 8064 39200 8176 40000 0 FreeSans 448 90 0 0 proj_in[57]
port 123 nsew signal tristate
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 proj_in[58]
port 124 nsew signal tristate
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 proj_in[59]
port 125 nsew signal tristate
flabel metal3 s 39200 30912 40000 31024 0 FreeSans 448 0 0 0 proj_in[5]
port 126 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 proj_in[60]
port 127 nsew signal tristate
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 proj_in[61]
port 128 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 proj_in[62]
port 129 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 proj_in[63]
port 130 nsew signal tristate
flabel metal3 s 0 14784 800 14896 0 FreeSans 448 0 0 0 proj_in[64]
port 131 nsew signal tristate
flabel metal3 s 0 12096 800 12208 0 FreeSans 448 0 0 0 proj_in[65]
port 132 nsew signal tristate
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 proj_in[66]
port 133 nsew signal tristate
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 proj_in[67]
port 134 nsew signal tristate
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 proj_in[68]
port 135 nsew signal tristate
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 proj_in[69]
port 136 nsew signal tristate
flabel metal3 s 39200 33600 40000 33712 0 FreeSans 448 0 0 0 proj_in[6]
port 137 nsew signal tristate
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 proj_in[70]
port 138 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 proj_in[71]
port 139 nsew signal tristate
flabel metal2 s 26208 39200 26320 40000 0 FreeSans 448 90 0 0 proj_in[72]
port 140 nsew signal tristate
flabel metal2 s 25536 39200 25648 40000 0 FreeSans 448 90 0 0 proj_in[73]
port 141 nsew signal tristate
flabel metal2 s 27552 39200 27664 40000 0 FreeSans 448 90 0 0 proj_in[74]
port 142 nsew signal tristate
flabel metal2 s 28224 39200 28336 40000 0 FreeSans 448 90 0 0 proj_in[75]
port 143 nsew signal tristate
flabel metal3 s 39200 26880 40000 26992 0 FreeSans 448 0 0 0 proj_in[76]
port 144 nsew signal tristate
flabel metal3 s 39200 22848 40000 22960 0 FreeSans 448 0 0 0 proj_in[77]
port 145 nsew signal tristate
flabel metal3 s 39200 22176 40000 22288 0 FreeSans 448 0 0 0 proj_in[78]
port 146 nsew signal tristate
flabel metal3 s 39200 20160 40000 20272 0 FreeSans 448 0 0 0 proj_in[79]
port 147 nsew signal tristate
flabel metal3 s 39200 21504 40000 21616 0 FreeSans 448 0 0 0 proj_in[7]
port 148 nsew signal tristate
flabel metal3 s 39200 4032 40000 4144 0 FreeSans 448 0 0 0 proj_in[80]
port 149 nsew signal tristate
flabel metal3 s 39200 6048 40000 6160 0 FreeSans 448 0 0 0 proj_in[81]
port 150 nsew signal tristate
flabel metal3 s 39200 16800 40000 16912 0 FreeSans 448 0 0 0 proj_in[82]
port 151 nsew signal tristate
flabel metal3 s 39200 10080 40000 10192 0 FreeSans 448 0 0 0 proj_in[83]
port 152 nsew signal tristate
flabel metal3 s 39200 14784 40000 14896 0 FreeSans 448 0 0 0 proj_in[84]
port 153 nsew signal tristate
flabel metal3 s 39200 12768 40000 12880 0 FreeSans 448 0 0 0 proj_in[85]
port 154 nsew signal tristate
flabel metal3 s 39200 13440 40000 13552 0 FreeSans 448 0 0 0 proj_in[86]
port 155 nsew signal tristate
flabel metal3 s 39200 11424 40000 11536 0 FreeSans 448 0 0 0 proj_in[87]
port 156 nsew signal tristate
flabel metal3 s 39200 28896 40000 29008 0 FreeSans 448 0 0 0 proj_in[88]
port 157 nsew signal tristate
flabel metal3 s 39200 25536 40000 25648 0 FreeSans 448 0 0 0 proj_in[89]
port 158 nsew signal tristate
flabel metal3 s 39200 4704 40000 4816 0 FreeSans 448 0 0 0 proj_in[8]
port 159 nsew signal tristate
flabel metal2 s 23520 39200 23632 40000 0 FreeSans 448 90 0 0 proj_in[90]
port 160 nsew signal tristate
flabel metal2 s 32256 39200 32368 40000 0 FreeSans 448 90 0 0 proj_in[91]
port 161 nsew signal tristate
flabel metal2 s 32928 39200 33040 40000 0 FreeSans 448 90 0 0 proj_in[92]
port 162 nsew signal tristate
flabel metal2 s 24864 39200 24976 40000 0 FreeSans 448 90 0 0 proj_in[93]
port 163 nsew signal tristate
flabel metal3 s 39200 27552 40000 27664 0 FreeSans 448 0 0 0 proj_in[94]
port 164 nsew signal tristate
flabel metal3 s 39200 23520 40000 23632 0 FreeSans 448 0 0 0 proj_in[95]
port 165 nsew signal tristate
flabel metal3 s 39200 32928 40000 33040 0 FreeSans 448 0 0 0 proj_in[96]
port 166 nsew signal tristate
flabel metal3 s 39200 34272 40000 34384 0 FreeSans 448 0 0 0 proj_in[97]
port 167 nsew signal tristate
flabel metal3 s 39200 19488 40000 19600 0 FreeSans 448 0 0 0 proj_in[98]
port 168 nsew signal tristate
flabel metal3 s 39200 17472 40000 17584 0 FreeSans 448 0 0 0 proj_in[99]
port 169 nsew signal tristate
flabel metal3 s 39200 18144 40000 18256 0 FreeSans 448 0 0 0 proj_in[9]
port 170 nsew signal tristate
flabel metal2 s 30240 39200 30352 40000 0 FreeSans 448 90 0 0 proj_rst_n[0]
port 171 nsew signal tristate
flabel metal2 s 12768 39200 12880 40000 0 FreeSans 448 90 0 0 proj_rst_n[1]
port 172 nsew signal tristate
flabel metal2 s 31584 39200 31696 40000 0 FreeSans 448 90 0 0 proj_rst_n[2]
port 173 nsew signal tristate
flabel metal2 s 13440 39200 13552 40000 0 FreeSans 448 90 0 0 proj_rst_n[3]
port 174 nsew signal tristate
flabel metal3 s 39200 28224 40000 28336 0 FreeSans 448 0 0 0 proj_rst_n[4]
port 175 nsew signal tristate
flabel metal2 s 21504 39200 21616 40000 0 FreeSans 448 90 0 0 proj_rst_n[5]
port 176 nsew signal tristate
flabel metal2 s 10080 39200 10192 40000 0 FreeSans 448 90 0 0 proj_rst_n[6]
port 177 nsew signal tristate
flabel metal3 s 39200 30240 40000 30352 0 FreeSans 448 0 0 0 proj_rst_n[7]
port 178 nsew signal tristate
flabel metal2 s 15456 39200 15568 40000 0 FreeSans 448 90 0 0 rst_n
port 179 nsew signal input
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 sel[0]
port 180 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 sel[1]
port 181 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 sel[2]
port 182 nsew signal input
flabel metal4 s 5846 3076 6166 36908 0 FreeSans 1280 90 0 0 vdd
port 183 nsew power bidirectional
flabel metal4 s 15170 3076 15490 36908 0 FreeSans 1280 90 0 0 vdd
port 183 nsew power bidirectional
flabel metal4 s 24494 3076 24814 36908 0 FreeSans 1280 90 0 0 vdd
port 183 nsew power bidirectional
flabel metal4 s 33818 3076 34138 36908 0 FreeSans 1280 90 0 0 vdd
port 183 nsew power bidirectional
flabel metal4 s 10508 3076 10828 36908 0 FreeSans 1280 90 0 0 vss
port 184 nsew ground bidirectional
flabel metal4 s 19832 3076 20152 36908 0 FreeSans 1280 90 0 0 vss
port 184 nsew ground bidirectional
flabel metal4 s 29156 3076 29476 36908 0 FreeSans 1280 90 0 0 vss
port 184 nsew ground bidirectional
flabel metal4 s 38480 3076 38800 36908 0 FreeSans 1280 90 0 0 vss
port 184 nsew ground bidirectional
rlabel metal1 19992 36848 19992 36848 0 vdd
rlabel via1 20072 36064 20072 36064 0 vss
rlabel metal2 22008 25872 22008 25872 0 _000_
rlabel metal2 21000 15232 21000 15232 0 _001_
rlabel metal2 20216 14112 20216 14112 0 _002_
rlabel metal2 20552 14168 20552 14168 0 _003_
rlabel metal2 28280 14224 28280 14224 0 _004_
rlabel metal2 24528 25704 24528 25704 0 _005_
rlabel metal3 21728 29176 21728 29176 0 _006_
rlabel metal2 24248 29904 24248 29904 0 _007_
rlabel metal2 25480 28280 25480 28280 0 _008_
rlabel metal2 21560 29904 21560 29904 0 _009_
rlabel metal2 26600 28616 26600 28616 0 _010_
rlabel metal2 23352 29848 23352 29848 0 _011_
rlabel metal2 27664 27944 27664 27944 0 _012_
rlabel metal2 21896 29848 21896 29848 0 _013_
rlabel metal2 29624 22568 29624 22568 0 _014_
rlabel metal2 30744 22680 30744 22680 0 _015_
rlabel metal2 31080 22848 31080 22848 0 _016_
rlabel metal2 31416 22232 31416 22232 0 _017_
rlabel metal2 32200 21840 32200 21840 0 _018_
rlabel metal2 27720 21224 27720 21224 0 _019_
rlabel metal3 32368 20664 32368 20664 0 _020_
rlabel metal3 30016 20776 30016 20776 0 _021_
rlabel metal2 29848 20328 29848 20328 0 _022_
rlabel metal3 30352 18424 30352 18424 0 _023_
rlabel metal3 29456 16744 29456 16744 0 _024_
rlabel metal2 30520 18928 30520 18928 0 _025_
rlabel metal2 31192 17808 31192 17808 0 _026_
rlabel metal2 31920 17528 31920 17528 0 _027_
rlabel metal2 27384 17472 27384 17472 0 _028_
rlabel metal2 32032 16856 32032 16856 0 _029_
rlabel metal3 28336 16856 28336 16856 0 _030_
rlabel metal2 30240 16856 30240 16856 0 _031_
rlabel metal2 27608 15232 27608 15232 0 _032_
rlabel metal2 28616 14448 28616 14448 0 _033_
rlabel metal2 29904 14392 29904 14392 0 _034_
rlabel metal2 27776 12152 27776 12152 0 _035_
rlabel metal2 28560 12152 28560 12152 0 _036_
rlabel metal2 27608 11592 27608 11592 0 _037_
rlabel metal3 28672 11256 28672 11256 0 _038_
rlabel metal2 23128 14560 23128 14560 0 _039_
rlabel metal2 28056 10472 28056 10472 0 _040_
rlabel metal2 27944 23744 27944 23744 0 _041_
rlabel metal2 24976 23800 24976 23800 0 _042_
rlabel metal2 20776 24808 20776 24808 0 _043_
rlabel metal3 24864 24696 24864 24696 0 _044_
rlabel metal2 14728 18872 14728 18872 0 _045_
rlabel metal2 15064 21952 15064 21952 0 _046_
rlabel via2 14504 25592 14504 25592 0 _047_
rlabel metal3 12712 26152 12712 26152 0 _048_
rlabel metal2 16632 22736 16632 22736 0 _049_
rlabel metal2 12712 25872 12712 25872 0 _050_
rlabel metal2 13552 26264 13552 26264 0 _051_
rlabel metal2 17080 14168 17080 14168 0 _052_
rlabel metal2 15904 15960 15904 15960 0 _053_
rlabel metal2 12432 24808 12432 24808 0 _054_
rlabel metal2 13496 25704 13496 25704 0 _055_
rlabel metal3 14448 26264 14448 26264 0 _056_
rlabel metal2 16632 18088 16632 18088 0 _057_
rlabel metal2 14504 19712 14504 19712 0 _058_
rlabel metal3 13328 23912 13328 23912 0 _059_
rlabel metal3 16688 27608 16688 27608 0 _060_
rlabel metal2 13944 27328 13944 27328 0 _061_
rlabel metal3 16240 28840 16240 28840 0 _062_
rlabel metal2 14392 28840 14392 28840 0 _063_
rlabel metal2 15064 27440 15064 27440 0 _064_
rlabel metal2 14056 29792 14056 29792 0 _065_
rlabel metal3 11536 23912 11536 23912 0 _066_
rlabel metal2 12040 22344 12040 22344 0 _067_
rlabel metal2 12096 22568 12096 22568 0 _068_
rlabel metal2 12600 23464 12600 23464 0 _069_
rlabel metal2 11536 21896 11536 21896 0 _070_
rlabel metal2 12824 21952 12824 21952 0 _071_
rlabel metal2 12376 22288 12376 22288 0 _072_
rlabel metal2 11592 22176 11592 22176 0 _073_
rlabel metal3 11480 21336 11480 21336 0 _074_
rlabel metal3 13216 21560 13216 21560 0 _075_
rlabel metal3 13496 20888 13496 20888 0 _076_
rlabel metal2 12936 20384 12936 20384 0 _077_
rlabel metal2 12712 18032 12712 18032 0 _078_
rlabel metal2 14056 15736 14056 15736 0 _079_
rlabel metal2 12376 16016 12376 16016 0 _080_
rlabel metal3 11760 15960 11760 15960 0 _081_
rlabel metal2 12264 18144 12264 18144 0 _082_
rlabel metal3 13384 18424 13384 18424 0 _083_
rlabel metal3 13496 16072 13496 16072 0 _084_
rlabel metal2 12600 17584 12600 17584 0 _085_
rlabel metal2 11928 18200 11928 18200 0 _086_
rlabel metal2 12712 16576 12712 16576 0 _087_
rlabel metal3 13328 16856 13328 16856 0 _088_
rlabel metal3 11592 16184 11592 16184 0 _089_
rlabel metal2 13048 15624 13048 15624 0 _090_
rlabel metal3 12320 14504 12320 14504 0 _091_
rlabel metal2 13720 13832 13720 13832 0 _092_
rlabel metal2 12712 13888 12712 13888 0 _093_
rlabel metal2 12824 14392 12824 14392 0 _094_
rlabel metal2 13552 22904 13552 22904 0 _095_
rlabel metal2 15624 13272 15624 13272 0 _096_
rlabel metal2 12824 12824 12824 12824 0 _097_
rlabel metal3 11312 12040 11312 12040 0 _098_
rlabel metal3 13048 11368 13048 11368 0 _099_
rlabel metal2 16296 12600 16296 12600 0 _100_
rlabel metal3 13776 12152 13776 12152 0 _101_
rlabel metal3 14280 23128 14280 23128 0 _102_
rlabel metal2 13944 23912 13944 23912 0 _103_
rlabel metal2 14392 24360 14392 24360 0 _104_
rlabel metal2 14392 22456 14392 22456 0 _105_
rlabel metal2 11704 24752 11704 24752 0 _106_
rlabel metal2 14728 24304 14728 24304 0 _107_
rlabel metal2 13552 24696 13552 24696 0 _108_
rlabel metal2 21448 16352 21448 16352 0 _109_
rlabel metal2 22344 23688 22344 23688 0 _110_
rlabel metal3 10192 26264 10192 26264 0 _111_
rlabel metal2 11368 26320 11368 26320 0 _112_
rlabel metal3 22344 23800 22344 23800 0 _113_
rlabel metal2 9800 25368 9800 25368 0 _114_
rlabel metal2 10192 26488 10192 26488 0 _115_
rlabel metal2 11704 25984 11704 25984 0 _116_
rlabel metal2 12600 27776 12600 27776 0 _117_
rlabel metal2 11928 26852 11928 26852 0 _118_
rlabel metal2 11368 20412 11368 20412 0 _119_
rlabel metal2 10696 24528 10696 24528 0 _120_
rlabel metal2 9968 26936 9968 26936 0 _121_
rlabel metal2 10192 24136 10192 24136 0 _122_
rlabel metal2 9688 23856 9688 23856 0 _123_
rlabel metal2 10584 24192 10584 24192 0 _124_
rlabel metal2 10472 22624 10472 22624 0 _125_
rlabel metal2 9968 21784 9968 21784 0 _126_
rlabel metal2 11032 20720 11032 20720 0 _127_
rlabel metal2 10696 21056 10696 21056 0 _128_
rlabel metal2 11368 15568 11368 15568 0 _129_
rlabel metal2 10136 17864 10136 17864 0 _130_
rlabel metal2 8904 16184 8904 16184 0 _131_
rlabel metal2 10136 16016 10136 16016 0 _132_
rlabel metal2 10920 17864 10920 17864 0 _133_
rlabel metal2 11368 17360 11368 17360 0 _134_
rlabel metal2 8792 17920 8792 17920 0 _135_
rlabel metal2 10864 16296 10864 16296 0 _136_
rlabel metal2 10808 15400 10808 15400 0 _137_
rlabel via2 10472 14840 10472 14840 0 _138_
rlabel metal3 9744 14504 9744 14504 0 _139_
rlabel metal3 10136 14392 10136 14392 0 _140_
rlabel metal2 10696 11760 10696 11760 0 _141_
rlabel metal2 11368 11816 11368 11816 0 _142_
rlabel metal2 11144 22568 11144 22568 0 _143_
rlabel metal2 11704 13608 11704 13608 0 _144_
rlabel metal4 18984 23800 18984 23800 0 _145_
rlabel metal2 18872 24360 18872 24360 0 _146_
rlabel metal2 19488 22344 19488 22344 0 _147_
rlabel metal2 19544 24192 19544 24192 0 _148_
rlabel metal2 16856 20608 16856 20608 0 _149_
rlabel metal2 16016 26488 16016 26488 0 _150_
rlabel metal2 13496 21056 13496 21056 0 _151_
rlabel metal2 14840 24416 14840 24416 0 _152_
rlabel metal2 16072 28224 16072 28224 0 _153_
rlabel metal2 14616 20720 14616 20720 0 _154_
rlabel metal2 14168 20720 14168 20720 0 _155_
rlabel metal2 15064 17248 15064 17248 0 _156_
rlabel metal2 14784 17864 14784 17864 0 _157_
rlabel metal2 15176 14168 15176 14168 0 _158_
rlabel metal3 15736 13160 15736 13160 0 _159_
rlabel metal3 22568 26264 22568 26264 0 _160_
rlabel metal2 24136 26040 24136 26040 0 _161_
rlabel metal2 25592 15512 25592 15512 0 _162_
rlabel metal2 26936 25872 26936 25872 0 _163_
rlabel metal2 25592 27608 25592 27608 0 _164_
rlabel metal2 25648 26936 25648 26936 0 _165_
rlabel metal2 26040 28336 26040 28336 0 _166_
rlabel metal2 26936 27328 26936 27328 0 _167_
rlabel metal2 27496 21672 27496 21672 0 _168_
rlabel metal2 28448 27832 28448 27832 0 _169_
rlabel metal2 27160 20384 27160 20384 0 _170_
rlabel metal2 26656 22232 26656 22232 0 _171_
rlabel metal2 27216 21784 27216 21784 0 _172_
rlabel metal2 28448 21560 28448 21560 0 _173_
rlabel metal2 26936 19544 26936 19544 0 _174_
rlabel metal2 27608 20440 27608 20440 0 _175_
rlabel metal2 27664 18536 27664 18536 0 _176_
rlabel metal3 28672 19096 28672 19096 0 _177_
rlabel metal2 28168 18648 28168 18648 0 _178_
rlabel metal2 28112 17528 28112 17528 0 _179_
rlabel metal2 26936 17024 26936 17024 0 _180_
rlabel metal2 27888 16856 27888 16856 0 _181_
rlabel metal2 27384 13832 27384 13832 0 _182_
rlabel metal2 28336 15288 28336 15288 0 _183_
rlabel metal2 28560 13720 28560 13720 0 _184_
rlabel metal2 27496 13216 27496 13216 0 _185_
rlabel metal2 26264 18200 26264 18200 0 _186_
rlabel metal2 27048 14784 27048 14784 0 _187_
rlabel metal2 27272 23464 27272 23464 0 _188_
rlabel metal2 27328 24696 27328 24696 0 _189_
rlabel metal2 21560 26684 21560 26684 0 _190_
rlabel metal2 23016 26264 23016 26264 0 _191_
rlabel metal2 22680 22904 22680 22904 0 _192_
rlabel metal2 22008 21896 22008 21896 0 _193_
rlabel metal2 22736 26936 22736 26936 0 _194_
rlabel metal2 23016 27328 23016 27328 0 _195_
rlabel metal2 23072 27832 23072 27832 0 _196_
rlabel metal2 23576 22288 23576 22288 0 _197_
rlabel metal2 23352 22848 23352 22848 0 _198_
rlabel metal2 23800 19936 23800 19936 0 _199_
rlabel metal2 24192 19992 24192 19992 0 _200_
rlabel metal2 24304 21784 24304 21784 0 _201_
rlabel metal2 24360 21280 24360 21280 0 _202_
rlabel metal2 24416 20216 24416 20216 0 _203_
rlabel metal2 23800 19152 23800 19152 0 _204_
rlabel metal2 24864 19432 24864 19432 0 _205_
rlabel metal2 24696 17472 24696 17472 0 _206_
rlabel metal3 25256 17640 25256 17640 0 _207_
rlabel metal2 25368 17192 25368 17192 0 _208_
rlabel metal2 25368 18144 25368 18144 0 _209_
rlabel metal2 25592 15960 25592 15960 0 _210_
rlabel metal3 21000 16968 21000 16968 0 _211_
rlabel metal2 23016 16240 23016 16240 0 _212_
rlabel metal2 24248 15624 24248 15624 0 _213_
rlabel metal2 22120 16800 22120 16800 0 _214_
rlabel metal2 22680 18480 22680 18480 0 _215_
rlabel metal2 23016 12824 23016 12824 0 _216_
rlabel metal2 23912 13216 23912 13216 0 _217_
rlabel metal2 24136 14056 24136 14056 0 _218_
rlabel metal2 21392 18984 21392 18984 0 _219_
rlabel metal2 22456 18928 22456 18928 0 _220_
rlabel metal2 22008 24696 22008 24696 0 _221_
rlabel metal3 17416 24696 17416 24696 0 _222_
rlabel metal2 18088 29008 18088 29008 0 _223_
rlabel metal3 18200 27048 18200 27048 0 _224_
rlabel metal2 19208 26936 19208 26936 0 _225_
rlabel metal2 18032 21560 18032 21560 0 _226_
rlabel metal2 18816 29624 18816 29624 0 _227_
rlabel metal2 19208 28728 19208 28728 0 _228_
rlabel metal2 19320 27832 19320 27832 0 _229_
rlabel metal2 18760 20832 18760 20832 0 _230_
rlabel metal2 19096 19600 19096 19600 0 _231_
rlabel metal2 19544 21504 19544 21504 0 _232_
rlabel metal2 18760 18368 18760 18368 0 _233_
rlabel metal2 19432 21056 19432 21056 0 _234_
rlabel metal2 19544 20440 19544 20440 0 _235_
rlabel metal2 19656 19096 19656 19096 0 _236_
rlabel metal2 17864 17080 17864 17080 0 _237_
rlabel metal2 18368 16856 18368 16856 0 _238_
rlabel metal2 19096 17192 19096 17192 0 _239_
rlabel metal2 17360 16856 17360 16856 0 _240_
rlabel metal2 18368 17080 18368 17080 0 _241_
rlabel metal2 18984 16072 18984 16072 0 _242_
rlabel metal3 18648 15288 18648 15288 0 _243_
rlabel metal2 17976 13272 17976 13272 0 _244_
rlabel metal3 17248 11368 17248 11368 0 _245_
rlabel metal2 18816 12936 18816 12936 0 _246_
rlabel metal2 16968 19208 16968 19208 0 _247_
rlabel metal2 18984 10864 18984 10864 0 _248_
rlabel metal2 18256 10584 18256 10584 0 _249_
rlabel metal2 19096 13664 19096 13664 0 _250_
rlabel metal2 18536 23912 18536 23912 0 _251_
rlabel metal2 28224 22232 28224 22232 0 _252_
rlabel metal2 27888 26264 27888 26264 0 _253_
rlabel metal2 27384 28840 27384 28840 0 _254_
rlabel metal2 25592 29064 25592 29064 0 _255_
rlabel metal2 25760 29624 25760 29624 0 _256_
rlabel metal2 27216 29624 27216 29624 0 _257_
rlabel metal2 28056 29904 28056 29904 0 _258_
rlabel metal2 31640 21616 31640 21616 0 _259_
rlabel metal2 30184 22848 30184 22848 0 _260_
rlabel metal2 31976 22848 31976 22848 0 _261_
rlabel metal2 31976 19936 31976 19936 0 _262_
rlabel metal2 30128 21000 30128 21000 0 _263_
rlabel metal3 30744 18200 30744 18200 0 _264_
rlabel metal2 30184 18760 30184 18760 0 _265_
rlabel metal2 31976 18928 31976 18928 0 _266_
rlabel metal2 32032 15960 32032 15960 0 _267_
rlabel metal2 30352 15960 30352 15960 0 _268_
rlabel metal3 25144 14392 25144 14392 0 _269_
rlabel metal2 25424 12936 25424 12936 0 _270_
rlabel metal2 25144 13440 25144 13440 0 _271_
rlabel metal3 26320 12376 26320 12376 0 _272_
rlabel metal2 26824 12096 26824 12096 0 _273_
rlabel metal3 28840 23800 28840 23800 0 _274_
rlabel metal2 28896 24696 28896 24696 0 _275_
rlabel metal2 22904 8400 22904 8400 0 _276_
rlabel metal2 22344 9352 22344 9352 0 _277_
rlabel metal2 27608 25872 27608 25872 0 _278_
rlabel metal2 25200 25368 25200 25368 0 _279_
rlabel metal2 26152 10360 26152 10360 0 _280_
rlabel metal2 27496 9408 27496 9408 0 _281_
rlabel metal3 20888 25704 20888 25704 0 _282_
rlabel metal2 15344 24696 15344 24696 0 _283_
rlabel metal2 25368 11928 25368 11928 0 _284_
rlabel metal2 24248 9296 24248 9296 0 _285_
rlabel metal2 23632 25368 23632 25368 0 _286_
rlabel metal2 24024 7952 24024 7952 0 _287_
rlabel metal2 27552 25368 27552 25368 0 _289_
rlabel metal2 20552 25760 20552 25760 0 _290_
rlabel metal2 18424 25984 18424 25984 0 _291_
rlabel metal2 28224 26488 28224 26488 0 _292_
rlabel metal2 34328 2030 34328 2030 0 clk
rlabel metal2 27272 10528 27272 10528 0 clknet_0__276_
rlabel metal3 25088 9688 25088 9688 0 clknet_0_clk
rlabel metal2 21784 10976 21784 10976 0 clknet_1_0__leaf__276_
rlabel metal3 21000 7448 21000 7448 0 clknet_1_0__leaf_clk
rlabel metal2 27832 9744 27832 9744 0 clknet_1_1__leaf__276_
rlabel metal2 27272 8624 27272 8624 0 clknet_1_1__leaf_clk
rlabel metal2 2744 37842 2744 37842 0 in[0]
rlabel metal2 5656 4256 5656 4256 0 in[10]
rlabel metal2 8008 2520 8008 2520 0 in[11]
rlabel metal2 10304 3304 10304 3304 0 in[12]
rlabel metal2 9408 4312 9408 4312 0 in[13]
rlabel metal2 8680 2520 8680 2520 0 in[14]
rlabel metal2 15568 3640 15568 3640 0 in[15]
rlabel metal2 6720 3192 6720 3192 0 in[16]
rlabel metal2 15288 36176 15288 36176 0 in[17]
rlabel metal2 5768 36736 5768 36736 0 in[1]
rlabel metal2 6664 36456 6664 36456 0 in[2]
rlabel metal2 4088 37842 4088 37842 0 in[3]
rlabel metal2 9576 35896 9576 35896 0 in[4]
rlabel metal2 5432 37562 5432 37562 0 in[5]
rlabel metal2 1736 33040 1736 33040 0 in[6]
rlabel metal2 1736 19768 1736 19768 0 in[7]
rlabel metal2 1736 18928 1736 18928 0 in[8]
rlabel metal2 35112 3024 35112 3024 0 in[9]
rlabel metal3 8400 26096 8400 26096 0 net1
rlabel metal2 16968 29120 16968 29120 0 net10
rlabel metal2 12376 5992 12376 5992 0 net100
rlabel metal2 11592 7896 11592 7896 0 net101
rlabel metal2 14168 22288 14168 22288 0 net102
rlabel metal2 13048 25256 13048 25256 0 net103
rlabel metal3 6888 25256 6888 25256 0 net104
rlabel metal2 12376 28280 12376 28280 0 net105
rlabel metal2 11480 30408 11480 30408 0 net106
rlabel metal2 9464 27384 9464 27384 0 net107
rlabel metal2 35336 35504 35336 35504 0 net108
rlabel metal3 6160 24808 6160 24808 0 net109
rlabel metal3 16296 29400 16296 29400 0 net11
rlabel metal2 2072 23576 2072 23576 0 net110
rlabel metal3 5656 22232 5656 22232 0 net111
rlabel metal3 8960 21672 8960 21672 0 net112
rlabel metal2 2184 12264 2184 12264 0 net113
rlabel metal2 11144 17024 11144 17024 0 net114
rlabel metal3 5264 17528 5264 17528 0 net115
rlabel metal2 10248 15400 10248 15400 0 net116
rlabel metal2 9576 13608 9576 13608 0 net117
rlabel metal2 10360 10136 10360 10136 0 net118
rlabel metal2 31304 24024 31304 24024 0 net119
rlabel metal3 18872 29960 18872 29960 0 net12
rlabel metal2 11032 10920 11032 10920 0 net120
rlabel metal3 6776 13832 6776 13832 0 net121
rlabel metal3 31920 24472 31920 24472 0 net122
rlabel metal2 19264 23800 19264 23800 0 net123
rlabel metal2 4200 31304 4200 31304 0 net124
rlabel metal2 8456 32144 8456 32144 0 net125
rlabel metal2 15624 29512 15624 29512 0 net126
rlabel metal2 14728 28168 14728 28168 0 net127
rlabel metal3 14728 21336 14728 21336 0 net128
rlabel metal3 12152 21112 12152 21112 0 net129
rlabel metal2 18144 23240 18144 23240 0 net13
rlabel metal2 32704 21672 32704 21672 0 net130
rlabel metal3 11704 21616 11704 21616 0 net131
rlabel metal3 8400 20440 8400 20440 0 net132
rlabel metal2 15176 17248 15176 17248 0 net133
rlabel metal3 8680 17584 8680 17584 0 net134
rlabel metal3 12824 16800 12824 16800 0 net135
rlabel metal2 2744 13048 2744 13048 0 net136
rlabel metal2 15288 13944 15288 13944 0 net137
rlabel metal2 15736 12376 15736 12376 0 net138
rlabel metal2 10248 7504 10248 7504 0 net139
rlabel metal3 6776 25144 6776 25144 0 net14
rlabel metal2 14392 3388 14392 3388 0 net140
rlabel metal3 34720 20664 34720 20664 0 net141
rlabel metal2 14616 22736 14616 22736 0 net142
rlabel metal3 8400 23744 8400 23744 0 net143
rlabel metal3 27188 36456 27188 36456 0 net144
rlabel metal2 26264 31192 26264 31192 0 net145
rlabel metal2 27216 26936 27216 26936 0 net146
rlabel metal2 29120 36456 29120 36456 0 net147
rlabel metal3 28560 22232 28560 22232 0 net148
rlabel metal2 27832 22400 27832 22400 0 net149
rlabel metal3 8400 20832 8400 20832 0 net15
rlabel metal2 37800 22008 37800 22008 0 net150
rlabel metal3 29512 20664 29512 20664 0 net151
rlabel metal2 29960 20580 29960 20580 0 net152
rlabel metal3 30744 18816 30744 18816 0 net153
rlabel metal3 37072 6664 37072 6664 0 net154
rlabel metal2 28616 17584 28616 17584 0 net155
rlabel metal2 28392 16408 28392 16408 0 net156
rlabel metal3 30380 15512 30380 15512 0 net157
rlabel metal2 29064 13664 29064 13664 0 net158
rlabel metal3 29876 12712 29876 12712 0 net159
rlabel metal3 8596 20104 8596 20104 0 net16
rlabel metal2 27272 14112 27272 14112 0 net160
rlabel metal3 28952 23352 28952 23352 0 net161
rlabel metal2 27832 24472 27832 24472 0 net162
rlabel metal2 30632 14112 30632 14112 0 net163
rlabel metal3 24192 33880 24192 33880 0 net164
rlabel metal2 33880 35952 33880 35952 0 net165
rlabel metal2 34440 36288 34440 36288 0 net166
rlabel metal2 23576 32200 23576 32200 0 net167
rlabel metal2 30408 23296 30408 23296 0 net168
rlabel metal2 35336 23128 35336 23128 0 net169
rlabel metal3 8232 18984 8232 18984 0 net17
rlabel metal2 32088 21784 32088 21784 0 net170
rlabel metal2 31528 28000 31528 28000 0 net171
rlabel metal3 31920 19936 31920 19936 0 net172
rlabel metal2 37912 17304 37912 17304 0 net173
rlabel metal2 32424 17976 32424 17976 0 net174
rlabel metal2 31416 32424 31416 32424 0 net175
rlabel metal2 14896 27608 14896 27608 0 net176
rlabel metal2 33096 29204 33096 29204 0 net177
rlabel metal2 14336 25256 14336 25256 0 net178
rlabel metal2 37688 26936 37688 26936 0 net179
rlabel metal3 31920 18088 31920 18088 0 net18
rlabel metal3 21448 36344 21448 36344 0 net180
rlabel metal2 9744 36456 9744 36456 0 net181
rlabel metal2 28672 26936 28672 26936 0 net182
rlabel metal2 20440 11312 20440 11312 0 net183
rlabel metal2 18704 11144 18704 11144 0 net184
rlabel metal2 24136 7952 24136 7952 0 net185
rlabel metal2 24248 7224 24248 7224 0 net186
rlabel metal3 25312 8232 25312 8232 0 net187
rlabel metal2 22848 7672 22848 7672 0 net188
rlabel metal2 17976 26040 17976 26040 0 net19
rlabel metal2 23688 17304 23688 17304 0 net2
rlabel metal2 21560 3304 21560 3304 0 net20
rlabel metal2 20776 10752 20776 10752 0 net21
rlabel metal2 19712 16072 19712 16072 0 net22
rlabel metal3 33656 4536 33656 4536 0 net23
rlabel metal2 27608 8344 27608 8344 0 net24
rlabel metal2 29960 5096 29960 5096 0 net25
rlabel metal2 32424 5040 32424 5040 0 net26
rlabel metal2 23352 5936 23352 5936 0 net27
rlabel metal2 30632 4256 30632 4256 0 net28
rlabel metal2 26152 5768 26152 5768 0 net29
rlabel metal2 14504 15680 14504 15680 0 net3
rlabel metal2 27496 4200 27496 4200 0 net30
rlabel metal2 37520 36456 37520 36456 0 net31
rlabel metal3 36960 3640 36960 3640 0 net32
rlabel metal3 36848 8232 36848 8232 0 net33
rlabel metal2 24584 15736 24584 15736 0 net34
rlabel metal2 23520 12376 23520 12376 0 net35
rlabel metal2 26768 3528 26768 3528 0 net36
rlabel metal2 25592 4144 25592 4144 0 net37
rlabel metal3 35336 6104 35336 6104 0 net38
rlabel metal2 23296 36456 23296 36456 0 net39
rlabel metal2 14560 15288 14560 15288 0 net4
rlabel metal3 16856 24920 16856 24920 0 net40
rlabel metal2 36232 36008 36232 36008 0 net41
rlabel metal2 37912 8288 37912 8288 0 net42
rlabel metal2 18760 30968 18760 30968 0 net43
rlabel metal3 18984 28504 18984 28504 0 net44
rlabel metal2 19824 28056 19824 28056 0 net45
rlabel metal3 18928 29400 18928 29400 0 net46
rlabel metal2 27048 23744 27048 23744 0 net47
rlabel metal2 20216 22176 20216 22176 0 net48
rlabel metal3 20440 18984 20440 18984 0 net49
rlabel metal2 17752 13104 17752 13104 0 net5
rlabel metal2 19208 14056 19208 14056 0 net50
rlabel metal2 14672 15512 14672 15512 0 net51
rlabel metal3 17304 15176 17304 15176 0 net52
rlabel metal2 30744 13384 30744 13384 0 net53
rlabel metal2 17976 4256 17976 4256 0 net54
rlabel metal2 18648 3304 18648 3304 0 net55
rlabel metal3 17752 10696 17752 10696 0 net56
rlabel metal2 17304 7112 17304 7112 0 net57
rlabel metal2 18872 14336 18872 14336 0 net58
rlabel metal3 17360 36344 17360 36344 0 net59
rlabel metal2 19768 11032 19768 11032 0 net6
rlabel metal2 32312 35056 32312 35056 0 net60
rlabel metal2 27384 34608 27384 34608 0 net61
rlabel metal3 29176 35336 29176 35336 0 net62
rlabel metal3 29176 33544 29176 33544 0 net63
rlabel metal2 30408 13664 30408 13664 0 net64
rlabel metal3 33768 23240 33768 23240 0 net65
rlabel metal2 32424 26712 32424 26712 0 net66
rlabel metal2 32256 21336 32256 21336 0 net67
rlabel metal3 34048 21672 34048 21672 0 net68
rlabel metal3 31612 18984 31612 18984 0 net69
rlabel metal2 16352 12040 16352 12040 0 net7
rlabel metal3 35112 7560 35112 7560 0 net70
rlabel metal2 32536 14728 32536 14728 0 net71
rlabel metal2 30856 16072 30856 16072 0 net72
rlabel metal2 28168 13608 28168 13608 0 net73
rlabel metal3 30688 11144 30688 11144 0 net74
rlabel metal2 37240 12544 37240 12544 0 net75
rlabel metal2 27160 11424 27160 11424 0 net76
rlabel metal2 27440 10360 27440 10360 0 net77
rlabel metal2 29512 24304 29512 24304 0 net78
rlabel metal2 29568 24920 29568 24920 0 net79
rlabel metal2 17248 22120 17248 22120 0 net8
rlabel metal2 29400 4032 29400 4032 0 net80
rlabel metal2 28616 5964 28616 5964 0 net81
rlabel metal3 37800 32536 37800 32536 0 net82
rlabel metal2 35336 25872 35336 25872 0 net83
rlabel metal3 10808 26488 10808 26488 0 net84
rlabel metal2 3640 32816 3640 32816 0 net85
rlabel metal2 21784 31584 21784 31584 0 net86
rlabel metal2 14336 29624 14336 29624 0 net87
rlabel metal2 13720 31864 13720 31864 0 net88
rlabel metal2 5096 24192 5096 24192 0 net89
rlabel metal2 17416 23856 17416 23856 0 net9
rlabel metal2 2184 22624 2184 22624 0 net90
rlabel metal3 7952 21784 7952 21784 0 net91
rlabel metal2 12600 19936 12600 19936 0 net92
rlabel metal3 8400 18368 8400 18368 0 net93
rlabel metal2 2632 8288 2632 8288 0 net94
rlabel metal2 2072 7728 2072 7728 0 net95
rlabel metal2 2072 11424 2072 11424 0 net96
rlabel metal2 23688 31584 23688 31584 0 net97
rlabel metal2 2072 14224 2072 14224 0 net98
rlabel metal2 10920 7616 10920 7616 0 net99
rlabel metal2 32984 2086 32984 2086 0 proj_clk[0]
rlabel metal2 32312 1358 32312 1358 0 proj_clk[1]
rlabel metal2 28952 1022 28952 1022 0 proj_clk[2]
rlabel metal2 30968 2086 30968 2086 0 proj_clk[3]
rlabel metal2 22904 2030 22904 2030 0 proj_clk[4]
rlabel metal2 29624 910 29624 910 0 proj_clk[5]
rlabel metal2 24920 2058 24920 2058 0 proj_clk[6]
rlabel metal2 26264 2058 26264 2058 0 proj_clk[7]
rlabel metal2 37352 36624 37352 36624 0 proj_in[0]
rlabel metal3 38738 3416 38738 3416 0 proj_in[100]
rlabel metal2 37576 7728 37576 7728 0 proj_in[101]
rlabel metal2 38304 15848 38304 15848 0 proj_in[102]
rlabel metal2 23576 1302 23576 1302 0 proj_in[103]
rlabel metal2 25592 854 25592 854 0 proj_in[104]
rlabel metal2 25256 3472 25256 3472 0 proj_in[105]
rlabel metal2 38248 5712 38248 5712 0 proj_in[106]
rlabel metal2 23016 36344 23016 36344 0 proj_in[107]
rlabel metal2 16352 35896 16352 35896 0 proj_in[108]
rlabel metal3 35504 36344 35504 36344 0 proj_in[109]
rlabel metal3 38738 8120 38738 8120 0 proj_in[10]
rlabel metal2 18200 37786 18200 37786 0 proj_in[110]
rlabel metal2 17528 37786 17528 37786 0 proj_in[111]
rlabel metal2 20216 37786 20216 37786 0 proj_in[112]
rlabel metal2 18872 37786 18872 37786 0 proj_in[113]
rlabel metal2 34440 35896 34440 35896 0 proj_in[114]
rlabel metal2 21000 36344 21000 36344 0 proj_in[115]
rlabel metal2 20888 2030 20888 2030 0 proj_in[116]
rlabel metal2 19544 2030 19544 2030 0 proj_in[117]
rlabel metal2 16856 2058 16856 2058 0 proj_in[118]
rlabel metal2 6104 2030 6104 2030 0 proj_in[119]
rlabel metal3 38584 9576 38584 9576 0 proj_in[11]
rlabel metal2 18200 2030 18200 2030 0 proj_in[120]
rlabel metal2 18872 2030 18872 2030 0 proj_in[121]
rlabel metal2 16296 4424 16296 4424 0 proj_in[122]
rlabel metal2 17528 2030 17528 2030 0 proj_in[123]
rlabel metal2 7448 2030 7448 2030 0 proj_in[124]
rlabel metal2 16408 36624 16408 36624 0 proj_in[125]
rlabel metal2 31192 37072 31192 37072 0 proj_in[126]
rlabel metal2 27160 36680 27160 36680 0 proj_in[127]
rlabel metal3 30128 36232 30128 36232 0 proj_in[128]
rlabel metal2 29736 37016 29736 37016 0 proj_in[129]
rlabel metal2 38304 11144 38304 11144 0 proj_in[12]
rlabel metal2 37576 35728 37576 35728 0 proj_in[130]
rlabel metal2 38248 29848 38248 29848 0 proj_in[131]
rlabel metal3 38248 25088 38248 25088 0 proj_in[132]
rlabel metal2 38248 21280 38248 21280 0 proj_in[133]
rlabel metal3 38584 18984 38584 18984 0 proj_in[134]
rlabel metal2 38248 7168 38248 7168 0 proj_in[135]
rlabel metal2 38248 8960 38248 8960 0 proj_in[136]
rlabel metal2 38248 16576 38248 16576 0 proj_in[137]
rlabel metal3 38584 14280 38584 14280 0 proj_in[138]
rlabel metal2 30296 854 30296 854 0 proj_in[139]
rlabel metal2 37576 12432 37576 12432 0 proj_in[13]
rlabel metal2 31640 2030 31640 2030 0 proj_in[140]
rlabel metal2 26936 2590 26936 2590 0 proj_in[141]
rlabel metal2 38248 35392 38248 35392 0 proj_in[142]
rlabel metal3 38402 31640 38402 31640 0 proj_in[143]
rlabel metal2 28280 2086 28280 2086 0 proj_in[14]
rlabel metal2 27608 854 27608 854 0 proj_in[15]
rlabel metal2 38248 32480 38248 32480 0 proj_in[16]
rlabel metal2 38192 26936 38192 26936 0 proj_in[17]
rlabel metal2 7448 37786 7448 37786 0 proj_in[18]
rlabel metal2 3416 37786 3416 37786 0 proj_in[19]
rlabel metal2 22344 36344 22344 36344 0 proj_in[1]
rlabel metal2 10696 36344 10696 36344 0 proj_in[20]
rlabel metal2 12040 36344 12040 36344 0 proj_in[21]
rlabel metal3 1246 30968 1246 30968 0 proj_in[22]
rlabel metal3 1246 22904 1246 22904 0 proj_in[23]
rlabel metal3 854 29624 854 29624 0 proj_in[24]
rlabel metal3 1246 32312 1246 32312 0 proj_in[25]
rlabel metal3 1246 18200 1246 18200 0 proj_in[26]
rlabel metal3 1582 7448 1582 7448 0 proj_in[27]
rlabel metal3 1246 8120 1246 8120 0 proj_in[28]
rlabel metal3 854 10808 854 10808 0 proj_in[29]
rlabel metal2 25256 36512 25256 36512 0 proj_in[2]
rlabel metal3 1246 14168 1246 14168 0 proj_in[30]
rlabel metal2 11480 2030 11480 2030 0 proj_in[31]
rlabel metal2 12824 2030 12824 2030 0 proj_in[32]
rlabel metal2 12152 2030 12152 2030 0 proj_in[33]
rlabel metal3 1582 26936 1582 26936 0 proj_in[34]
rlabel metal3 1246 25592 1246 25592 0 proj_in[35]
rlabel metal3 1302 26264 1302 26264 0 proj_in[36]
rlabel metal3 1246 28280 1246 28280 0 proj_in[37]
rlabel metal2 11368 36344 11368 36344 0 proj_in[38]
rlabel metal3 1246 27608 1246 27608 0 proj_in[39]
rlabel metal2 34888 37016 34888 37016 0 proj_in[3]
rlabel metal3 1246 24248 1246 24248 0 proj_in[40]
rlabel metal3 1246 23576 1246 23576 0 proj_in[41]
rlabel metal3 1246 22232 1246 22232 0 proj_in[42]
rlabel metal3 1246 30296 1246 30296 0 proj_in[43]
rlabel metal3 1246 11480 1246 11480 0 proj_in[44]
rlabel metal3 854 15512 854 15512 0 proj_in[45]
rlabel metal3 1246 17528 1246 17528 0 proj_in[46]
rlabel metal3 1246 9464 1246 9464 0 proj_in[47]
rlabel metal3 1246 12824 1246 12824 0 proj_in[48]
rlabel metal3 1246 8792 1246 8792 0 proj_in[49]
rlabel metal2 38248 24528 38248 24528 0 proj_in[4]
rlabel metal3 1246 10136 1246 10136 0 proj_in[50]
rlabel metal3 1246 13496 1246 13496 0 proj_in[51]
rlabel metal2 36680 36512 36680 36512 0 proj_in[52]
rlabel metal2 19544 37786 19544 37786 0 proj_in[53]
rlabel metal2 4704 36344 4704 36344 0 proj_in[54]
rlabel metal2 8792 37786 8792 37786 0 proj_in[55]
rlabel metal2 14112 36344 14112 36344 0 proj_in[56]
rlabel metal2 8120 37786 8120 37786 0 proj_in[57]
rlabel metal3 854 21560 854 21560 0 proj_in[58]
rlabel metal3 1582 31640 1582 31640 0 proj_in[59]
rlabel metal2 38304 31528 38304 31528 0 proj_in[5]
rlabel metal3 1246 20888 1246 20888 0 proj_in[60]
rlabel metal3 1246 20216 1246 20216 0 proj_in[61]
rlabel metal3 1246 16184 1246 16184 0 proj_in[62]
rlabel metal3 1582 16856 1582 16856 0 proj_in[63]
rlabel metal3 1246 14840 1246 14840 0 proj_in[64]
rlabel metal3 1582 12152 1582 12152 0 proj_in[65]
rlabel metal2 14840 2030 14840 2030 0 proj_in[66]
rlabel metal2 13440 3416 13440 3416 0 proj_in[67]
rlabel metal2 10808 1190 10808 1190 0 proj_in[68]
rlabel metal2 14168 2030 14168 2030 0 proj_in[69]
rlabel metal2 38248 33936 38248 33936 0 proj_in[6]
rlabel metal3 1246 28952 1246 28952 0 proj_in[70]
rlabel metal3 1246 24920 1246 24920 0 proj_in[71]
rlabel metal2 27272 36624 27272 36624 0 proj_in[72]
rlabel metal2 26600 36512 26600 36512 0 proj_in[73]
rlabel metal2 28392 36736 28392 36736 0 proj_in[74]
rlabel metal3 28784 36232 28784 36232 0 proj_in[75]
rlabel metal2 37576 26992 37576 26992 0 proj_in[76]
rlabel metal2 38248 23072 38248 23072 0 proj_in[77]
rlabel metal3 38738 22232 38738 22232 0 proj_in[78]
rlabel metal2 38304 20552 38304 20552 0 proj_in[79]
rlabel metal2 37576 21840 37576 21840 0 proj_in[7]
rlabel metal2 38248 4256 38248 4256 0 proj_in[80]
rlabel metal2 38248 6328 38248 6328 0 proj_in[81]
rlabel metal2 37576 17136 37576 17136 0 proj_in[82]
rlabel metal2 38248 10416 38248 10416 0 proj_in[83]
rlabel metal2 38248 15120 38248 15120 0 proj_in[84]
rlabel metal3 38738 12824 38738 12824 0 proj_in[85]
rlabel metal2 38248 13664 38248 13664 0 proj_in[86]
rlabel metal2 38248 11872 38248 11872 0 proj_in[87]
rlabel metal2 38248 29232 38248 29232 0 proj_in[88]
rlabel metal2 38248 25984 38248 25984 0 proj_in[89]
rlabel metal3 38584 4872 38584 4872 0 proj_in[8]
rlabel metal2 24584 36400 24584 36400 0 proj_in[90]
rlabel metal2 33544 37072 33544 37072 0 proj_in[91]
rlabel metal3 33600 36344 33600 36344 0 proj_in[92]
rlabel metal2 25928 36624 25928 36624 0 proj_in[93]
rlabel metal2 38248 27776 38248 27776 0 proj_in[94]
rlabel metal3 38584 23688 38584 23688 0 proj_in[95]
rlabel metal3 38584 33096 38584 33096 0 proj_in[96]
rlabel metal2 38304 34664 38304 34664 0 proj_in[97]
rlabel metal2 38248 19824 38248 19824 0 proj_in[98]
rlabel metal3 38738 17528 38738 17528 0 proj_in[99]
rlabel metal2 38248 18368 38248 18368 0 proj_in[9]
rlabel metal2 31080 37016 31080 37016 0 proj_rst_n[0]
rlabel metal2 12600 37016 12600 37016 0 proj_rst_n[1]
rlabel metal2 31640 38066 31640 38066 0 proj_rst_n[2]
rlabel metal2 13440 36344 13440 36344 0 proj_rst_n[3]
rlabel metal3 38584 28392 38584 28392 0 proj_rst_n[4]
rlabel metal2 21672 36344 21672 36344 0 proj_rst_n[5]
rlabel metal2 10024 36344 10024 36344 0 proj_rst_n[6]
rlabel metal2 38248 30688 38248 30688 0 proj_rst_n[7]
rlabel metal2 15568 36456 15568 36456 0 rst_n
rlabel metal2 21840 3080 21840 3080 0 sel[0]
rlabel metal2 22456 2520 22456 2520 0 sel[1]
rlabel metal2 20328 4200 20328 4200 0 sel[2]
rlabel metal2 23240 10416 23240 10416 0 sel_reg\[0\]
rlabel metal2 24192 11480 24192 11480 0 sel_reg\[1\]
rlabel metal2 22120 7728 22120 7728 0 sel_reg\[2\]
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
