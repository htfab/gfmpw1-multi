* NGSPICE file created from cells9.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2 D RN SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__mux2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__mux2_1 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2 D SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlya_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlya_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_16 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_16 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 D SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffq_1 D SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2 D RN SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyc_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyc_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__mux2_4 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlya_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlya_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__addf_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__addf_2 A B CI CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffq_4 D SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__invz_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__invz_2 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1 D RN SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_1 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latq_2 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4 D RN SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__icgtp_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__icgtp_4 CLK E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latrnq_2 D E RN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_4 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latsnq_1 D E SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_16 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_16 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_20 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyd_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyd_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_12 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_12 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 D RN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyb_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyb_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__invz_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__invz_8 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1 D SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latsnq_4 D E SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai33_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai33_4 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1 D RN SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2 D RN SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1 D SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffsnq_1 D SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1 D RN SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4 D SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyc_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4 D RN SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4 D SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__addf_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__addf_1 A B CI CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_16 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 D SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4 D RN SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__invz_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__invz_1 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyc_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyc_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_12 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_12 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__addh_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__addh_2 A B CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latrsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latrsnq_2 D E RN SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__icgtn_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__icgtn_2 CLKN E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__addf_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__addf_4 A B CI CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__invz_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__invz_4 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latrnq_1 D E RN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_3 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_3 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_20 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_20 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyd_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnq_2 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latq_4 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1 D RN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latrnq_4 D E RN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1 D RN SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyd_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyd_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4 D RN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or3_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4 D RN SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__hold abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__hold Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_16 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_16 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__icgtp_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__icgtp_2 CLK E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffq_2 D SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__invz_12 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__invz_12 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__addh_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__addh_1 A B CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latrsnq_1 D E RN SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__icgtn_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__icgtn_1 CLKN E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__invz_3 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__invz_3 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2 D RN SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_2 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__addh_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__addh_4 A B CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latrsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latrsnq_4 D E RN SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__icgtn_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__icgtn_4 CLKN E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_20 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_20 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnq_1 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyb_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyb_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latsnq_2 D E SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai33_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai33_2 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnq_4 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_12 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_12 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2 D SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_8 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

.subckt cells9 clk in[0] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[1]
+ in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] out[0] out[10] out[11] out[1] out[2]
+ out[3] out[4] out[5] out[6] out[7] out[8] out[9] rst_n vdd vss
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_415 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_501_ _005_ in[0] cm_inst.page\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XANTENNA__365__S _133_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nor3_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_432_ _107_ _197_ _031_ _198_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XTAP_TAPCELL_ROW_51_481 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_51_470 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_294_ cm_inst.cc_inst.out_notouch_\[65\] cm_inst.cc_inst.out_notouch_\[73\] cm_inst.cc_inst.out_notouch_\[81\]
+ cm_inst.cc_inst.out_notouch_\[89\] _060_ _064_ _065_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA__424__S1 _095_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_23_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_363_ cm_inst.cc_inst.out_notouch_\[131\] cm_inst.cc_inst.out_notouch_\[139\] cm_inst.cc_inst.out_notouch_\[147\]
+ cm_inst.cc_inst.out_notouch_\[155\] _094_ _095_ _132_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.oai33_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_2_inst_B3 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_170 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.oai31_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_214 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_10_453 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__249__I _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.buf_3_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_263 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.dffrsnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[154\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2
XTAP_TAPCELL_ROW_5_151 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__506__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_415_ _179_ _181_ _030_ _182_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_346_ _106_ _110_ _045_ _115_ _116_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
XFILLER_0_51_342 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.aoi221_1_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_36_361 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_277_ cm_inst.cc_inst.out_notouch_\[160\] cm_inst.cc_inst.out_notouch_\[168\] cm_inst.cc_inst.out_notouch_\[176\]
+ cm_inst.cc_inst.out_notouch_\[184\] _048_ _023_ _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XPHY_EDGE_ROW_20_Left_72 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_6_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_6_255 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.xor3_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_42_375 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__492__A3 in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_37_158 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_289 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_350 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_16_223 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[20\].div_flop ro_inst.counter_n\[20\] in[0] ro_inst.counter_n\[19\]
+ ro_inst.counter\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
X_329_ _098_ _046_ _099_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
XFILLER_0_51_172 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_3_236 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.dlyd_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffq_4_inst_SE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_51_70 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA__262__I _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_42_183 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_367 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_38_381 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_434 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_412 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_13_204 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_172 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_29_434 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.and3_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and3_2
XFILLER_0_29_467 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nand2_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_12_312 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_389 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.icgtp_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.nor4_4_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_35_362 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_35_415 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.sdffsnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[169\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xcm_inst.cc_inst.mux2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[117\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_30_131 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.nand4_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.clkbuf_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[191\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_4
XPHY_EDGE_ROW_51_Left_103 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_ro_inst.gcount\[30\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.latq_4_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_41_398 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_34_470 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai222_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_49_454 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_32_61 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_17_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_44_289 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.dffq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.aoi222_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_7_191 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi222_4_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.latrnq_1_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_46_435 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.invz_1_inst_EN cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_4_183 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dlya_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[176\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlya_1
XFILLER_0_13_440 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_13_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.xnor3_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor3_2
X_500_ _004_ in[0] cm_inst.page\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XFILLER_0_48_381 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_416 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_362_ cm_inst.cc_inst.out_notouch_\[163\] cm_inst.cc_inst.out_notouch_\[171\] cm_inst.cc_inst.out_notouch_\[179\]
+ cm_inst.cc_inst.out_notouch_\[187\] _094_ _078_ _131_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_431_ cm_inst.cc_inst.out_notouch_\[70\] cm_inst.cc_inst.out_notouch_\[78\] _038_
+ _197_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_51_502 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_471 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_293_ _063_ _064_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA_cm_inst.cc_inst.oai33_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_3_18 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_8_171 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nand3_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_3_29 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_14_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_ro_inst.gcount\[9\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_9_286 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_207 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__376__S _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_5_152 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.clkinv_12_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_345_ _112_ _114_ _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XFILLER_0_28_307 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
X_414_ cm_inst.cc_inst.out_notouch_\[69\] cm_inst.cc_inst.out_notouch_\[77\] cm_inst.cc_inst.out_notouch_\[85\]
+ cm_inst.cc_inst.out_notouch_\[93\] _142_ _180_ _181_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_276_ _019_ _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
Xro_inst.gcount\[10\].div_flop ro_inst.counter_n\[10\] in[0] ro_inst.counter_n\[9\]
+ ro_inst.counter\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_51_376 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.aoi221_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi221_1_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_395 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_11_207 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_42_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_95 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.xor3_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.mux4_2_inst_S0 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_2_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_251 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_295 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA__492__A4 in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.addf_1_inst_CI cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_33_354 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_33_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.oai21_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_115 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_224 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_328_ _061_ _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
X_259_ _030_ _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.clkinv_16_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[202\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_16
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dffsnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[157\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffsnq_2
XFILLER_0_30_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_343 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_15_398 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_30_379 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_38_382 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SE cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_446 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_424 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_13_205 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_21_260 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_184 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA__402__B _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_446 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_307 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_63 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nand2_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.sdffq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[159\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffq_1
XANTENNA_cm_inst.cc_inst.dffnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_47_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_35_449 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.nand4_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_198 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dffnrsnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[142\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2
XANTENNA_cm_inst.cc_inst.latq_4_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__454__S0 _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_41_399 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_26_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_21_132 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_49_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_49_455 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_243 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_221 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.oai32_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[90\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai32_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_4_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_12_187 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_35_268 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_493 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_18 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.latrsnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_46_436 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.latrnq_1_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_224 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.inv_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_2
XFILLER_0_1_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_22_430 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.mux2_1_inst_I0 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_202 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_257 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_51_472 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_43_417 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_292_ cm_inst.page\[1\] _063_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_361_ _130_ ro_inst.counter\[2\] _016_ out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_430_ _102_ cm_inst.cc_inst.out_notouch_\[86\] _195_ _037_ _196_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi211_1
Xro_inst.gcount\[7\].div_flop ro_inst.counter_n\[7\] in[0] ro_inst.counter_n\[6\]
+ ro_inst.counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_8_172 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nand3_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_9_298 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_271 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_413_ _063_ _180_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA_cm_inst.cc_inst.aoi21_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi221_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_344_ cm_inst.cc_inst.out_notouch_\[98\] cm_inst.cc_inst.out_notouch_\[106\] cm_inst.cc_inst.out_notouch_\[114\]
+ cm_inst.cc_inst.out_notouch_\[122\] _085_ _113_ _114_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_275_ _017_ _047_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XTAP_TAPCELL_ROW_11_188 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_19_244 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_42_333 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.mux4_2_inst_S1 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_SE cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_10_263 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_33_300 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_18_374 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai21_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_16_225 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[8\].div_flop_inv ro_inst.counter\[8\] ro_inst.counter_n\[8\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
Xcm_inst.cc_inst.mux4_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[121\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_2
XFILLER_0_36_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_258_ _029_ _030_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_24_366 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_333 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_24_280 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_327_ _092_ _096_ _051_ _097_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA_ro_inst.gcount\[26\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.inv_16_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_347 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_383 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_13_206 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_130 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_21_261 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_196 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xro_inst.gcount\[33\].div_flop_inv ro_inst.counter\[33\] ro_inst.counter_n\[33\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.and2_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_403 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_24_174 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_24_152 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[14\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.aoi21_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[68\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_4
XFILLER_0_20_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_43_450 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_417 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_483 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.nand4_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.dffrnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dlyb_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_233 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_494 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_461 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dlyc_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[183\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyc_2
XTAP_TAPCELL_ROW_49_456 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_29_277 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_255 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_40_453 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_155 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_12_199 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai211_2_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_35_203 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_31_431 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_160 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_46_437 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.oai222_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[103\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai222_2
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__509__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.mux2_1_inst_I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_225 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_269 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_40_294 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_37_Left_89 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_51_473 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_43_418 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_291_ cm_inst.cc_inst.out_notouch_\[97\] cm_inst.cc_inst.out_notouch_\[105\] cm_inst.cc_inst.out_notouch_\[113\]
+ cm_inst.cc_inst.out_notouch_\[121\] _060_ _061_ _062_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_360_ _047_ _101_ _128_ _129_ _130_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
Xro_inst.gcount\[26\].div_flop_inv ro_inst.counter\[26\] ro_inst.counter_n\[26\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_31_294 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_23_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_48_Left_100 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_8_173 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nand3_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_501 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_489_ in[7] cm_inst.cc_inst.in\[5\] _238_ _011_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_38_51 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_22_294 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_49_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_9_266 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
X_412_ cm_inst.cc_inst.out_notouch_\[101\] cm_inst.cc_inst.out_notouch_\[109\] cm_inst.cc_inst.out_notouch_\[117\]
+ cm_inst.cc_inst.out_notouch_\[125\] _142_ _138_ _179_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.aoi21_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_375 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_36_364 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.addf_4_inst_A cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__472__I in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_343_ _022_ _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_24_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_189 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_274_ _044_ _045_ _046_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XANTENNA__494__I0 in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_19_245 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_42_367 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__382__I _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_507 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_27_364 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_236 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_15_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__485__I0 in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_33_323 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_33_312 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__292__I cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.mux2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[119\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_4
XANTENNA__476__I0 in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_3_inst_I cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_326_ cm_inst.cc_inst.out_notouch_\[130\] cm_inst.cc_inst.out_notouch_\[138\] cm_inst.cc_inst.out_notouch_\[146\]
+ cm_inst.cc_inst.out_notouch_\[154\] _094_ _095_ _096_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XTAP_TAPCELL_ROW_16_226 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_257_ cm_inst.page\[2\] _029_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
XFILLER_0_24_389 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_24_281 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_24_Left_76 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_3_228 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_12_507 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.and4_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_183 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_359 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_337 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_30_326 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_38_404 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[19\].div_flop_inv ro_inst.counter\[19\] ro_inst.counter_n\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XTAP_TAPCELL_ROW_13_207 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_109 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_21_262 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.and2_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_415 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__377__A2 _145_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_309_ _077_ _079_ _051_ _080_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_21_10 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi211_2_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.dlya_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[178\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlya_4
XANTENNA_cm_inst.cc_inst.nand4_4_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_134 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.inv_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.or2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[46\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or2_2
XTAP_TAPCELL_ROW_49_457 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_223 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_32_335 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_8_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_12_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai211_2_inst_C cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.nor2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[36\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__381__S1 _095_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_11_Left_63 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_35_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xcm_inst.cc_inst.addf_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[107\] cm_inst.cc_inst.out_notouch_\[108\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu9t5v0__addf_2
XANTENNA__372__S1 _064_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.nand2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XTAP_TAPCELL_ROW_46_438 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__363__S1 _095_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_8_inst_EN cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_443 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_51_474 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.latsnq_2_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_290_ cm_inst.page\[1\] _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_8_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_16_281 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_16_292 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_488_ in[6] cm_inst.cc_inst.in\[4\] _240_ _010_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_42_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_218 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_251 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.mux2_2_inst_S cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_245 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.addf_4_inst_B cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_342_ _111_ _112_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
X_411_ _173_ _176_ _177_ _155_ _178_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_273_ cm_inst.page\[3\] _045_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XANTENNA__263__S0 _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_19_246 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_42_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_379 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_335 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.sdffq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[161\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffq_4
XANTENNA__485__I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_2_125 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.aoi222_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[79\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi222_2
XFILLER_0_18_343 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_18_354 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_36_162 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_24_282 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_325_ _022_ _095_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XTAP_TAPCELL_ROW_16_227 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_256_ cm_inst.cc_inst.out_notouch_\[0\] cm_inst.cc_inst.out_notouch_\[8\] cm_inst.cc_inst.out_notouch_\[16\]
+ cm_inst.cc_inst.out_notouch_\[24\] _021_ _024_ _028_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA__432__B _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_76 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_47_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffq_4_inst_SI cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.oai32_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[92\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai32_4
XANTENNA_cm_inst.cc_inst.and4_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_305 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.aoi211_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_41_Left_93 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_38_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_13_208 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_176 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_21_263 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.oai21_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[81\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XANTENNA__478__I in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_154 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_4_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_308_ cm_inst.cc_inst.out_notouch_\[129\] cm_inst.cc_inst.out_notouch_\[137\] cm_inst.cc_inst.out_notouch_\[145\]
+ cm_inst.cc_inst.out_notouch_\[153\] _020_ _078_ _079_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
Xro_inst.gcount\[4\].div_flop_inv ro_inst.counter\[4\] ro_inst.counter_n\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.aoi211_2_inst_C cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_463 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_452 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_43_430 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_30_168 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.icgtn_1_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_224 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_452 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_474 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_1_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_21_124 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_458 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_32_336 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_257 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_235 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_40_391 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_37_290 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.invz_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[174\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__invz_2
XFILLER_0_25_430 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_40_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.bufz_4_inst_EN cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.sdffrsnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[165\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1
XANTENNA_cm_inst.cc_inst.addh_2_inst_A cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_411 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_7_195 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_190 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_439 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_500 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_22_400 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_22_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_187 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[6\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_51_506 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_51_475 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.latsnq_2_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_31_274 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.or2_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_39_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_487_ in[5] cm_inst.cc_inst.in\[3\] _240_ _009_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_6_419 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xcm_inst.cc_inst.bufz_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[171\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_1
XFILLER_0_38_86 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_22_296 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_224 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_257 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_263 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_36_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_410_ cm_inst.cc_inst.out_notouch_\[197\] cm_inst.cc_inst.out_notouch_\[205\] _039_
+ _177_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_341_ cm_inst.page\[2\] _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
X_272_ _029_ _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XANTENNA__263__S1 _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_290 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.dffq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[22\].div_flop_inv ro_inst.counter\[22\] ro_inst.counter_n\[22\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
Xcm_inst.cc_inst.and2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
XTAP_TAPCELL_ROW_19_247 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_42_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_39_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_27_366 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_27_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_27_300 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_24_77 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_6_216 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_222 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_255 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_2_126 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_10_299 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[6\].div_flop ro_inst.counter_n\[6\] in[0] ro_inst.counter_n\[5\]
+ ro_inst.counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_18_300 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_18_333 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_33_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_5_293 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_366 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_16_228 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_24_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_24_283 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_324_ _093_ _094_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_255_ cm_inst.cc_inst.out_notouch_\[32\] cm_inst.cc_inst.out_notouch_\[40\] cm_inst.cc_inst.out_notouch_\[48\]
+ cm_inst.cc_inst.out_notouch_\[56\] _021_ _024_ _027_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.buf_20_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_358 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_108 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.and4_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_2_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_23_380 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai21_4_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi211_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SI cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.clkbuf_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_428 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_141 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_21_328 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_21_264 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.nor4_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor4_2
XTAP_TAPCELL_ROW_29_320 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_417 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_24_100 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_24_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_307_ _022_ _078_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XANTENNA_cm_inst.cc_inst.clkbuf_16_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__385__I1 _152_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.nand4_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand4_2
XFILLER_0_20_394 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_35_356 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_43_442 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_7_399 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_15_155 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.oai211_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[97\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_2
Xcm_inst.cc_inst.xnor2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[54\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor2_1
XFILLER_0_34_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[15\].div_flop_inv ro_inst.counter\[15\] ro_inst.counter_n\[15\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.xnor2_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_49_459 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.latrnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_32_337 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_392 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.addh_2_inst_B cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_453 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_497 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_434 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_261 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_25_250 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_17_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or4_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_294 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_412 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_51_476 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_8_461 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.or2_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_42_410 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_342 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_486_ in[4] cm_inst.cc_inst.in\[2\] _240_ _008_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_9_236 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_5_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__488__I0 in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_5_146 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_13_275 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_271_ cm_inst.cc_inst.out_notouch_\[208\] _040_ _042_ _037_ _043_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi22_1
X_340_ _107_ _109_ _031_ _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XANTENNA_cm_inst.cc_inst.inv_8_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_45 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_19_248 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_183 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_27_323 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_469_ _232_ ro_inst.signal vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_50_381 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_49_20 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_2_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_181 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_2_127 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_SI cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_18_378 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_33_326 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[23\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_5_261 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xcm_inst.cc_inst.aoi22_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[69\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XANTENNA_cm_inst.cc_inst.nor3_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_16_229 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_36_164 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_36_131 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_323_ cm_inst.page\[0\] _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XTAP_TAPCELL_ROW_24_284 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_24_337 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_209 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_254_ cm_inst.cc_inst.out_notouch_\[64\] cm_inst.cc_inst.out_notouch_\[72\] cm_inst.cc_inst.out_notouch_\[80\]
+ cm_inst.cc_inst.out_notouch_\[88\] _021_ _024_ _026_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.and4_2_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.nor2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[38\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_4
XANTENNA_ro_inst.gcount\[11\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_46_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.nand2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_4
XFILLER_0_37_440 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_407 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_306_ cm_inst.cc_inst.out_notouch_\[161\] cm_inst.cc_inst.out_notouch_\[169\] cm_inst.cc_inst.out_notouch_\[177\]
+ cm_inst.cc_inst.out_notouch_\[185\] _048_ _023_ _077_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.buf_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_35_357 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_28_495 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_356 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_487 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_340 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_11_362 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_34_498 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_34_454 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.clkinv_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[197\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_2
XANTENNA_cm_inst.cc_inst.xnor2_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_44_229 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_338 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_32_45 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_25_443 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_432 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.nor2_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_40_393 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai32_2_inst_B1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_273 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_35_207 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_31_424 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_16_443 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.latsnq_1_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[29\].div_flop ro_inst.counter_n\[29\] in[0] ro_inst.counter_n\[28\]
+ ro_inst.counter\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_27_78 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_27_56 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_430 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_43_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai222_1_inst_C1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_273 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_402 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_17_229 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.or4_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.buf_3_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_3
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_15_Left_67 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.and4_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and4_2
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_51_477 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_51_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_16_295 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_42_411 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_485_ in[3] cm_inst.cc_inst.in\[1\] _240_ _007_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_27_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_254 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.bufz_16_inst_EN cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.aoi211_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[73\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_2
XFILLER_0_45_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_33_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__497__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__488__I1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_5_147 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.latq_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[124\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latq_2
XANTENNA__309__S _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_379 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_36_368 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_36_357 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_24_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_270_ cm_inst.cc_inst.out_notouch_\[192\] cm_inst.cc_inst.out_notouch_\[200\] _041_
+ _042_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
Xcm_inst.cc_inst.oai21_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[83\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_4
XANTENNA_cm_inst.cc_inst.dffsnq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_162 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_468_ _228_ _229_ _230_ _231_ ro_sel\[2\] ro_sel\[1\] _232_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.oai33_1_inst_B1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_19_249 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.inv_8_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_8
X_399_ _081_ _166_ _121_ _167_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_10_182 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_15_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_49_65 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.latrnq_2_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_2_128 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_18_Left_70 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SETN cm_inst.cc_inst.in\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nor3_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_322_ cm_inst.cc_inst.out_notouch_\[162\] cm_inst.cc_inst.out_notouch_\[170\] cm_inst.cc_inst.out_notouch_\[178\]
+ cm_inst.cc_inst.out_notouch_\[186\] _020_ _078_ _092_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XTAP_TAPCELL_ROW_24_285 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_24_349 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.dlyb_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[179\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyb_1
X_253_ cm_inst.cc_inst.out_notouch_\[96\] cm_inst.cc_inst.out_notouch_\[104\] cm_inst.cc_inst.out_notouch_\[112\]
+ cm_inst.cc_inst.out_notouch_\[120\] _021_ _024_ _025_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_32_371 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_27_187 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_23_393 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai221_2_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.sdffrsnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[167\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4
XFILLER_0_38_408 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_38_377 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_165 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_3_Left_55 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_14_382 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_474 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.oai221_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[99\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai221_1
XTAP_TAPCELL_ROW_12_200 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_305_ _075_ _076_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_37_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_32_190 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_21_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_35_358 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_43_455 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.xor3_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_430 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.icgtp_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[209\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__icgtp_4
XPHY_EDGE_ROW_45_Left_97 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_30_127 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_30_138 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.latrnq_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[127\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latrnq_2
XFILLER_0_19_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[19\].div_flop ro_inst.counter_n\[19\] in[0] ro_inst.counter_n\[18\]
+ ro_inst.counter\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XTAP_TAPCELL_ROW_40_394 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_37_293 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_271 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_339 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nor2_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.bufz_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[172\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_4
XANTENNA_cm_inst.cc_inst.oai32_2_inst_B2 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai32_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_48_450 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_43_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_411 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai221_4_inst_C cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_491 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.and2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_4
XTAP_TAPCELL_ROW_45_431 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai222_1_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai222_1_inst_C2 cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnq_2_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffsnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.or4_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_296 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.bufz_12_inst_EN cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_436 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_447 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[11\].div_flop_inv ro_inst.counter\[11\] ro_inst.counter_n\[11\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_40_255 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__420__S _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_21_480 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_48_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_51_478 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_8_463 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_16_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.latsnq_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[132\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latsnq_1
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.xor2_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_12_491 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_8_167 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.clkbuf_8_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__330__S _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_39_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_39_322 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_32_Left_84 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
X_484_ _238_ _240_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_ro_inst.gcount\[19\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_22_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_38_45 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_9_216 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_249 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_18_506 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.bufz_16_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[173\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_16
XANTENNA_cm_inst.cc_inst.latrsnq_1_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_5_148 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_36_303 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.oai33_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[93\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai33_1
XANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.oai33_1_inst_B2 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dffq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[148\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_2
X_398_ cm_inst.cc_inst.out_notouch_\[4\] cm_inst.cc_inst.out_notouch_\[12\] _119_
+ _166_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_467_ _210_ _224_ _225_ _231_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_380 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_10_183 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.latrnq_2_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_2_129 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_33_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.xnor2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[56\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor2_4
XANTENNA_cm_inst.cc_inst.nor3_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_321_ _091_ ro_inst.counter\[1\] _016_ out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_252_ _023_ _024_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.buf_20_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_20
XANTENNA__473__B in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_133 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_15_220 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_372 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai221_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai221_2_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.invz_8_inst_EN cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_38_378 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_114 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_37_431 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_304_ _032_ _075_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_201 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[5\].div_flop ro_inst.counter_n\[5\] in[0] ro_inst.counter_n\[4\]
+ ro_inst.counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_21_26 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.aoi221_4_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_47_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_359 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_43_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_43_467 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_43_434 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.xor3_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__502__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_34_478 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi221_4_inst_C cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_40_395 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_32_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai32_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_12_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_48_451 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_7_199 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_11_194 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_297 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[3\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_45_432 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai222_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai222_1_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.or4_2_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_51_479 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_51_468 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.aoi221_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[75\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi221_1
XANTENNA_cm_inst.cc_inst.xor2_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_453 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_442 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_31_278 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_256 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_8_168 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.aoi22_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[71\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_4
XANTENNA_cm_inst.cc_inst.clkinv_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_356 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_39_334 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_483_ in[2] cm_inst.cc_inst.in\[0\] _239_ _006_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_22_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SE cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dlyb_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_228 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xcm_inst.cc_inst.dlyd_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[186\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyd_2
XFILLER_0_13_201 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_13_267 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_278 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_5_149 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_44_370 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai33_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_1_inst_B3 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_42_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_39_175 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_39_164 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_397_ _083_ cm_inst.cc_inst.out_notouch_\[20\] _164_ _105_ _165_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi211_1
X_466_ _130_ _147_ ro_sel\[0\] _230_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XTAP_TAPCELL_ROW_10_184 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_10_259 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__426__S _133_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_18_240 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.invz_4_inst_EN cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_5_286 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_51_104 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_36_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_36_123 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
X_320_ _058_ _074_ _090_ _091_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor3_1
X_251_ _022_ _023_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_24_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nand3_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_15_221 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_449_ cm_inst.cc_inst.out_notouch_\[39\] cm_inst.cc_inst.out_notouch_\[47\] cm_inst.cc_inst.out_notouch_\[55\]
+ cm_inst.cc_inst.out_notouch_\[63\] _184_ _180_ _214_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_23_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_38_379 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai221_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_123 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_41_192 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.icgtp_4_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_37_476 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_303_ _059_ _073_ _074_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
XFILLER_0_32_170 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi221_4_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi221_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.xor3_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_11_398 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_38_229 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.addf_4_inst_CI cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_432 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_40_396 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_435 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_502 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.oai32_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_48_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_452 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nand2_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_4_inst_I cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_31_330 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_43_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_427 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.clkinv_12_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[201\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_12
XFILLER_0_22_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dffnrnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[139\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2
XFILLER_0_45_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.oai222_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_36_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_51_469 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_221 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_265 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_169 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__339__S _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai22_2_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_482_ _235_ _239_ _055_ _237_ _005_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
Xcm_inst.cc_inst.dlyb_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[181\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyb_4
XANTENNA_ro_inst.gcount\[32\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.inv_3_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.invz_8_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[175\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__invz_8
Xcm_inst.cc_inst.or3_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or3_2
XFILLER_0_13_257 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_21_290 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[28\].div_flop ro_inst.counter_n\[28\] in[0] ro_inst.counter_n\[27\]
+ ro_inst.counter\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_36_349 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_51_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_44_382 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.oai221_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[101\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai221_4
XANTENNA_cm_inst.cc_inst.oai33_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_465_ _172_ _189_ _225_ _229_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
Xcm_inst.cc_inst.nor3_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor3_1
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_35_360 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[20\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_327 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dffnsnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[144\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1
X_396_ _038_ cm_inst.cc_inst.out_notouch_\[28\] _164_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
XFILLER_0_49_57 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_185 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.nand3_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand3_1
XTAP_TAPCELL_ROW_18_241 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.mux2_4_inst_I0 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[29\].div_flop_inv ro_inst.counter\[29\] ro_inst.counter_n\[29\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XTAP_TAPCELL_ROW_1_120 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_51_138 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_36_179 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_250_ cm_inst.page\[1\] _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA_cm_inst.cc_inst.nand3_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_51_36 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_7_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_15_222 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_448_ _211_ _212_ _030_ _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_379_ ro_inst.enable _148_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_50_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_50_Left_102 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.mux4_1_inst_S0 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_157 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_258 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_29_314 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_302_ _067_ _072_ _033_ _073_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_37_444 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi221_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_333 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_344 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_499 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_28_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_11_344 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_366 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.dffrnq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_34_350 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_411 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_46_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.latsnq_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[134\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latsnq_4
XPHY_EDGE_ROW_7_Left_59 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_40_397 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_447 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_48_453 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nand2_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_222 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_200 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_31_331 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_28_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.aoi22_2_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.oai33_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[95\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai33_4
XFILLER_0_19_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_34_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_34_255 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_483 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_277 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_200 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA__270__S _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_23_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.oai22_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[84\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai22_1
Xro_inst.gcount\[18\].div_flop ro_inst.counter_n\[18\] in[0] ro_inst.counter_n\[17\]
+ ro_inst.counter\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_31_214 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_16_288 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_16_299 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_193 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_3_182 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai22_2_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_481_ _234_ _239_ _089_ _237_ _004_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XANTENNA_cm_inst.cc_inst.oai22_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_22_258 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_13_203 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_8_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.dlyc_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_36_Left_88 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.dffrnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_4_140 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_464_ _225_ _056_ _227_ _228_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XFILLER_0_42_309 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.mux4_2_inst_I0 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_199 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_35_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_395_ _158_ _160_ _045_ _162_ _163_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
XFILLER_0_49_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_49_25 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xcm_inst.cc_inst.dffrsnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[153\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1
XFILLER_0_10_228 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_10_186 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_18_242 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_45_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__505__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_339 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_5_277 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.mux2_4_inst_I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_1_121 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_36_103 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_32_375 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xcm_inst.cc_inst.sdffrnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[163\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2
XANTENNA_cm_inst.cc_inst.nand3_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_378_ _047_ _136_ _146_ _129_ _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
X_516_ out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tiel
X_447_ cm_inst.cc_inst.out_notouch_\[71\] cm_inst.cc_inst.out_notouch_\[79\] cm_inst.cc_inst.out_notouch_\[87\]
+ cm_inst.cc_inst.out_notouch_\[95\] _184_ _124_ _212_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_42_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_23_397 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_23_386 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_46_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_26_191 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.mux4_1_inst_S1 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_21_259 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_397 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_29_315 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_301_ _068_ _071_ _066_ _072_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XTAP_TAPCELL_ROW_37_370 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.dffq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_39_Left_91 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_43_459 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_434 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_401 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_23_Left_75 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_23_150 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.and3_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and3_1
XTAP_TAPCELL_ROW_34_351 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.aoi221_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[77\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi221_4
XFILLER_0_6_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_361 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_297 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai211_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.sdffsnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[168\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1
Xcm_inst.cc_inst.clkbuf_3_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[190\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_3
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.icgtn_1_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_ro_inst.gcount\[28\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_31_332 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_7_158 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_415 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.invz_1_inst_I cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_197 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[4\].div_flop ro_inst.counter_n\[4\] in[0] ro_inst.counter_n\[3\]
+ ro_inst.counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XANTENNA_cm_inst.cc_inst.aoi22_2_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi22_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_234 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_19_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_286 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_495 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.clkbuf_3_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[7\].div_flop_inv ro_inst.counter\[7\] ro_inst.counter_n\[7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_21_484 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[16\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_8_401 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_8_445 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_10_Left_62 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_12_495 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_42_405 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_326 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai22_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_480_ _233_ _239_ _173_ _237_ _003_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
Xcm_inst.cc_inst.clkinv_8_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[200\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_8
XFILLER_0_38_49 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.xnor3_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor3_1
Xro_inst.gcount\[32\].div_flop_inv ro_inst.counter\[32\] ro_inst.counter_n\[32\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XTAP_TAPCELL_ROW_7_160 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__319__A2 _080_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_44_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_36_307 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_381 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_286 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.and3_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_4_141 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_394_ _112_ _161_ _162_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
X_463_ _129_ _226_ _074_ _090_ _227_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or4_1
XANTENNA__366__S _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dffrnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[151\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_2
XANTENNA_cm_inst.cc_inst.mux4_2_inst_I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_340 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_10_187 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_18_243 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_5_201 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_41_398 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_41_343 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_289 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_1_122 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_44_181 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_24_279 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_515_ out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tiel
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_377_ _059_ _145_ _146_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
XANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_446_ cm_inst.cc_inst.out_notouch_\[103\] cm_inst.cc_inst.out_notouch_\[111\] cm_inst.cc_inst.out_notouch_\[119\]
+ cm_inst.cc_inst.out_notouch_\[127\] _184_ _180_ _211_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_35_170 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_23_376 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_14_310 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_18_137 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.tiel_inst cm_inst.cc_inst.out_notouch_\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tiel
XANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_316 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_300_ cm_inst.cc_inst.out_notouch_\[1\] cm_inst.cc_inst.out_notouch_\[9\] cm_inst.cc_inst.out_notouch_\[17\]
+ cm_inst.cc_inst.out_notouch_\[25\] _070_ _064_ _071_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_37_435 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_424 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_37_402 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_37_371 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.dffsnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[156\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffsnq_1
Xro_inst.gcount\[25\].div_flop_inv ro_inst.counter\[25\] ro_inst.counter_n\[25\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_20_335 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_43_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_429_ _103_ cm_inst.cc_inst.out_notouch_\[94\] _195_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
XANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_11_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.and4_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_34_352 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_6_373 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_40_Left_92 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai211_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.inv_12_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dffnrsnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[141\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1
XTAP_TAPCELL_ROW_31_333 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_28_221 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_31_419 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_16_449 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.latrsnq_1_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.aoi22_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi211_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_474 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.nor3_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor3_4
Xcm_inst.cc_inst.dffnsnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[146\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_25_235 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.nand3_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand3_4
XFILLER_0_21_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.inv_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_24_290 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_430 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_12_441 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_42_406 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_338 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_50_461 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_35_500 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xro_inst.gcount\[18\].div_flop_inv ro_inst.counter\[18\] ro_inst.counter_n\[18\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XTAP_TAPCELL_ROW_7_161 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SI cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_21_260 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_61 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_44_374 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_8_298 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_17_500 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.and3_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.xor2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[61\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor2_2
XTAP_TAPCELL_ROW_4_142 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_179 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_393_ cm_inst.cc_inst.out_notouch_\[100\] cm_inst.cc_inst.out_notouch_\[108\] cm_inst.cc_inst.out_notouch_\[116\]
+ cm_inst.cc_inst.out_notouch_\[124\] _085_ _113_ _161_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_27_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_462_ ro_sel\[0\] _226_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
XFILLER_0_50_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.mux4_2_inst_I2 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_1_123 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_363 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_514_ out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tiel
X_376_ _140_ _144_ _033_ _145_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_445_ _210_ ro_inst.counter\[34\] _148_ out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_23_333 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dlya_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[27\].div_flop ro_inst.counter_n\[27\] in[0] ro_inst.counter_n\[26\]
+ ro_inst.counter\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_25_95 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_25_51 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai31_1_inst_B cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.mux4_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[120\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_37_372 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_29_317 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_37_414 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_32_196 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_17_193 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_428_ _173_ _192_ _193_ _155_ _194_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XFILLER_0_7_319 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_417 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_359_ cm_inst.page\[5\] _129_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_23_152 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_51_494 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_11_336 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_358 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.oai22_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[86\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai22_4
XFILLER_0_36_61 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.and4_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_34_353 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_6_341 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_42_461 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_288 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_439 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_417 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_506 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_31_334 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_417 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_43_269 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.dlyc_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[182\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyc_1
XFILLER_0_24_461 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.latrsnq_1_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_11_144 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.aoi211_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_453 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_431 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_45_426 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__385__S _133_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_258 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_25_269 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dffrsnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[155\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.oai222_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[102\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai222_1
XFILLER_0_17_96 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_33_62 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA__508__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_3_inst_EN cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_225 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_3_174 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA__269__I _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_42_407 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_50_462 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_7_162 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.bufz_16_inst_I cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[3\].div_flop_inv ro_inst.counter\[3\] ro_inst.counter_n\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_21_272 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_73 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.dffsnq_2_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.and3_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_461_ ro_sel\[0\] _225_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XTAP_TAPCELL_ROW_4_143 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.mux4_2_inst_I3 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_39_158 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_35_364 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_35_342 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_23_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_392_ _107_ _159_ _031_ _160_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XANTENNA__493__I0 in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[17\].div_flop ro_inst.counter_n\[17\] in[0] ro_inst.counter_n\[16\]
+ ro_inst.counter\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_41_345 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_38_191 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_41 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_5_203 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_1_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__308__S0 _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_1_124 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xcm_inst.cc_inst.and3_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and3_4
XANTENNA_cm_inst.cc_inst.dffsnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrnq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_342 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_32_367 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__475__I0 in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_ro_inst.gcount\[8\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_444_ _018_ _194_ _209_ _058_ _210_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
X_513_ out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tiel
Xcm_inst.cc_inst.sdffsnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[170\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4
X_375_ _141_ _143_ _066_ _144_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA_cm_inst.cc_inst.icgtn_4_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_23_389 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_63 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.dffnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_29_318 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_37_373 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_37_437 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_32_131 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_20_251 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_32_164 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
X_427_ cm_inst.cc_inst.out_notouch_\[198\] cm_inst.cc_inst.out_notouch_\[206\] _039_
+ _193_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_358_ _116_ _127_ _017_ _128_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_1
XFILLER_0_36_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_289_ cm_inst.page\[0\] _060_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.and4_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_415 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_34_354 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_6_353 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_42_473 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or3_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_37_267 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_484 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__470__I in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.xnor3_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor3_4
XPHY_EDGE_ROW_27_Left_79 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xro_inst.gcount\[21\].div_flop_inv ro_inst.counter\[21\] ro_inst.counter_n\[21\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_43_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_204 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_ro_inst.slow_clock_inv_I in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.or2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[45\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or2_1
XFILLER_0_24_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_19_234 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__290__I cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_278 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_487 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_443 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_45_427 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.addf_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[105\] cm_inst.cc_inst.out_notouch_\[106\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu9t5v0__addf_1
XFILLER_0_25_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.latrnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_476 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_42 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_24_292 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_3_186 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_12_487 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_50_463 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_42_408 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_50_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_7_470 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_163 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.buf_16_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_16
XANTENNA_cm_inst.cc_inst.nor2_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[3\].div_flop ro_inst.counter_n\[3\] in[0] ro_inst.counter_n\[2\]
+ ro_inst.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XANTENNA_cm_inst.cc_inst.clkinv_20_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.icgtn_2_inst_TE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_44_332 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or4_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_14_Left_66 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_4_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_12_262 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_4_144 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__326__S1 _095_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_460_ _224_ ro_inst.saved_signal ro_inst.enable out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_391_ cm_inst.cc_inst.out_notouch_\[68\] cm_inst.cc_inst.out_notouch_\[76\] _108_
+ _159_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA_cm_inst.cc_inst.dffq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dffsnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[158\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffsnq_4
XFILLER_0_35_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.icgtp_4_inst_TE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_49_18 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[14\].div_flop_inv ro_inst.counter\[14\] ro_inst.counter_n\[14\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_41_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai222_4_inst_C1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_29_170 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.xnor3_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_374_ cm_inst.cc_inst.out_notouch_\[3\] cm_inst.cc_inst.out_notouch_\[11\] cm_inst.cc_inst.out_notouch_\[19\]
+ cm_inst.cc_inst.out_notouch_\[27\] _142_ _138_ _143_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_27_129 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_27_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_512_ _243_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tiel
X_443_ _201_ _208_ _059_ _209_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_1
XTAP_TAPCELL_ROW_15_216 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_368 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_23_335 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.aoi222_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[78\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi222_1
XFILLER_0_11_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.clkinv_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dffnrsnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[143\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4
XANTENNA__383__I _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_302 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_41_198 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_335 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_29_319 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_49_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_37_427 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_37_374 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_20_252 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_43_419 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_426_ _190_ _191_ _133_ _192_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_28_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_357_ _118_ _122_ _075_ _126_ _127_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
XANTENNA_cm_inst.cc_inst.oai33_4_inst_B1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_288_ cm_inst.page\[4\] _059_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_23_198 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_11_349 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.oai211_4_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_41 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_34_355 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.and4_1_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.inv_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_4
XFILLER_0_6_365 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.or3_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_37_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_37_246 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_ro_inst.gcount\[25\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_419 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_0_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_2_Left_54 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_48_447 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_409_ _174_ _175_ _133_ _176_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_24_441 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_44_Left_96 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.invz_1_inst cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[173\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__invz_1
XANTENNA_cm_inst.cc_inst.clkbuf_12_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_ro_inst.gcount\[13\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_45_428 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_290 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_260 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_10 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_8_449 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai32_1_inst_B1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_12_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_433 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_499 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__340__B _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_42_409 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_319 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_50_464 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.nor4_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_22_208 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_7_164 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__421__A2 _187_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nor2_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_5_419 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_21_274 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_44_366 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or4_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.mux4_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[122\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_4
XFILLER_0_29_385 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_4_145 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_390_ _102_ cm_inst.cc_inst.out_notouch_\[84\] _157_ _105_ _158_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi211_1
XPHY_EDGE_ROW_31_Left_83 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_5_216 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.oai222_4_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai222_4_inst_C2 cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_44_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_193 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_160 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.aoi21_1_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.xor2_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.xnor3_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_511_ _015_ in[0] ro_sel\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
X_373_ _069_ _142_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_442_ _203_ _205_ _034_ _207_ _208_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
XTAP_TAPCELL_ROW_23_272 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_15_217 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_31_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi211_4_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_76 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_10 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.dlyc_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[184\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyc_4
XFILLER_0_41_188 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai31_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_37_375 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_37_406 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.inv_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_32_133 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_32_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xcm_inst.cc_inst.or4_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or4_2
XTAP_TAPCELL_ROW_20_253 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.bufz_12_inst cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[172\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_12
XANTENNA_cm_inst.cc_inst.oai33_4_inst_B2 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_409 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.latsnq_4_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_425_ cm_inst.cc_inst.out_notouch_\[134\] cm_inst.cc_inst.out_notouch_\[142\] cm_inst.cc_inst.out_notouch_\[150\]
+ cm_inst.cc_inst.out_notouch_\[158\] _150_ _151_ _191_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_356_ _111_ _125_ _126_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
X_287_ cm_inst.page\[5\] _058_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_23_166 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xcm_inst.cc_inst.addh_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[113\]
+ cm_inst.cc_inst.out_notouch_\[114\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__addh_2
XANTENNA_cm_inst.cc_inst.oai211_4_inst_C cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.nor4_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor4_1
Xcm_inst.cc_inst.oai222_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[104\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai222_4
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai221_1_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnq_1_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.nand4_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand4_1
XANTENNA_cm_inst.cc_inst.or3_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[26\].div_flop ro_inst.counter_n\[26\] in[0] ro_inst.counter_n\[25\]
+ ro_inst.counter\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XTAP_TAPCELL_ROW_48_448 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.oai211_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[96\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
X_408_ cm_inst.cc_inst.out_notouch_\[133\] cm_inst.cc_inst.out_notouch_\[141\] cm_inst.cc_inst.out_notouch_\[149\]
+ cm_inst.cc_inst.out_notouch_\[157\] _119_ _151_ _175_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_339_ cm_inst.cc_inst.out_notouch_\[66\] cm_inst.cc_inst.out_notouch_\[74\] _108_
+ _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_11_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_37_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.latsnq_4_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_163 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_15_453 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_45_429 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_280 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.latrsnq_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[130\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latrsnq_2
XANTENNA_cm_inst.cc_inst.mux2_4_inst_S cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_17_88 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_16_217 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai32_1_inst_B2 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai32_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.icgtn_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[205\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__icgtn_2
XFILLER_0_24_272 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_412 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_12_445 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nor4_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_50_465 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_7_461 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_450 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_15_261 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_30_253 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_30_231 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_7_165 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_331 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.buf_16_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dlyd_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.or4_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA__487__I0 in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_356 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_345 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi222_2_inst_C1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_18_237 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_183 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_172 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_389 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_26_345 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai222_4_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai222_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_348 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_172 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_44_197 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.xor2_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_367 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_356 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.xnor3_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_441_ _111_ _206_ _207_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
X_510_ _014_ in[0] ro_sel\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
X_372_ cm_inst.cc_inst.out_notouch_\[35\] cm_inst.cc_inst.out_notouch_\[43\] cm_inst.cc_inst.out_notouch_\[51\]
+ cm_inst.cc_inst.out_notouch_\[59\] _070_ _064_ _141_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.latq_1_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_109 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_23_273 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_15_218 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.aoi211_4_inst_C cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_55 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xro_inst.gcount\[10\].div_flop_inv ro_inst.counter\[10\] ro_inst.counter_n\[10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA__303__A2 _073_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai31_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.or2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[47\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or2_4
XFILLER_0_22_381 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_37_376 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_37_418 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[16\].div_flop ro_inst.counter_n\[16\] in[0] ro_inst.counter_n\[15\]
+ ro_inst.counter\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_17_197 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_20_254 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_424_ cm_inst.cc_inst.out_notouch_\[166\] cm_inst.cc_inst.out_notouch_\[174\] cm_inst.cc_inst.out_notouch_\[182\]
+ cm_inst.cc_inst.out_notouch_\[190\] _150_ _095_ _190_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
Xcm_inst.cc_inst.addf_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[109\] cm_inst.cc_inst.out_notouch_\[110\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu9t5v0__addf_4
XFILLER_0_28_418 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_28_310 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai33_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_4_inst_B3 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_51_410 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_36_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_355_ cm_inst.cc_inst.out_notouch_\[34\] cm_inst.cc_inst.out_notouch_\[42\] cm_inst.cc_inst.out_notouch_\[50\]
+ cm_inst.cc_inst.out_notouch_\[58\] _123_ _124_ _125_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_286_ _016_ _056_ _057_ out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XANTENNA_cm_inst.cc_inst.dffrnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_54 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.addh_4_inst_A cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_407 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_42_465 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai221_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai221_1_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_18_440 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_20_115 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_48_449 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_407_ cm_inst.cc_inst.out_notouch_\[165\] cm_inst.cc_inst.out_notouch_\[173\] cm_inst.cc_inst.out_notouch_\[181\]
+ cm_inst.cc_inst.out_notouch_\[189\] _150_ _151_ _174_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_28_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_338_ _060_ _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_51_240 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_24_465 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_269_ _020_ _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.clkinv_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[196\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.latsnq_4_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_435 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.latrsnq_4_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_10_181 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_502 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_424 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_44_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai32_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffsnq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_3_189 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.clkinv_8_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nor4_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_50_466 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_15_273 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.buf_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_2
XTAP_TAPCELL_ROW_7_166 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.and4_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and4_1
XTAP_TAPCELL_ROW_41_400 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.aoi222_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[80\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi222_4
XFILLER_0_41_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.or4_1_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nand2_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_376 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA__487__I1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.aoi211_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[72\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
XANTENNA_cm_inst.cc_inst.icgtn_2_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_390 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.invz_2_inst_I cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__496__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_23_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.aoi222_2_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_2_inst_C2 cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.latq_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[123\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latq_1
XTAP_TAPCELL_ROW_18_238 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_26_293 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai222_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_ro_inst.gcount\[5\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SE cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_49_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.clkbuf_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_324 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[2\].div_flop ro_inst.counter_n\[2\] in[0] ro_inst.counter_n\[1\]
+ ro_inst.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
X_371_ _137_ _139_ _066_ _140_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_440_ cm_inst.cc_inst.out_notouch_\[38\] cm_inst.cc_inst.out_notouch_\[46\] cm_inst.cc_inst.out_notouch_\[54\]
+ cm_inst.cc_inst.out_notouch_\[62\] _123_ _113_ _206_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XTAP_TAPCELL_ROW_15_219 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.latq_1_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_176 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_110 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_274 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__511__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_12 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_25_78 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_25_67 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_143 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_1_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai31_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.invz_3_inst_EN cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__357__B _075_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.invz_4_inst cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[174\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__invz_4
XTAP_TAPCELL_ROW_20_255 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_13_360 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_28_311 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_354_ _063_ _124_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_423_ _189_ ro_inst.counter\[5\] _148_ out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA_cm_inst.cc_inst.oai33_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_51_444 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_285_ ro_inst.counter\[0\] ro_inst.enable _057_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XFILLER_0_23_135 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_3_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_36_99 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.addh_4_inst_B cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_290 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai221_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_357 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_419 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_6_379 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_205 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_33_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_208 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.latrnq_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[126\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latrnq_1
XTAP_TAPCELL_ROW_31_328 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_24_400 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_406_ _075_ _173_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_337_ _098_ _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_51_274 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_268_ _037_ _039_ _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_19_205 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_238 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.mux4_4_inst_S0 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_403 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.bufz_3_inst cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[171\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_3
XANTENNA_cm_inst.cc_inst.sdffq_2_inst_SE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_6_Left_58 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_18_271 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_44_420 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai32_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_50_467 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nor4_2_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_7_463 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nand4_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_41_401 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_26_506 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_28_45 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_44_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_322 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.nand2_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_238 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_44_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_44_336 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_336 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_43_380 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.inv_20_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_20
XANTENNA_cm_inst.cc_inst.aoi222_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.latrsnq_2_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_2_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai22_1_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_163 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_294 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_9_Left_61 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_18_239 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_41_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_38_174 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_39_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.nor4_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor4_4
XTAP_TAPCELL_ROW_1_118 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_130 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.dffq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[147\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XFILLER_0_17_336 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.nand4_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand4_4
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_370_ cm_inst.cc_inst.out_notouch_\[67\] cm_inst.cc_inst.out_notouch_\[75\] cm_inst.cc_inst.out_notouch_\[83\]
+ cm_inst.cc_inst.out_notouch_\[91\] _070_ _138_ _139_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XPHY_EDGE_ROW_35_Left_87 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_23_275 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.oai211_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[98\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_4
XANTENNA_ro_inst.gcount\[34\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_499_ _003_ in[0] cm_inst.page\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XFILLER_0_26_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_41_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_14_306 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_333 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_45_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_17_100 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_199 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_20_256 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.sig_cmp ro_inst.signal ro_inst.saved_signal ro_inst.running vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__xnor2_1
XTAP_TAPCELL_ROW_28_312 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_353_ _069_ _123_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_422_ _018_ _178_ _188_ _058_ _189_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
X_284_ _018_ _035_ _054_ _055_ _056_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
XFILLER_0_51_478 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_ro_inst.gcount\[22\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.xor3_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[64\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor3_2
XFILLER_0_36_56 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_27_442 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_169 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__501__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_31_329 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_24_445 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_24_423 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_405_ _172_ ro_inst.counter\[4\] _148_ out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_267_ _038_ _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XANTENNA_ro_inst.gcount\[10\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai21_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_336_ _102_ cm_inst.cc_inst.out_notouch_\[82\] _104_ _105_ _106_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi211_1
XFILLER_0_22_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_38_Left_90 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_47_440 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_47_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_22_Left_74 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.mux4_4_inst_S1 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_155 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.dlya_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_10_161 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[28\].div_flop_inv ro_inst.counter\[28\] ro_inst.counter_n\[28\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
Xro_inst.slow_clock_inv in[0] ro_inst.slow_clk_n vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SE cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai31_2_inst_B cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_294 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.addf_1_inst_A cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_33_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_17_58 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_421 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_46 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_24_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_253 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_12_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_12_437 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.clkbuf_20_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[195\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_20
XFILLER_0_16_209 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_319_ _076_ _080_ _088_ _089_ _090_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
Xro_inst.gcount\[25\].div_flop ro_inst.counter_n\[25\] in[0] ro_inst.counter_n\[24\]
+ ro_inst.counter\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_7_442 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.aoi22_1_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_7_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_15_231 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nand4_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_402 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.latrnq_4_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_256 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_389 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_378 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_345 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_356 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_4_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.oai31_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[88\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai31_2
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.dlyd_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[185\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyd_1
XFILLER_0_7_272 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.latrsnq_2_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai22_1_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai22_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.latrsnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_26_295 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__305__I _075_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_1_119 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_44_189 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_370 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_40_395 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_48_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_35_134 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_31_362 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_23_276 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dffnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[136\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnq_2
XFILLER_0_16_392 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_395 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_25_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.mux4_1_inst_I0 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_498_ _002_ in[0] cm_inst.page\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XFILLER_0_26_189 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_123 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_26_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_210 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.clkinv_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[199\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_4
XFILLER_0_22_373 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_189 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_20_257 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_28_313 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_421_ _059_ _187_ _188_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
XANTENNA_cm_inst.cc_inst.aoi21_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_454 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_36_443 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_352_ _081_ _120_ _121_ _122_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
X_283_ cm_inst.page\[5\] _055_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
XFILLER_0_36_46 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_349 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_39_292 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__368__S1 _064_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_10_376 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_181 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_SE cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_37_207 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_33_413 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_18_432 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_424 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.and4_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and4_4
Xro_inst.ring_osc_0 ro_inst.ring\[0\] ro_inst.enable ro_inst.ring\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
X_404_ _018_ _156_ _171_ _129_ _172_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
XANTENNA_cm_inst.cc_inst.invz_8_inst_I cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_295 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_36_240 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_266_ _019_ _038_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA_cm_inst.cc_inst.oai21_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_335_ _036_ _105_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xro_inst.gcount\[15\].div_flop ro_inst.counter_n\[15\] in[0] ro_inst.counter_n\[14\]
+ ro_inst.counter\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XTAP_TAPCELL_ROW_47_441 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_27_240 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_30_427 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_173 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.aoi211_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[74\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_4
XANTENNA_cm_inst.cc_inst.addf_1_inst_B cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__499__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.and2_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.latq_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[125\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latq_4
Xcm_inst.cc_inst.tieh_inst cm_inst.cc_inst.out_notouch_\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tieh
XANTENNA_cm_inst.cc_inst.oai211_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_44_422 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_318_ cm_inst.page\[4\] _089_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
X_249_ _020_ _021_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_12_449 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dffnrnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[138\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1
XFILLER_0_47_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_35_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_7_454 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.and4_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_202 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.aoi22_1_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi22_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_265 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nand4_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_41_403 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_26_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.dffrnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.latrnq_4_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_139 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_393 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_43_360 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__392__B _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.or3_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or3_1
XANTENNA_cm_inst.cc_inst.oai22_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_187 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_296 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_1_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_17_230 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_382 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_ro_inst.gcount\[18\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.and3_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__406__I _075_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_23_277 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xcm_inst.cc_inst.latrnq_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[128\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latrnq_4
XANTENNA_cm_inst.cc_inst.mux4_1_inst_I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_14_211 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_497_ _001_ in[0] cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XFILLER_0_6_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xro_inst.gcount\[6\].div_flop_inv ro_inst.counter\[6\] ro_inst.counter_n\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_22_341 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_17_146 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_32_127 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_31_80 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi21_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_420_ _182_ _186_ _033_ _187_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_351_ _044_ _121_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_36_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_282_ _043_ _046_ _047_ _053_ _054_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
Xro_inst.gcount\[31\].div_flop_inv ro_inst.counter\[31\] ro_inst.counter_n\[31\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_27_444 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xro_inst.gcount\[1\].div_flop ro_inst.counter_n\[1\] in[0] ro_inst.counter_n\[0\]
+ ro_inst.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_42_469 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffsnq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_349 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_193 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_444 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_41_480 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.ring_osc_1 ro_inst.ring\[1\] ro_inst.ring\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
X_403_ _163_ _170_ _017_ _171_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_1
X_334_ _103_ cm_inst.cc_inst.out_notouch_\[90\] _104_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
XFILLER_0_36_263 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_265_ _036_ _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XTAP_TAPCELL_ROW_47_442 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_27_296 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_233 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_439 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.clkinv_3_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_506 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_18_263 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.dlyb_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_44_423 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.and2_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai211_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_317_ _084_ _087_ _046_ _088_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_1
XFILLER_0_24_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.sdffq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__324__I _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_248_ _019_ _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_20_461 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dffq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[149\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_4
XANTENNA_cm_inst.cc_inst.and4_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_7_466 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_277 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi22_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.nand4_2_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_41_404 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_236 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[24\].div_flop_inv ro_inst.counter\[24\] ro_inst.counter_n\[24\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.icgtp_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_44_306 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_29_347 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_20_291 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[2\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai21_1_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_372 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_38_155 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_297 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SI cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_166 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_144 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_17_231 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_17_328 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_40_397 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_494 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_110 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__322__S0 _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__504__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.and3_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_23_278 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_16_361 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_31_364 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_496_ _000_ in[0] cm_inst.page\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XTAP_TAPCELL_ROW_14_212 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.mux4_1_inst_I2 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[34\].div_flop ro_inst.counter_n\[34\] in[0] ro_inst.counter_n\[33\]
+ ro_inst.counter\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_10_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_49_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.sdffrnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[162\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1
XFILLER_0_9_347 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_342 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_350_ cm_inst.cc_inst.out_notouch_\[2\] cm_inst.cc_inst.out_notouch_\[10\] _119_
+ _120_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_36_423 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xro_inst.gcount\[17\].div_flop_inv ro_inst.counter\[17\] ro_inst.counter_n\[17\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_281_ _034_ _052_ _053_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
X_479_ _238_ _239_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_10_378 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_18_423 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.aoi21_2_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_264_ cm_inst.page\[1\] _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
X_402_ _165_ _167_ _034_ _169_ _170_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
Xro_inst.ring_osc_2 ro_inst.ring\[2\] ro_inst.ring\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
X_333_ _093_ _103_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_24_437 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_404 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_47_443 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_209 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_30_321 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_286 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffq_2_inst_SI cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.clkbuf_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[189\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_2
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffsnq_1_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dlyd_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[187\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyd_4
XFILLER_0_18_275 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_44_424 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_247_ cm_inst.page\[0\] _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XPHY_EDGE_ROW_26_Left_78 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_24_201 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_316_ _037_ _086_ _087_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XANTENNA__281__A1 _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.and4_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__451__S _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__250__I cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_46_381 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_29_326 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_44_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_195 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.bufz_2_inst_EN cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_93 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_28_370 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_31_502 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xro_inst.gcount\[24\].div_flop ro_inst.counter_n\[24\] in[0] ro_inst.counter_n\[23\]
+ ro_inst.counter\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_38_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_26_298 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.buf_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.latrnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dffrnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[150\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XTAP_TAPCELL_ROW_17_232 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_40_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_29_Left_81 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_25_362 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_234 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_ro_inst.gcount\[31\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_92 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_13_Left_65 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_0_111 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_35_126 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xcm_inst.cc_inst.buf_8_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_8
XFILLER_0_31_310 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.and3_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_31_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or2_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.mux4_1_inst_I3 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_39_390 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_495_ in[4] ro_sel\[2\] _242_ _015_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XTAP_TAPCELL_ROW_14_213 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_22_332 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xcm_inst.cc_inst.buf_12_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_12
XANTENNA_cm_inst.cc_inst.or4_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dlyd_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_280_ _049_ _050_ _051_ _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_39_295 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_39_273 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_478_ in[1] _238_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_6_307 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_368 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xcm_inst.cc_inst.dffnrnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[140\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4
Xro_inst.gcount\[2\].div_flop_inv ro_inst.counter\[2\] ro_inst.counter_n\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_45_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_33_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_401_ _111_ _168_ _169_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XFILLER_0_36_232 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_24_427 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
X_263_ _025_ _026_ _027_ _028_ _031_ _034_ _035_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_332_ _082_ _102_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_47_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_47_444 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.latq_2_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__338__I _060_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_419 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_322 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_10_165 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_81 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_33_202 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SI cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.or3_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or3_4
XANTENNA_cm_inst.cc_inst.or3_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_298 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_44_425 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_1_Left_53 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
X_315_ cm_inst.cc_inst.out_notouch_\[193\] cm_inst.cc_inst.out_notouch_\[201\] _085_
+ _086_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_24_268 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_257 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_246_ _017_ _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XTAP_TAPCELL_ROW_9_180 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_7_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.and4_4_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_11_441 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_43_Left_95 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xro_inst.gcount\[14\].div_flop ro_inst.counter_n\[14\] in[0] ro_inst.counter_n\[13\]
+ ro_inst.counter\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_14_290 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.xnor2_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_12_196 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_221 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_102 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_26_299 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_382 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.xor2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[60\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor2_1
XFILLER_0_9_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_17_233 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[20\].div_flop_inv ro_inst.counter\[20\] ro_inst.counter_n\[20\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.oai32_4_inst_B1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_4_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.icgtn_1_inst_TE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_0_112 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_396 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.or2_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_12_inst_I cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
X_494_ in[3] ro_sel\[1\] _242_ _014_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XTAP_TAPCELL_ROW_14_214 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_34_193 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_30_Left_82 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_22_377 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_9_349 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.or4_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_149 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_48_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_36_447 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_36_403 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.xnor3_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai221_1_inst_C cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.invz_3_inst_I cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_477_ in[4] _112_ _236_ _002_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_10_303 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_342 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_SI cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_436 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_447 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_5_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_400_ cm_inst.cc_inst.out_notouch_\[36\] cm_inst.cc_inst.out_notouch_\[44\] cm_inst.cc_inst.out_notouch_\[52\]
+ cm_inst.cc_inst.out_notouch_\[60\] _123_ _124_ _168_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_331_ _076_ _097_ _099_ _100_ _101_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XFILLER_0_36_299 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_36_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_262_ _033_ _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_24_406 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.nor3_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.aoi21_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[67\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_2
XTAP_TAPCELL_ROW_47_445 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[13\].div_flop_inv ro_inst.counter\[13\] ro_inst.counter_n\[13\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.latq_2_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SETN cm_inst.cc_inst.in\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_30_323 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_155 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__264__I cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.or3_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_277 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_314_ _019_ _085_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_245_ cm_inst.page\[4\] _017_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_24_203 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__349__I _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_23_62 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.oai221_4_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_11_453 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_3_61 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__507__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_ro_inst.gcount\[27\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.xnor2_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_40_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_197 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.sdffrnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[164\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4
XFILLER_0_20_272 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_283 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_47_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_43_364 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_501 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.nor4_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_3_132 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_169 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_ro_inst.gcount\[15\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_22_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_17_234 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_40_312 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai32_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai32_4_inst_B2 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__483__I0 in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_113 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_48_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_16_353 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi221_1_inst_C cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_493_ in[2] _225_ _242_ _013_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
Xcm_inst.cc_inst.hold_inst cm_inst.cc_inst.out_notouch_\[173\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__hold
XFILLER_0_39_456 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_215 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_191 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_22_270 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_1_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_15_96 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or4_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_31_84 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_334 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_356 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.mux2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[118\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_2
XTAP_TAPCELL_ROW_28_307 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.xnor3_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_120 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_16_161 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_476_ in[3] _107_ _236_ _001_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_50_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_26_73 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_33_343 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_41_484 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai31_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_197 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[33\].div_flop ro_inst.counter_n\[33\] in[0] ro_inst.counter_n\[32\]
+ ro_inst.counter\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
X_330_ cm_inst.cc_inst.out_notouch_\[194\] cm_inst.cc_inst.out_notouch_\[202\] _041_
+ _100_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_261_ _032_ _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XANTENNA_cm_inst.cc_inst.nor3_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_47_446 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_30_324 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_459_ _058_ _218_ _223_ _224_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor3_1
XFILLER_0_6_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_42_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.dlya_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[177\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlya_2
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_37_83 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.inv_16_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_16
XANTENNA_cm_inst.cc_inst.or3_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_244_ ro_inst.enable _016_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
X_313_ _081_ _083_ cm_inst.cc_inst.out_notouch_\[209\] _084_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand3_1
XANTENNA__391__S _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_465 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dffrnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[152\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_4
XFILLER_0_7_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_7_415 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai221_4_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai221_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.xor3_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_270 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_21_207 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__386__S _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xro_inst.clock_gate ro_inst.ring\[0\] ro_inst.running _243_ ro_inst.counter\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__icgtp_2
XTAP_TAPCELL_ROW_12_198 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_41 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_376 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nor4_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_104 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_3_133 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_17_235 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.addf_2_inst_A cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_25_290 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_343 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_25_332 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_4_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_4_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai32_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_51 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_31_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA__483__I1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_0_114 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_48_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_16_343 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnq_4_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_492_ in[5] in[6] in[7] in[1] _242_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand4_1
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.aoi222_1_inst_C1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_22_271 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_10_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.sdffq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[160\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffq_2
XFILLER_0_45_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_38_490 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or4_4_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_1_inst_I cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_17_Left_69 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.invz_12_inst cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[175\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__invz_12
XFILLER_0_13_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[23\].div_flop ro_inst.counter_n\[23\] in[0] ro_inst.counter_n\[22\]
+ ro_inst.counter\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_36_363 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_28_308 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.xnor3_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_395 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_31_132 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.clkbuf_16_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[194\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_16
XFILLER_0_39_243 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.oai32_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[91\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai32_2
X_475_ in[2] _039_ _237_ _000_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA__455__S0 _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_2_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SE cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.inv_20_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_33_344 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai31_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_427 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_260_ cm_inst.page\[3\] _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
Xcm_inst.cc_inst.inv_3_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_3
XFILLER_0_8_192 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nor3_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_30_325 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_458_ _173_ _221_ _222_ _155_ _089_ _223_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi221_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_389_ _103_ cm_inst.cc_inst.out_notouch_\[92\] _157_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
XFILLER_0_23_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_23_430 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__284__A2 _035_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.clkinv_16_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_5_195 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_441 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_500 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_312_ _082_ _083_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XANTENNA__471__I in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.xor2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[62\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor2_4
XANTENNA_cm_inst.cc_inst.aoi221_2_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai221_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.xor3_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_11_433 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_500 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XPHY_EDGE_ROW_5_Left_57 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_6_153 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_199 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_20_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.dffsnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_374 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_47_Left_99 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_43_388 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_506 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_268 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nor4_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_3_134 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_19_341 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_25_291 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_17_236 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.addf_2_inst_B cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_366 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai32_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[13\].div_flop ro_inst.counter_n\[13\] in[0] ro_inst.counter_n\[12\]
+ ro_inst.counter\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_104 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_0_115 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_196 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_358 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xro_inst.sig_latch ro_inst.signal ro_inst.slow_clk_n ro_inst.saved_signal vdd vdd
+ vss vss gf180mcu_fd_sc_mcu9t5v0__latq_1
XANTENNA_cm_inst.cc_inst.buf_12_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_458 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_491_ _241_ _012_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.aoi222_1_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_1_inst_C2 cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_174 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_22_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_22_369 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_8_Left_60 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_25_196 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_28_309 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_36_364 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_12_380 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_34_Left_86 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.oai22_4_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_277 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_39_233 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_474_ _236_ _237_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_27_428 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.or4_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or4_1
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_33_345 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_ro_inst.gcount\[7\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_33_409 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai31_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_453 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.invz_2_inst_EN cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_144 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.addh_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[111\]
+ cm_inst.cc_inst.out_notouch_\[112\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__addh_1
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_51_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_44_280 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_32_464 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.nand3_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_30_326 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_203 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_23_442 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_388_ _076_ _153_ _154_ _155_ _156_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
X_457_ _102_ cm_inst.cc_inst.out_notouch_\[199\] _222_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
XFILLER_0_10_169 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_37_63 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.dlyc_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_453 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_311_ _048_ _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
XANTENNA_cm_inst.cc_inst.aoi221_2_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi221_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_509_ _013_ in[0] ro_sel\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XFILLER_0_11_412 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_21_Left_73 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.xor3_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.latrsnq_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[129\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latrsnq_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_3_20 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_11_445 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_309 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffq_1_inst_SE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_461 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.addf_2_inst_CI cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_294 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.icgtn_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[204\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__icgtn_1
XFILLER_0_21_209 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_6_154 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__495__I0 in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_7_214 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_43_356 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_11_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.clkbuf_8_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[192\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_8
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__486__I0 in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nor4_1_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_3_135 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_34_301 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_386 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.nand4_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__477__I0 in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.clkinv_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_25_292 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_378 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.dffq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_0_105 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_0_116 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_17_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_28_183 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_389 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_3_250 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi22_4_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_39_384 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_490_ _238_ _016_ _236_ _241_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XANTENNA_cm_inst.cc_inst.aoi222_1_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_183 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_197 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.clock_gate_inv ro_inst.counter\[0\] ro_inst.counter_n\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_15_88 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_31_65 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_429 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_36_407 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_36_365 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_29_481 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_44_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_31_178 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_375 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.oai22_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai22_4_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_223 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_473_ _233_ _234_ _235_ in[1] _236_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai31_1
XANTENNA_cm_inst.cc_inst.oai21_2_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_10_307 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.nor2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[37\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_2
XTAP_TAPCELL_ROW_33_346 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_429 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_41_476 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_41_410 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.mux2_2_inst_I0 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.nand2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_2
XFILLER_0_8_194 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xro_inst.gcount\[9\].div_flop_inv ro_inst.counter\[9\] ro_inst.counter_n\[9\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.mux4_4_inst_I0 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nand3_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_456_ _219_ _220_ _121_ _221_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_35_270 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_30_327 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_248 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_387_ _099_ _155_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_37_20 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_419 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_310_ _078_ _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XANTENNA__291__S0 _060_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_32_251 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xro_inst.gcount\[34\].div_flop_inv ro_inst.counter\[34\] ro_inst.counter_n\[34\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_174 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.invz_12_inst_I cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi221_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai21_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_ro_inst.gcount\[24\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[32\].div_flop ro_inst.counter_n\[32\] in[0] ro_inst.counter_n\[31\]
+ ro_inst.counter\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
X_508_ _012_ in[0] ro_inst.enable vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
X_439_ _081_ _204_ _121_ _205_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XFILLER_0_23_251 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_6_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_262 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SE cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_6_155 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_40_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.buf_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_18_77 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_20_287 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_65 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[12\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_368 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_28_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_11_190 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA__486__I1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_3_136 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_49_Left_101 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.nand4_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_379 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_22_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.oai211_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_324 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_13_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_10 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__442__B _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_98 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_106 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_0_117 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_357 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.oai21_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[82\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_2
XANTENNA_cm_inst.cc_inst.aoi22_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi22_4_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_405 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_39_385 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[27\].div_flop_inv ro_inst.counter\[27\] ro_inst.counter_n\[27\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.aoi222_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_195 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.latrsnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_338 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA__510__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_36_366 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_471 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA__302__S _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai22_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_472_ in[7] _235_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
XTAP_TAPCELL_ROW_27_300 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.invz_3_inst cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[174\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__invz_3
Xcm_inst.cc_inst.sdffrsnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[166\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2
XTAP_TAPCELL_ROW_33_347 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_41_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.buf_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_463 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.mux2_2_inst_I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_44_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_44_271 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_430 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.and3_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi21_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.mux4_4_inst_I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[22\].div_flop ro_inst.counter_n\[22\] in[0] ro_inst.counter_n\[21\]
+ ro_inst.counter\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XANTENNA_cm_inst.cc_inst.nand3_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.clkbuf_20_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_386_ cm_inst.cc_inst.out_notouch_\[196\] cm_inst.cc_inst.out_notouch_\[204\] _041_
+ _154_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_455_ cm_inst.cc_inst.out_notouch_\[135\] cm_inst.cc_inst.out_notouch_\[143\] cm_inst.cc_inst.out_notouch_\[151\]
+ cm_inst.cc_inst.out_notouch_\[159\] _108_ _098_ _220_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_50_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.icgtp_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[208\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__icgtp_2
XFILLER_0_26_271 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_SE cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__291__S1 _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_482 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.bufz_2_inst cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[171\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_2
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_9_175 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_20_436 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai21_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_369_ _063_ _138_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_438_ cm_inst.cc_inst.out_notouch_\[6\] cm_inst.cc_inst.out_notouch_\[14\] _119_
+ _204_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_507_ _011_ in[0] cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XFILLER_0_7_419 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_46_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_34_506 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_14_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_14_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_6_156 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.and2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_2
XFILLER_0_9_290 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.and2_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_45 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_43_347 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_191 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_11_266 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_3_137 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_42_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nand4_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai211_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.or4_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or4_4
XFILLER_0_25_358 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_336 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_88 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_107 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_303 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_369 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xcm_inst.cc_inst.addh_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[115\]
+ cm_inst.cc_inst.out_notouch_\[116\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__addh_4
XANTENNA_cm_inst.cc_inst.aoi22_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_39_386 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_14_209 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_34_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_30_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffrnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_22_328 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_450 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_494 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_36_367 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.xnor2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[55\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor2_2
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_29_450 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_399 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_372 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_27_301 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.invz_12_inst_EN cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_203 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_471_ in[6] _234_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
Xro_inst.gcount\[12\].div_flop ro_inst.counter_n\[12\] in[0] ro_inst.counter_n\[11\]
+ ro_inst.counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_50_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SI cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_45_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_348 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.latrsnq_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[131\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latrsnq_4
Xcm_inst.cc_inst.xor3_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor3_1
XANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_36_228 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.icgtn_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[206\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__icgtn_4
XFILLER_0_8_141 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.clkinv_20_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[203\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_20
XANTENNA_cm_inst.cc_inst.and3_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_12_191 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi21_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.mux4_4_inst_I2 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_454_ cm_inst.cc_inst.out_notouch_\[167\] cm_inst.cc_inst.out_notouch_\[175\] cm_inst.cc_inst.out_notouch_\[183\]
+ cm_inst.cc_inst.out_notouch_\[191\] _108_ _098_ _219_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_385_ _149_ _152_ _133_ _153_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA__500__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_23_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_23_434 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_10_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_37_88 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_37_77 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_37_55 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_14_401 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_445 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_32_297 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_17_261 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_9_176 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_506_ _010_ in[0] cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XFILLER_0_23_46 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_368_ cm_inst.cc_inst.out_notouch_\[99\] cm_inst.cc_inst.out_notouch_\[107\] cm_inst.cc_inst.out_notouch_\[115\]
+ cm_inst.cc_inst.out_notouch_\[123\] _070_ _064_ _137_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_299_ _069_ _070_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_15_209 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xro_inst.gcount\[5\].div_flop_inv ro_inst.counter\[5\] ro_inst.counter_n\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
X_437_ _083_ cm_inst.cc_inst.out_notouch_\[22\] _202_ _105_ _203_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi211_1
XFILLER_0_23_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_11_437 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.icgtn_4_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai221_2_inst_C cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.invz_4_inst_I cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_464 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA__489__I0 in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_6_157 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.and2_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_256 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_25_Left_77 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xro_inst.gcount\[30\].div_flop_inv ro_inst.counter\[30\] ro_inst.counter_n\[30\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_34_45 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_217 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_378 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_11_201 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_11_192 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.aoi22_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[70\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_2
XTAP_TAPCELL_ROW_3_138 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.aoi211_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_261 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_345 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_378 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nand4_1_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_37_120 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xcm_inst.cc_inst.oai31_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[87\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai31_1
XFILLER_0_33_370 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_67 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_108 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_24_392 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_370 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_3_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_39_387 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[9\].div_flop ro_inst.counter_n\[9\] in[0] ro_inst.counter_n\[8\]
+ ro_inst.counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_22_265 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_30_395 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_318 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xcm_inst.cc_inst.dffnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[135\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnq_1
XFILLER_0_21_373 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_36_368 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_28_Left_80 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_8_323 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_12_Left_64 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_16_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.clkinv_3_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[198\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_3
XFILLER_0_12_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_ro_inst.gcount\[4\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_27_302 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_470_ in[5] _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xro_inst.gcount\[23\].div_flop_inv ro_inst.counter\[23\] ro_inst.counter_n\[23\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA__300__S1 _064_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_41_402 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_465 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_41_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_49_460 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_17_410 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_44_273 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_32_435 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.and3_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.mux4_4_inst_I3 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_453_ _047_ _217_ _218_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
X_384_ cm_inst.cc_inst.out_notouch_\[132\] cm_inst.cc_inst.out_notouch_\[140\] cm_inst.cc_inst.out_notouch_\[148\]
+ cm_inst.cc_inst.out_notouch_\[156\] _150_ _151_ _152_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA__294__S0 _060_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_35_295 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.buf_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_4
XFILLER_0_23_446 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.aoi221_2_inst_C cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_37_67 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_46_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.icgtn_2_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_273 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_9_177 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_505_ _009_ in[0] cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
X_436_ _103_ cm_inst.cc_inst.out_notouch_\[30\] _202_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
XFILLER_0_43_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_298_ cm_inst.page\[0\] _069_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XANTENNA__498__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_367_ _076_ _134_ _135_ _099_ _136_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XFILLER_0_23_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_449 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__409__S _133_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffq_1_inst_SI cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.latrsnq_4_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_298 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__489__I1 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_6_158 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xro_inst.gcount\[16\].div_flop_inv ro_inst.counter\[16\] ro_inst.counter_n\[16\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XPHY_EDGE_ROW_0_Left_52 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_20_268 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_419_ _183_ _185_ _030_ _186_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_7_207 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_11_193 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.buf_8_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi211_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_305 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_42_371 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_42_Left_94 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xro_inst.gcount\[31\].div_flop ro_inst.counter_n\[31\] in[0] ro_inst.counter_n\[30\]
+ ro_inst.counter\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XANTENNA_cm_inst.cc_inst.or3_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dlyb_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[180\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyb_2
XANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_500 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_109 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai211_1_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_187 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_24_382 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.bufz_1_inst_EN cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_39_388 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.oai221_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[100\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai221_2
XFILLER_0_19_132 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_34_168 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_34_135 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_187 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_22_266 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_30_363 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_31_14 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_25_146 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_36_369 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_430 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_8_302 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_485 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_16_157 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_80 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_39_216 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_27_303 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__327__S _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffsnq_4_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.or2_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.icgtp_2_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_293 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.dlya_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.icgtn_4_inst_TE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai31_4_inst_B cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_260 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_44_285 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_44_263 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_ro_inst.gcount\[33\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_383_ _061_ _151_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA__294__S1 _064_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_452_ _213_ _216_ _075_ _217_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_23_458 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.latsnq_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[133\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latsnq_2
XFILLER_0_41_233 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_ro_inst.gcount\[21\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_2_inst_I cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.xnor3_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_9_178 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_43_412 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_504_ _008_ in[0] cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
X_435_ _196_ _198_ _045_ _200_ _201_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
X_366_ cm_inst.cc_inst.out_notouch_\[195\] cm_inst.cc_inst.out_notouch_\[203\] _041_
+ _135_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_297_ cm_inst.cc_inst.out_notouch_\[33\] cm_inst.cc_inst.out_notouch_\[41\] cm_inst.cc_inst.out_notouch_\[49\]
+ cm_inst.cc_inst.out_notouch_\[57\] _060_ _061_ _068_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_11_406 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_3_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.oai33_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[94\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai33_2
XANTENNA_cm_inst.cc_inst.latrsnq_4_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_222 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[21\].div_flop ro_inst.counter_n\[21\] in[0] ro_inst.counter_n\[20\]
+ ro_inst.counter\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_14_233 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_14_255 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_14_266 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_159 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SI cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi211_1_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_339 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
X_349_ _093_ _119_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_28_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_303 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_418_ cm_inst.cc_inst.out_notouch_\[5\] cm_inst.cc_inst.out_notouch_\[13\] cm_inst.cc_inst.out_notouch_\[21\]
+ cm_inst.cc_inst.out_notouch_\[29\] _184_ _180_ _185_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_36_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_11_194 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[1\].div_flop_inv ro_inst.counter\[1\] ro_inst.counter_n\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XTAP_TAPCELL_ROW_19_250 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_42_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.inv_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.or3_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_339 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_286 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_14 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.xnor2_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.oai211_1_inst_C cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.xor3_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[65\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor3_4
XTAP_TAPCELL_ROW_39_389 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_47_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_19_144 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_19_199 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_267 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_30_353 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_30_375 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_38_420 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_442 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__503__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_25_125 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_40_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_180 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nor2_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_375 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_475 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_29_442 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_44_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.latsnq_1_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SETN cm_inst.cc_inst.in\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_31_128 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_39_239 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_39_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_27_304 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nor4_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_194 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or2_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.icgtp_2_inst_TE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_22_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.mux2_1_inst_S cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_434 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai222_2_inst_C1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_32_340 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_17_434 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_382_ _093_ _150_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_451_ _214_ _215_ _051_ _216_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_35_297 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_35_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_23_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_37_14 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.aoi221_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[76\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi221_2
XFILLER_0_41_278 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_275 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_437 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[11\].div_flop ro_inst.counter_n\[11\] in[0] ro_inst.counter_n\[10\]
+ ro_inst.counter\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_SI cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.xnor3_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_286 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_32_267 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_191 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_9_179 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.clkbuf_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[188\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_503_ _007_ in[0] cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XANTENNA_cm_inst.cc_inst.nor3_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_43_413 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.oai31_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[89\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai31_4
X_296_ _062_ _065_ _066_ _067_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_434_ _112_ _199_ _200_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XFILLER_0_28_507 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_365_ _131_ _132_ _133_ _134_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai33_2_inst_B1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai31_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.latsnq_2_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_9_261 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.aoi211_1_inst_C cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
X_417_ _069_ _184_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
X_348_ _083_ cm_inst.cc_inst.out_notouch_\[18\] _117_ _036_ _118_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi211_1
Xcm_inst.cc_inst.dffnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[137\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnq_4
X_279_ _044_ _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_19_337 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.or3_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_220 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA__492__A1 in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_2_130 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.inv_12_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_12
XTAP_TAPCELL_ROW_25_287 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.dlyc_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_370 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.xnor2_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_123 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xro_inst.gcount\[12\].div_flop_inv ro_inst.counter\[12\] ro_inst.counter_n\[12\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_16_307 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.addh_1_inst_A cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_24_362 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_351 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_34_137 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_22_268 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_454 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_13_202 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_38_498 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[29\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_31_49 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_25_148 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_33_192 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nor2_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.latsnq_1_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_304 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_398 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.nor4_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_35_360 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_27_305 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__297__S0 _060_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_ro_inst.gcount\[17\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_34_490 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.oai222_2_inst_C2 cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai222_2_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__333__I _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_16_Left_68 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xro_inst.gcount\[8\].div_flop ro_inst.counter_n\[8\] in[0] ro_inst.counter_n\[7\]
+ ro_inst.counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_44_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_32_341 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_17_402 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_12_195 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.xor2_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_381_ cm_inst.cc_inst.out_notouch_\[164\] cm_inst.cc_inst.out_notouch_\[172\] cm_inst.cc_inst.out_notouch_\[180\]
+ cm_inst.cc_inst.out_notouch_\[188\] _094_ _095_ _149_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_450_ cm_inst.cc_inst.out_notouch_\[7\] cm_inst.cc_inst.out_notouch_\[15\] cm_inst.cc_inst.out_notouch_\[23\]
+ cm_inst.cc_inst.out_notouch_\[31\] _123_ _124_ _215_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_23_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi222_4_inst_C1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_46_433 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__328__I _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_202 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_405 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_14_449 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_49_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_37_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.xnor3_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_243 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_17_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_40_290 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_43_414 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_433_ cm_inst.cc_inst.out_notouch_\[102\] cm_inst.cc_inst.out_notouch_\[110\] cm_inst.cc_inst.out_notouch_\[118\]
+ cm_inst.cc_inst.out_notouch_\[126\] _085_ _113_ _199_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_502_ _006_ in[0] cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XANTENNA_cm_inst.cc_inst.nor3_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_51_480 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_295_ _029_ _066_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_364_ _044_ _133_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA_cm_inst.cc_inst.oai33_2_inst_B2 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_31_290 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.clkbuf_12_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[193\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_12
XANTENNA_cm_inst.cc_inst.clkbuf_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.oai31_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.nor3_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor3_2
XPHY_EDGE_ROW_19_Left_71 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.dffnsnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[145\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2
XFILLER_0_9_240 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_227 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.nand3_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand3_2
XTAP_TAPCELL_ROW_5_150 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_34_49 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_416_ cm_inst.cc_inst.out_notouch_\[37\] cm_inst.cc_inst.out_notouch_\[45\] cm_inst.cc_inst.out_notouch_\[53\]
+ cm_inst.cc_inst.out_notouch_\[61\] _142_ _138_ _183_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_36_371 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_278_ cm_inst.cc_inst.out_notouch_\[128\] cm_inst.cc_inst.out_notouch_\[136\] cm_inst.cc_inst.out_notouch_\[144\]
+ cm_inst.cc_inst.out_notouch_\[152\] _048_ _023_ _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_11_205 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_347_ _038_ cm_inst.cc_inst.out_notouch_\[26\] _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
XFILLER_0_24_93 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.xor3_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_349 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_30_503 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_6_265 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__452__S _075_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__492__A2 in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_2_131 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_4_Left_56 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_25_288 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.bufz_8_inst cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[172\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_8
XFILLER_0_18_382 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_16 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_8_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.addh_1_inst_B cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_396 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_374 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_24_341 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.latrsnq_2_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_3_246 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_503 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_46_Left_98 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_34_127 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_15_341 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_124 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_269 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_30_399 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_322 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.bufz_8_inst_I cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_396 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_400 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_38_380 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_ro_inst.gcount\[1\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_13_203 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_127 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_29_411 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xro_inst.gcount\[30\].div_flop ro_inst.counter_n\[30\] in[0] ro_inst.counter_n\[29\]
+ ro_inst.counter\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_29_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_327 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_12_333 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_27_306 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nor4_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_219 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_35_361 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.aoi21_4_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_447 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_360 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__297__S1 _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_406 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai222_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai222_2_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.xor2_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_12_163 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_380_ _147_ ro_inst.counter\[3\] _148_ out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA_cm_inst.cc_inst.aoi222_4_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_4_inst_C2 cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_33_Left_85 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.oai22_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[85\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai22_2
XTAP_TAPCELL_ROW_46_434 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_26_222 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffrnq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__280__S _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.aoi21_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[66\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_1
.ends

