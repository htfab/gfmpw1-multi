magic
tech gf180mcuD
magscale 1 5
timestamp 1702448219
<< obsm1 >>
rect 672 1971 19400 18189
<< metal2 >>
rect 7392 19600 7448 20000
rect 7728 19600 7784 20000
<< obsm2 >>
rect 2030 19570 7362 19600
rect 7478 19570 7698 19600
rect 7814 19570 19386 19600
rect 2030 1997 19386 19570
<< metal3 >>
rect 19600 12768 20000 12824
rect 19600 12432 20000 12488
rect 0 12096 400 12152
rect 19600 12096 20000 12152
rect 0 11760 400 11816
rect 19600 11760 20000 11816
rect 0 11424 400 11480
rect 19600 11424 20000 11480
rect 0 11088 400 11144
rect 19600 11088 20000 11144
rect 0 10752 400 10808
rect 19600 10752 20000 10808
rect 0 10416 400 10472
rect 19600 10416 20000 10472
rect 0 10080 400 10136
rect 19600 10080 20000 10136
rect 0 9744 400 9800
rect 19600 9744 20000 9800
rect 0 9408 400 9464
rect 19600 9408 20000 9464
rect 0 9072 400 9128
rect 19600 9072 20000 9128
rect 0 8736 400 8792
rect 19600 8736 20000 8792
rect 0 8400 400 8456
rect 19600 8400 20000 8456
rect 0 8064 400 8120
rect 19600 8064 20000 8120
rect 19600 7728 20000 7784
rect 19600 7392 20000 7448
<< obsm3 >>
rect 400 12854 19600 18158
rect 400 12738 19570 12854
rect 400 12518 19600 12738
rect 400 12402 19570 12518
rect 400 12182 19600 12402
rect 430 12066 19570 12182
rect 400 11846 19600 12066
rect 430 11730 19570 11846
rect 400 11510 19600 11730
rect 430 11394 19570 11510
rect 400 11174 19600 11394
rect 430 11058 19570 11174
rect 400 10838 19600 11058
rect 430 10722 19570 10838
rect 400 10502 19600 10722
rect 430 10386 19570 10502
rect 400 10166 19600 10386
rect 430 10050 19570 10166
rect 400 9830 19600 10050
rect 430 9714 19570 9830
rect 400 9494 19600 9714
rect 430 9378 19570 9494
rect 400 9158 19600 9378
rect 430 9042 19570 9158
rect 400 8822 19600 9042
rect 430 8706 19570 8822
rect 400 8486 19600 8706
rect 430 8370 19570 8486
rect 400 8150 19600 8370
rect 430 8034 19570 8150
rect 400 7814 19600 8034
rect 400 7698 19570 7814
rect 400 7478 19600 7698
rect 400 7362 19570 7478
rect 400 2002 19600 7362
<< metal4 >>
rect 2923 1986 3083 18174
rect 5254 1986 5414 18174
rect 7585 1986 7745 18174
rect 9916 1986 10076 18174
rect 12247 1986 12407 18174
rect 14578 1986 14738 18174
rect 16909 1986 17069 18174
rect 19240 1986 19400 18174
<< labels >>
rlabel metal2 s 7392 19600 7448 20000 6 clk
port 1 nsew signal input
rlabel metal3 s 0 8064 400 8120 6 in[0]
port 2 nsew signal input
rlabel metal3 s 19600 7392 20000 7448 6 in[10]
port 3 nsew signal input
rlabel metal3 s 19600 12768 20000 12824 6 in[11]
port 4 nsew signal input
rlabel metal3 s 19600 8400 20000 8456 6 in[12]
port 5 nsew signal input
rlabel metal3 s 19600 8736 20000 8792 6 in[13]
port 6 nsew signal input
rlabel metal3 s 19600 9408 20000 9464 6 in[14]
port 7 nsew signal input
rlabel metal3 s 19600 8064 20000 8120 6 in[15]
port 8 nsew signal input
rlabel metal3 s 19600 9744 20000 9800 6 in[16]
port 9 nsew signal input
rlabel metal3 s 19600 10080 20000 10136 6 in[17]
port 10 nsew signal input
rlabel metal3 s 0 9744 400 9800 6 in[1]
port 11 nsew signal input
rlabel metal3 s 0 12096 400 12152 6 in[2]
port 12 nsew signal input
rlabel metal3 s 0 9072 400 9128 6 in[3]
port 13 nsew signal input
rlabel metal3 s 0 8400 400 8456 6 in[4]
port 14 nsew signal input
rlabel metal3 s 0 10080 400 10136 6 in[5]
port 15 nsew signal input
rlabel metal3 s 0 8736 400 8792 6 in[6]
port 16 nsew signal input
rlabel metal3 s 0 11424 400 11480 6 in[7]
port 17 nsew signal input
rlabel metal3 s 0 11760 400 11816 6 in[8]
port 18 nsew signal input
rlabel metal3 s 0 11088 400 11144 6 in[9]
port 19 nsew signal input
rlabel metal2 s 7728 19600 7784 20000 6 out[0]
port 20 nsew signal output
rlabel metal3 s 19600 9072 20000 9128 6 out[10]
port 21 nsew signal output
rlabel metal3 s 19600 11760 20000 11816 6 out[11]
port 22 nsew signal output
rlabel metal3 s 0 10752 400 10808 6 out[1]
port 23 nsew signal output
rlabel metal3 s 0 10416 400 10472 6 out[2]
port 24 nsew signal output
rlabel metal3 s 19600 12096 20000 12152 6 out[3]
port 25 nsew signal output
rlabel metal3 s 19600 11088 20000 11144 6 out[4]
port 26 nsew signal output
rlabel metal3 s 19600 11424 20000 11480 6 out[5]
port 27 nsew signal output
rlabel metal3 s 19600 7728 20000 7784 6 out[6]
port 28 nsew signal output
rlabel metal3 s 19600 12432 20000 12488 6 out[7]
port 29 nsew signal output
rlabel metal3 s 19600 10752 20000 10808 6 out[8]
port 30 nsew signal output
rlabel metal3 s 19600 10416 20000 10472 6 out[9]
port 31 nsew signal output
rlabel metal3 s 0 9408 400 9464 6 rst_n
port 32 nsew signal input
rlabel metal4 s 2923 1986 3083 18174 6 vdd
port 33 nsew power bidirectional
rlabel metal4 s 7585 1986 7745 18174 6 vdd
port 33 nsew power bidirectional
rlabel metal4 s 12247 1986 12407 18174 6 vdd
port 33 nsew power bidirectional
rlabel metal4 s 16909 1986 17069 18174 6 vdd
port 33 nsew power bidirectional
rlabel metal4 s 5254 1986 5414 18174 6 vss
port 34 nsew ground bidirectional
rlabel metal4 s 9916 1986 10076 18174 6 vss
port 34 nsew ground bidirectional
rlabel metal4 s 14578 1986 14738 18174 6 vss
port 34 nsew ground bidirectional
rlabel metal4 s 19240 1986 19400 18174 6 vss
port 34 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 280892
string GDS_FILE /home/htamas/progs/gfmpw1-multi.v3/openlane/loopback9/runs/23_12_13_07_15/results/signoff/loopback9.magic.gds
string GDS_START 75428
<< end >>

