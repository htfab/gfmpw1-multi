VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO input_mux
  CLASS BLOCK ;
  FOREIGN input_mux ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 4.000 ;
    END
  END clk
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 196.000 14.000 200.000 ;
    END
  END in[0]
  PIN in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 0.000 27.440 4.000 ;
    END
  END in[10]
  PIN in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 0.000 40.880 4.000 ;
    END
  END in[11]
  PIN in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END in[12]
  PIN in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 0.000 47.600 4.000 ;
    END
  END in[13]
  PIN in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END in[14]
  PIN in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END in[15]
  PIN in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END in[16]
  PIN in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 196.000 74.480 200.000 ;
    END
  END in[17]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 196.000 30.800 200.000 ;
    END
  END in[1]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 196.000 34.160 200.000 ;
    END
  END in[2]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 196.000 20.720 200.000 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 196.000 47.600 200.000 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 196.000 27.440 200.000 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.440 4.000 98.000 ;
    END
  END in[7]
  PIN in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END in[8]
  PIN in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END in[9]
  PIN proj_clk[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END proj_clk[0]
  PIN proj_clk[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END proj_clk[1]
  PIN proj_clk[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END proj_clk[2]
  PIN proj_clk[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 0.000 155.120 4.000 ;
    END
  END proj_clk[3]
  PIN proj_clk[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 4.000 ;
    END
  END proj_clk[4]
  PIN proj_clk[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 0.000 148.400 4.000 ;
    END
  END proj_clk[5]
  PIN proj_clk[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END proj_clk[6]
  PIN proj_clk[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END proj_clk[7]
  PIN proj_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 196.000 182.000 200.000 ;
    END
  END proj_in[0]
  PIN proj_in[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 16.800 200.000 17.360 ;
    END
  END proj_in[100]
  PIN proj_in[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 36.960 200.000 37.520 ;
    END
  END proj_in[101]
  PIN proj_in[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 77.280 200.000 77.840 ;
    END
  END proj_in[102]
  PIN proj_in[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 4.000 ;
    END
  END proj_in[103]
  PIN proj_in[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 0.000 128.240 4.000 ;
    END
  END proj_in[104]
  PIN proj_in[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 0.000 121.520 4.000 ;
    END
  END proj_in[105]
  PIN proj_in[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 26.880 200.000 27.440 ;
    END
  END proj_in[106]
  PIN proj_in[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 196.000 114.800 200.000 ;
    END
  END proj_in[107]
  PIN proj_in[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 196.000 81.200 200.000 ;
    END
  END proj_in[108]
  PIN proj_in[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 196.000 175.280 200.000 ;
    END
  END proj_in[109]
  PIN proj_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 40.320 200.000 40.880 ;
    END
  END proj_in[10]
  PIN proj_in[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 196.000 91.280 200.000 ;
    END
  END proj_in[110]
  PIN proj_in[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 196.000 87.920 200.000 ;
    END
  END proj_in[111]
  PIN proj_in[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 196.000 101.360 200.000 ;
    END
  END proj_in[112]
  PIN proj_in[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 196.000 94.640 200.000 ;
    END
  END proj_in[113]
  PIN proj_in[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 196.000 171.920 200.000 ;
    END
  END proj_in[114]
  PIN proj_in[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 196.000 104.720 200.000 ;
    END
  END proj_in[115]
  PIN proj_in[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END proj_in[116]
  PIN proj_in[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END proj_in[117]
  PIN proj_in[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END proj_in[118]
  PIN proj_in[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 4.000 ;
    END
  END proj_in[119]
  PIN proj_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 47.040 200.000 47.600 ;
    END
  END proj_in[11]
  PIN proj_in[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END proj_in[120]
  PIN proj_in[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 4.000 ;
    END
  END proj_in[121]
  PIN proj_in[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 4.000 ;
    END
  END proj_in[122]
  PIN proj_in[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 4.000 ;
    END
  END proj_in[123]
  PIN proj_in[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 4.000 ;
    END
  END proj_in[124]
  PIN proj_in[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 196.000 84.560 200.000 ;
    END
  END proj_in[125]
  PIN proj_in[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 196.000 155.120 200.000 ;
    END
  END proj_in[126]
  PIN proj_in[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 196.000 134.960 200.000 ;
    END
  END proj_in[127]
  PIN proj_in[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 196.000 148.400 200.000 ;
    END
  END proj_in[128]
  PIN proj_in[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 196.000 145.040 200.000 ;
    END
  END proj_in[129]
  PIN proj_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 53.760 200.000 54.320 ;
    END
  END proj_in[12]
  PIN proj_in[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 178.080 200.000 178.640 ;
    END
  END proj_in[130]
  PIN proj_in[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 147.840 200.000 148.400 ;
    END
  END proj_in[131]
  PIN proj_in[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 124.320 200.000 124.880 ;
    END
  END proj_in[132]
  PIN proj_in[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 104.160 200.000 104.720 ;
    END
  END proj_in[133]
  PIN proj_in[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 94.080 200.000 94.640 ;
    END
  END proj_in[134]
  PIN proj_in[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 33.600 200.000 34.160 ;
    END
  END proj_in[135]
  PIN proj_in[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 43.680 200.000 44.240 ;
    END
  END proj_in[136]
  PIN proj_in[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 80.640 200.000 81.200 ;
    END
  END proj_in[137]
  PIN proj_in[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 70.560 200.000 71.120 ;
    END
  END proj_in[138]
  PIN proj_in[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 4.000 ;
    END
  END proj_in[139]
  PIN proj_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 60.480 200.000 61.040 ;
    END
  END proj_in[13]
  PIN proj_in[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END proj_in[140]
  PIN proj_in[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 0.000 134.960 4.000 ;
    END
  END proj_in[141]
  PIN proj_in[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 174.720 200.000 175.280 ;
    END
  END proj_in[142]
  PIN proj_in[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 157.920 200.000 158.480 ;
    END
  END proj_in[143]
  PIN proj_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 0.000 141.680 4.000 ;
    END
  END proj_in[14]
  PIN proj_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 0.000 138.320 4.000 ;
    END
  END proj_in[15]
  PIN proj_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 161.280 200.000 161.840 ;
    END
  END proj_in[16]
  PIN proj_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 131.040 200.000 131.600 ;
    END
  END proj_in[17]
  PIN proj_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 196.000 37.520 200.000 ;
    END
  END proj_in[18]
  PIN proj_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 196.000 17.360 200.000 ;
    END
  END proj_in[19]
  PIN proj_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 196.000 111.440 200.000 ;
    END
  END proj_in[1]
  PIN proj_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 196.000 54.320 200.000 ;
    END
  END proj_in[20]
  PIN proj_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 196.000 61.040 200.000 ;
    END
  END proj_in[21]
  PIN proj_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END proj_in[22]
  PIN proj_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END proj_in[23]
  PIN proj_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.840 4.000 148.400 ;
    END
  END proj_in[24]
  PIN proj_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.280 4.000 161.840 ;
    END
  END proj_in[25]
  PIN proj_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END proj_in[26]
  PIN proj_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.960 4.000 37.520 ;
    END
  END proj_in[27]
  PIN proj_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.320 4.000 40.880 ;
    END
  END proj_in[28]
  PIN proj_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 4.000 54.320 ;
    END
  END proj_in[29]
  PIN proj_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 196.000 121.520 200.000 ;
    END
  END proj_in[2]
  PIN proj_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.560 4.000 71.120 ;
    END
  END proj_in[30]
  PIN proj_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 4.000 ;
    END
  END proj_in[31]
  PIN proj_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END proj_in[32]
  PIN proj_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 4.000 ;
    END
  END proj_in[33]
  PIN proj_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END proj_in[34]
  PIN proj_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END proj_in[35]
  PIN proj_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 4.000 131.600 ;
    END
  END proj_in[36]
  PIN proj_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END proj_in[37]
  PIN proj_in[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 196.000 57.680 200.000 ;
    END
  END proj_in[38]
  PIN proj_in[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 4.000 138.320 ;
    END
  END proj_in[39]
  PIN proj_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 196.000 168.560 200.000 ;
    END
  END proj_in[3]
  PIN proj_in[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END proj_in[40]
  PIN proj_in[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END proj_in[41]
  PIN proj_in[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END proj_in[42]
  PIN proj_in[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END proj_in[43]
  PIN proj_in[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 4.000 57.680 ;
    END
  END proj_in[44]
  PIN proj_in[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.280 4.000 77.840 ;
    END
  END proj_in[45]
  PIN proj_in[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END proj_in[46]
  PIN proj_in[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.040 4.000 47.600 ;
    END
  END proj_in[47]
  PIN proj_in[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 63.840 4.000 64.400 ;
    END
  END proj_in[48]
  PIN proj_in[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 4.000 44.240 ;
    END
  END proj_in[49]
  PIN proj_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 120.960 200.000 121.520 ;
    END
  END proj_in[4]
  PIN proj_in[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.400 4.000 50.960 ;
    END
  END proj_in[50]
  PIN proj_in[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 67.200 4.000 67.760 ;
    END
  END proj_in[51]
  PIN proj_in[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 196.000 178.640 200.000 ;
    END
  END proj_in[52]
  PIN proj_in[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 196.000 98.000 200.000 ;
    END
  END proj_in[53]
  PIN proj_in[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 196.000 24.080 200.000 ;
    END
  END proj_in[54]
  PIN proj_in[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 196.000 44.240 200.000 ;
    END
  END proj_in[55]
  PIN proj_in[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 196.000 71.120 200.000 ;
    END
  END proj_in[56]
  PIN proj_in[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 196.000 40.880 200.000 ;
    END
  END proj_in[57]
  PIN proj_in[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.520 4.000 108.080 ;
    END
  END proj_in[58]
  PIN proj_in[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 4.000 158.480 ;
    END
  END proj_in[59]
  PIN proj_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 154.560 200.000 155.120 ;
    END
  END proj_in[5]
  PIN proj_in[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 4.000 104.720 ;
    END
  END proj_in[60]
  PIN proj_in[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END proj_in[61]
  PIN proj_in[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.640 4.000 81.200 ;
    END
  END proj_in[62]
  PIN proj_in[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 4.000 84.560 ;
    END
  END proj_in[63]
  PIN proj_in[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 73.920 4.000 74.480 ;
    END
  END proj_in[64]
  PIN proj_in[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 4.000 61.040 ;
    END
  END proj_in[65]
  PIN proj_in[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END proj_in[66]
  PIN proj_in[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 0.000 67.760 4.000 ;
    END
  END proj_in[67]
  PIN proj_in[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 4.000 ;
    END
  END proj_in[68]
  PIN proj_in[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END proj_in[69]
  PIN proj_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 168.000 200.000 168.560 ;
    END
  END proj_in[6]
  PIN proj_in[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 4.000 145.040 ;
    END
  END proj_in[70]
  PIN proj_in[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END proj_in[71]
  PIN proj_in[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 196.000 131.600 200.000 ;
    END
  END proj_in[72]
  PIN proj_in[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 196.000 128.240 200.000 ;
    END
  END proj_in[73]
  PIN proj_in[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 196.000 138.320 200.000 ;
    END
  END proj_in[74]
  PIN proj_in[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 196.000 141.680 200.000 ;
    END
  END proj_in[75]
  PIN proj_in[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 134.400 200.000 134.960 ;
    END
  END proj_in[76]
  PIN proj_in[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 114.240 200.000 114.800 ;
    END
  END proj_in[77]
  PIN proj_in[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 110.880 200.000 111.440 ;
    END
  END proj_in[78]
  PIN proj_in[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 100.800 200.000 101.360 ;
    END
  END proj_in[79]
  PIN proj_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 107.520 200.000 108.080 ;
    END
  END proj_in[7]
  PIN proj_in[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 20.160 200.000 20.720 ;
    END
  END proj_in[80]
  PIN proj_in[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 30.240 200.000 30.800 ;
    END
  END proj_in[81]
  PIN proj_in[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 84.000 200.000 84.560 ;
    END
  END proj_in[82]
  PIN proj_in[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 50.400 200.000 50.960 ;
    END
  END proj_in[83]
  PIN proj_in[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 73.920 200.000 74.480 ;
    END
  END proj_in[84]
  PIN proj_in[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 63.840 200.000 64.400 ;
    END
  END proj_in[85]
  PIN proj_in[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 67.200 200.000 67.760 ;
    END
  END proj_in[86]
  PIN proj_in[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 57.120 200.000 57.680 ;
    END
  END proj_in[87]
  PIN proj_in[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 144.480 200.000 145.040 ;
    END
  END proj_in[88]
  PIN proj_in[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 127.680 200.000 128.240 ;
    END
  END proj_in[89]
  PIN proj_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 23.520 200.000 24.080 ;
    END
  END proj_in[8]
  PIN proj_in[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 196.000 118.160 200.000 ;
    END
  END proj_in[90]
  PIN proj_in[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 196.000 161.840 200.000 ;
    END
  END proj_in[91]
  PIN proj_in[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 196.000 165.200 200.000 ;
    END
  END proj_in[92]
  PIN proj_in[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 196.000 124.880 200.000 ;
    END
  END proj_in[93]
  PIN proj_in[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 137.760 200.000 138.320 ;
    END
  END proj_in[94]
  PIN proj_in[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 117.600 200.000 118.160 ;
    END
  END proj_in[95]
  PIN proj_in[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 164.640 200.000 165.200 ;
    END
  END proj_in[96]
  PIN proj_in[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 171.360 200.000 171.920 ;
    END
  END proj_in[97]
  PIN proj_in[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 97.440 200.000 98.000 ;
    END
  END proj_in[98]
  PIN proj_in[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 87.360 200.000 87.920 ;
    END
  END proj_in[99]
  PIN proj_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 90.720 200.000 91.280 ;
    END
  END proj_in[9]
  PIN proj_rst_n[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 196.000 151.760 200.000 ;
    END
  END proj_rst_n[0]
  PIN proj_rst_n[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 196.000 64.400 200.000 ;
    END
  END proj_rst_n[1]
  PIN proj_rst_n[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 196.000 158.480 200.000 ;
    END
  END proj_rst_n[2]
  PIN proj_rst_n[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 196.000 67.760 200.000 ;
    END
  END proj_rst_n[3]
  PIN proj_rst_n[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 141.120 200.000 141.680 ;
    END
  END proj_rst_n[4]
  PIN proj_rst_n[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 196.000 108.080 200.000 ;
    END
  END proj_rst_n[5]
  PIN proj_rst_n[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 196.000 50.960 200.000 ;
    END
  END proj_rst_n[6]
  PIN proj_rst_n[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 151.200 200.000 151.760 ;
    END
  END proj_rst_n[7]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 196.000 77.840 200.000 ;
    END
  END rst_n
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 0.000 108.080 4.000 ;
    END
  END sel[0]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END sel[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 29.230 15.380 30.830 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 75.850 15.380 77.450 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.470 15.380 124.070 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 169.090 15.380 170.690 184.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 52.540 15.380 54.140 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.160 15.380 100.760 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 145.780 15.380 147.380 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 192.400 15.380 194.000 184.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 4.630 194.000 189.130 ;
      LAYER Metal2 ;
        RECT 8.540 195.700 13.140 196.000 ;
        RECT 14.300 195.700 16.500 196.000 ;
        RECT 17.660 195.700 19.860 196.000 ;
        RECT 21.020 195.700 23.220 196.000 ;
        RECT 24.380 195.700 26.580 196.000 ;
        RECT 27.740 195.700 29.940 196.000 ;
        RECT 31.100 195.700 33.300 196.000 ;
        RECT 34.460 195.700 36.660 196.000 ;
        RECT 37.820 195.700 40.020 196.000 ;
        RECT 41.180 195.700 43.380 196.000 ;
        RECT 44.540 195.700 46.740 196.000 ;
        RECT 47.900 195.700 50.100 196.000 ;
        RECT 51.260 195.700 53.460 196.000 ;
        RECT 54.620 195.700 56.820 196.000 ;
        RECT 57.980 195.700 60.180 196.000 ;
        RECT 61.340 195.700 63.540 196.000 ;
        RECT 64.700 195.700 66.900 196.000 ;
        RECT 68.060 195.700 70.260 196.000 ;
        RECT 71.420 195.700 73.620 196.000 ;
        RECT 74.780 195.700 76.980 196.000 ;
        RECT 78.140 195.700 80.340 196.000 ;
        RECT 81.500 195.700 83.700 196.000 ;
        RECT 84.860 195.700 87.060 196.000 ;
        RECT 88.220 195.700 90.420 196.000 ;
        RECT 91.580 195.700 93.780 196.000 ;
        RECT 94.940 195.700 97.140 196.000 ;
        RECT 98.300 195.700 100.500 196.000 ;
        RECT 101.660 195.700 103.860 196.000 ;
        RECT 105.020 195.700 107.220 196.000 ;
        RECT 108.380 195.700 110.580 196.000 ;
        RECT 111.740 195.700 113.940 196.000 ;
        RECT 115.100 195.700 117.300 196.000 ;
        RECT 118.460 195.700 120.660 196.000 ;
        RECT 121.820 195.700 124.020 196.000 ;
        RECT 125.180 195.700 127.380 196.000 ;
        RECT 128.540 195.700 130.740 196.000 ;
        RECT 131.900 195.700 134.100 196.000 ;
        RECT 135.260 195.700 137.460 196.000 ;
        RECT 138.620 195.700 140.820 196.000 ;
        RECT 141.980 195.700 144.180 196.000 ;
        RECT 145.340 195.700 147.540 196.000 ;
        RECT 148.700 195.700 150.900 196.000 ;
        RECT 152.060 195.700 154.260 196.000 ;
        RECT 155.420 195.700 157.620 196.000 ;
        RECT 158.780 195.700 160.980 196.000 ;
        RECT 162.140 195.700 164.340 196.000 ;
        RECT 165.500 195.700 167.700 196.000 ;
        RECT 168.860 195.700 171.060 196.000 ;
        RECT 172.220 195.700 174.420 196.000 ;
        RECT 175.580 195.700 177.780 196.000 ;
        RECT 178.940 195.700 181.140 196.000 ;
        RECT 182.300 195.700 193.860 196.000 ;
        RECT 8.540 4.300 193.860 195.700 ;
        RECT 8.540 4.000 26.580 4.300 ;
        RECT 27.740 4.000 29.940 4.300 ;
        RECT 31.100 4.000 33.300 4.300 ;
        RECT 34.460 4.000 36.660 4.300 ;
        RECT 37.820 4.000 40.020 4.300 ;
        RECT 41.180 4.000 43.380 4.300 ;
        RECT 44.540 4.000 46.740 4.300 ;
        RECT 47.900 4.000 50.100 4.300 ;
        RECT 51.260 4.000 53.460 4.300 ;
        RECT 54.620 4.000 56.820 4.300 ;
        RECT 57.980 4.000 60.180 4.300 ;
        RECT 61.340 4.000 63.540 4.300 ;
        RECT 64.700 4.000 66.900 4.300 ;
        RECT 68.060 4.000 70.260 4.300 ;
        RECT 71.420 4.000 73.620 4.300 ;
        RECT 74.780 4.000 76.980 4.300 ;
        RECT 78.140 4.000 80.340 4.300 ;
        RECT 81.500 4.000 83.700 4.300 ;
        RECT 84.860 4.000 87.060 4.300 ;
        RECT 88.220 4.000 90.420 4.300 ;
        RECT 91.580 4.000 93.780 4.300 ;
        RECT 94.940 4.000 97.140 4.300 ;
        RECT 98.300 4.000 100.500 4.300 ;
        RECT 101.660 4.000 103.860 4.300 ;
        RECT 105.020 4.000 107.220 4.300 ;
        RECT 108.380 4.000 110.580 4.300 ;
        RECT 111.740 4.000 113.940 4.300 ;
        RECT 115.100 4.000 117.300 4.300 ;
        RECT 118.460 4.000 120.660 4.300 ;
        RECT 121.820 4.000 124.020 4.300 ;
        RECT 125.180 4.000 127.380 4.300 ;
        RECT 128.540 4.000 130.740 4.300 ;
        RECT 131.900 4.000 134.100 4.300 ;
        RECT 135.260 4.000 137.460 4.300 ;
        RECT 138.620 4.000 140.820 4.300 ;
        RECT 141.980 4.000 144.180 4.300 ;
        RECT 145.340 4.000 147.540 4.300 ;
        RECT 148.700 4.000 150.900 4.300 ;
        RECT 152.060 4.000 154.260 4.300 ;
        RECT 155.420 4.000 157.620 4.300 ;
        RECT 158.780 4.000 160.980 4.300 ;
        RECT 162.140 4.000 164.340 4.300 ;
        RECT 165.500 4.000 167.700 4.300 ;
        RECT 168.860 4.000 171.060 4.300 ;
        RECT 172.220 4.000 193.860 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 178.940 196.000 184.660 ;
        RECT 4.000 177.780 195.700 178.940 ;
        RECT 4.000 175.580 196.000 177.780 ;
        RECT 4.000 174.420 195.700 175.580 ;
        RECT 4.000 172.220 196.000 174.420 ;
        RECT 4.000 171.060 195.700 172.220 ;
        RECT 4.000 168.860 196.000 171.060 ;
        RECT 4.000 167.700 195.700 168.860 ;
        RECT 4.000 165.500 196.000 167.700 ;
        RECT 4.300 164.340 195.700 165.500 ;
        RECT 4.000 162.140 196.000 164.340 ;
        RECT 4.300 160.980 195.700 162.140 ;
        RECT 4.000 158.780 196.000 160.980 ;
        RECT 4.300 157.620 195.700 158.780 ;
        RECT 4.000 155.420 196.000 157.620 ;
        RECT 4.300 154.260 195.700 155.420 ;
        RECT 4.000 152.060 196.000 154.260 ;
        RECT 4.300 150.900 195.700 152.060 ;
        RECT 4.000 148.700 196.000 150.900 ;
        RECT 4.300 147.540 195.700 148.700 ;
        RECT 4.000 145.340 196.000 147.540 ;
        RECT 4.300 144.180 195.700 145.340 ;
        RECT 4.000 141.980 196.000 144.180 ;
        RECT 4.300 140.820 195.700 141.980 ;
        RECT 4.000 138.620 196.000 140.820 ;
        RECT 4.300 137.460 195.700 138.620 ;
        RECT 4.000 135.260 196.000 137.460 ;
        RECT 4.300 134.100 195.700 135.260 ;
        RECT 4.000 131.900 196.000 134.100 ;
        RECT 4.300 130.740 195.700 131.900 ;
        RECT 4.000 128.540 196.000 130.740 ;
        RECT 4.300 127.380 195.700 128.540 ;
        RECT 4.000 125.180 196.000 127.380 ;
        RECT 4.300 124.020 195.700 125.180 ;
        RECT 4.000 121.820 196.000 124.020 ;
        RECT 4.300 120.660 195.700 121.820 ;
        RECT 4.000 118.460 196.000 120.660 ;
        RECT 4.300 117.300 195.700 118.460 ;
        RECT 4.000 115.100 196.000 117.300 ;
        RECT 4.300 113.940 195.700 115.100 ;
        RECT 4.000 111.740 196.000 113.940 ;
        RECT 4.300 110.580 195.700 111.740 ;
        RECT 4.000 108.380 196.000 110.580 ;
        RECT 4.300 107.220 195.700 108.380 ;
        RECT 4.000 105.020 196.000 107.220 ;
        RECT 4.300 103.860 195.700 105.020 ;
        RECT 4.000 101.660 196.000 103.860 ;
        RECT 4.300 100.500 195.700 101.660 ;
        RECT 4.000 98.300 196.000 100.500 ;
        RECT 4.300 97.140 195.700 98.300 ;
        RECT 4.000 94.940 196.000 97.140 ;
        RECT 4.300 93.780 195.700 94.940 ;
        RECT 4.000 91.580 196.000 93.780 ;
        RECT 4.300 90.420 195.700 91.580 ;
        RECT 4.000 88.220 196.000 90.420 ;
        RECT 4.300 87.060 195.700 88.220 ;
        RECT 4.000 84.860 196.000 87.060 ;
        RECT 4.300 83.700 195.700 84.860 ;
        RECT 4.000 81.500 196.000 83.700 ;
        RECT 4.300 80.340 195.700 81.500 ;
        RECT 4.000 78.140 196.000 80.340 ;
        RECT 4.300 76.980 195.700 78.140 ;
        RECT 4.000 74.780 196.000 76.980 ;
        RECT 4.300 73.620 195.700 74.780 ;
        RECT 4.000 71.420 196.000 73.620 ;
        RECT 4.300 70.260 195.700 71.420 ;
        RECT 4.000 68.060 196.000 70.260 ;
        RECT 4.300 66.900 195.700 68.060 ;
        RECT 4.000 64.700 196.000 66.900 ;
        RECT 4.300 63.540 195.700 64.700 ;
        RECT 4.000 61.340 196.000 63.540 ;
        RECT 4.300 60.180 195.700 61.340 ;
        RECT 4.000 57.980 196.000 60.180 ;
        RECT 4.300 56.820 195.700 57.980 ;
        RECT 4.000 54.620 196.000 56.820 ;
        RECT 4.300 53.460 195.700 54.620 ;
        RECT 4.000 51.260 196.000 53.460 ;
        RECT 4.300 50.100 195.700 51.260 ;
        RECT 4.000 47.900 196.000 50.100 ;
        RECT 4.300 46.740 195.700 47.900 ;
        RECT 4.000 44.540 196.000 46.740 ;
        RECT 4.300 43.380 195.700 44.540 ;
        RECT 4.000 41.180 196.000 43.380 ;
        RECT 4.300 40.020 195.700 41.180 ;
        RECT 4.000 37.820 196.000 40.020 ;
        RECT 4.300 36.660 195.700 37.820 ;
        RECT 4.000 34.460 196.000 36.660 ;
        RECT 4.000 33.300 195.700 34.460 ;
        RECT 4.000 31.100 196.000 33.300 ;
        RECT 4.000 29.940 195.700 31.100 ;
        RECT 4.000 27.740 196.000 29.940 ;
        RECT 4.000 26.580 195.700 27.740 ;
        RECT 4.000 24.380 196.000 26.580 ;
        RECT 4.000 23.220 195.700 24.380 ;
        RECT 4.000 21.020 196.000 23.220 ;
        RECT 4.000 19.860 195.700 21.020 ;
        RECT 4.000 17.660 196.000 19.860 ;
        RECT 4.000 16.500 195.700 17.660 ;
        RECT 4.000 4.620 196.000 16.500 ;
      LAYER Metal4 ;
        RECT 50.540 22.490 52.240 147.190 ;
        RECT 54.440 22.490 75.550 147.190 ;
        RECT 77.750 22.490 98.860 147.190 ;
        RECT 101.060 22.490 122.170 147.190 ;
        RECT 124.370 22.490 124.740 147.190 ;
  END
END input_mux
END LIBRARY

