* NGSPICE file created from cells9.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2 D RN SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2 D SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__mux2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__mux2_1 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlya_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlya_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_16 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_16 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 D SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffq_1 D SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2 D RN SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyc_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyc_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__mux2_4 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlya_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlya_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__addf_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__addf_2 A B CI CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffq_4 D SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__invz_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__invz_2 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1 D RN SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__icgtp_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__icgtp_1 CLK E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_1 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latq_2 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4 D RN SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__icgtp_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__icgtp_4 CLK E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latrnq_2 D E RN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_4 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latsnq_1 D E SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_16 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_16 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_20 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyd_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyd_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_12 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_12 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 D RN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyb_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyb_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__invz_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__invz_8 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1 D SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latsnq_4 D E SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai33_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai33_4 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1 D RN SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2 D RN SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1 D SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffsnq_1 D SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1 D RN SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4 D SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyc_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4 D RN SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4 D SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__addf_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__addf_1 A B CI CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_16 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 D SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4 D RN SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__invz_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__invz_1 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyc_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyc_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_12 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_12 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__addh_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__addh_2 A B CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latrsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latrsnq_2 D E RN SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__icgtn_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__icgtn_2 CLKN E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__addf_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__addf_4 A B CI CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__invz_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__invz_4 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latrnq_1 D E RN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_3 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_3 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_20 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_20 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyd_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnq_2 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latq_4 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1 D RN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latrnq_4 D E RN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1 D RN SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyd_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyd_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4 D RN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or3_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4 D RN SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__hold abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__hold Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_16 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_16 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffq_2 D SE SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__invz_12 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__invz_12 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__addh_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__addh_1 A B CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latrsnq_1 D E RN SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__icgtn_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__icgtn_1 CLKN E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__invz_3 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__invz_3 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2 D RN SE SETN SI CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__icgtp_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__icgtp_2 CLK E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_2 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__addh_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__addh_4 A B CO S VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latrsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latrsnq_4 D E RN SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__icgtn_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__icgtn_4 CLKN E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_20 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_20 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnq_1 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dlyb_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dlyb_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__latsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__latsnq_2 D E SETN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai33_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai33_2 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__xor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__xor3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnq_4 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__inv_12 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__inv_12 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2 D SETN CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__bufz_8 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_8 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu9t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu9t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

.subckt cells9 clk in[0] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[1]
+ in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] out[0] out[10] out[11] out[1] out[2]
+ out[3] out[4] out[5] out[6] out[7] out[8] out[9] rst_n vdd vss
XFILLER_0_9_444 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA__254__I _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_4_193 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_409 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_40_291 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_415 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_501_ _005_ in[0] cm_inst.page\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XANTENNA_cm_inst.cc_inst.nor3_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_432_ _107_ _197_ _034_ _198_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XTAP_TAPCELL_ROW_51_481 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_51_470 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_294_ _064_ _065_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_363_ _046_ _132_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA__329__A1 _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_2_inst_B3 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_170 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_39_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai31_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_497 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA__249__I _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_37_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.buf_3_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.dffrsnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[154\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2
XFILLER_0_20_239 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_34_28 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_5_151 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__506__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_339 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_415_ _046_ _182_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_346_ _100_ cm_inst.cc_inst.out_notouch_\[26\] _116_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
XFILLER_0_51_342 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_36_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi221_1_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_277_ cm_inst.page\[4\] _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XPHY_EDGE_ROW_20_Left_72 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.xor3_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_42_342 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_299 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA__492__A3 in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_10_294 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_25_289 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_309 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_16_223 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[20\].div_flop ro_inst.counter_n\[20\] in[0] ro_inst.counter_n\[19\]
+ ro_inst.counter\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_28_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_329_ _098_ _048_ _099_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
XFILLER_0_51_172 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.dlyd_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffq_4_inst_SE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_51_70 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_30_312 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__262__I _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_397 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_183 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_356 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_38_381 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_128 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_204 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_150 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_217 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_18_191 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.and3_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and3_2
XFILLER_0_8_306 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.nand2_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_12_323 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.icgtp_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.nor4_4_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_35_362 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_35_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.sdffsnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[169\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_30_120 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.mux2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[117\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_7_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.clkbuf_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[191\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_4
XANTENNA_cm_inst.cc_inst.nand4_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_51_Left_103 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_ro_inst.gcount\[30\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_231 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.latq_4_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_41_398 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_38_253 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_38_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai222_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_49_454 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_17_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_32_429 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_17_459 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_201 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_180 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.aoi222_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_4_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.latrnq_1_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_46_435 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_41_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_418 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.invz_1_inst_EN cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_17_234 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_278 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dlya_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[176\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlya_1
X_500_ _004_ in[0] cm_inst.page\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
Xcm_inst.cc_inst.xnor3_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor3_2
XFILLER_0_48_381 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_416 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_362_ cm_inst.cc_inst.out_notouch_\[131\] cm_inst.cc_inst.out_notouch_\[139\] cm_inst.cc_inst.out_notouch_\[147\]
+ cm_inst.cc_inst.out_notouch_\[155\] _130_ _095_ _131_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_431_ cm_inst.cc_inst.out_notouch_\[70\] cm_inst.cc_inst.out_notouch_\[78\] _041_
+ _197_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_51_502 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_471 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_293_ cm_inst.page\[1\] _064_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA_cm_inst.cc_inst.oai33_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_8_171 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nand3_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_ro_inst.gcount\[9\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_14_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_465 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_37_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA__265__I _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_9_286 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_18 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_152 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[10\].div_flop ro_inst.counter_n\[10\] in[0] ro_inst.counter_n\[9\]
+ ro_inst.counter\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
X_276_ _046_ _047_ _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
X_414_ cm_inst.cc_inst.out_notouch_\[69\] cm_inst.cc_inst.out_notouch_\[77\] cm_inst.cc_inst.out_notouch_\[85\]
+ cm_inst.cc_inst.out_notouch_\[93\] _179_ _180_ _181_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.clkinv_12_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_345_ _106_ _109_ _047_ _114_ _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
XFILLER_0_51_376 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_36_373 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi221_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi221_1_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_307 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_27_362 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_223 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.xor3_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.mux4_2_inst_S0 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_2_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_251 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_273 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA__492__A4 in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.addf_1_inst_CI cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_33_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_33_310 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_28_104 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.oai21_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_16_224 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_36_181 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_328_ _022_ _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_24_343 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_24_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_3_204 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_259_ cm_inst.cc_inst.out_notouch_\[0\] cm_inst.cc_inst.out_notouch_\[8\] cm_inst.cc_inst.out_notouch_\[16\]
+ cm_inst.cc_inst.out_notouch_\[24\] _028_ _024_ _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_29_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.clkinv_16_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[202\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_16
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xcm_inst.cc_inst.dffsnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[157\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffsnq_2
XFILLER_0_15_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_382 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SE cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_424 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_13_205 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_21_260 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_12_302 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_12_335 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.nand2_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_96 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.sdffq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[159\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffq_1
XANTENNA_cm_inst.cc_inst.dffnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_47_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_7_340 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.nand4_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dffnrsnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[142\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2
XANTENNA_cm_inst.cc_inst.latq_4_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__384__S _132_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_41_399 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_21_187 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_49_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_49_455 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_232 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.oai32_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[90\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai32_1
XFILLER_0_40_452 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_31_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.latrsnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_46_436 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.latrnq_1_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.inv_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_2
XFILLER_0_22_430 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.mux2_1_inst_I0 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_479 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA__418__S0 _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_4_195 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_51_472 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_43_417 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_361_ _060_ _130_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_292_ _019_ _063_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_430_ _085_ cm_inst.cc_inst.out_notouch_\[86\] _195_ _040_ _196_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi211_1
Xro_inst.gcount\[7\].div_flop ro_inst.counter_n\[7\] in[0] ro_inst.counter_n\[6\]
+ ro_inst.counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_172 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nand3_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_500 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_10_411 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_433 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_221 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_45_363 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_413_ _064_ _180_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA_cm_inst.cc_inst.aoi21_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_344_ _111_ _113_ _114_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XANTENNA_cm_inst.cc_inst.aoi221_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_275_ cm_inst.page\[3\] _047_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XTAP_TAPCELL_ROW_11_188 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_19_244 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_42_333 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.mux4_2_inst_S1 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_SE cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_10_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_363 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_344 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_33_333 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.oai21_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[8\].div_flop_inv ro_inst.counter\[8\] ro_inst.counter_n\[8\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XTAP_TAPCELL_ROW_16_225 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_36_193 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.mux4_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[121\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_2
XFILLER_0_24_377 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_300 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_24_280 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_327_ _094_ _096_ _033_ _097_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_12_506 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_258_ cm_inst.cc_inst.out_notouch_\[32\] cm_inst.cc_inst.out_notouch_\[40\] cm_inst.cc_inst.out_notouch_\[48\]
+ cm_inst.cc_inst.out_notouch_\[56\] _028_ _024_ _030_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_ro_inst.gcount\[26\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.inv_16_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_300 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_38_383 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_447 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_403 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_13_206 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_21_261 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[33\].div_flop_inv ro_inst.counter\[33\] ro_inst.counter_n\[33\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_33_196 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.and2_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_414 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_ro_inst.gcount\[14\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.aoi21_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[68\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_4
XFILLER_0_41_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.nand4_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.dffrnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dlyb_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_26_406 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dlyc_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[183\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyc_2
XFILLER_0_34_461 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_155 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_49_456 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_222 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_44_269 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_32_85 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_17_417 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.oai211_2_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_203 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_31_453 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_23_409 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_46_437 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.oai222_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[103\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai222_2
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__509__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_447 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_17_203 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__418__S1 _122_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.mux2_1_inst_I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_4_163 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_37_Left_89 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_51_473 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_43_418 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_291_ cm_inst.cc_inst.out_notouch_\[97\] cm_inst.cc_inst.out_notouch_\[105\] cm_inst.cc_inst.out_notouch_\[113\]
+ cm_inst.cc_inst.out_notouch_\[121\] _060_ _061_ _062_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_360_ cm_inst.cc_inst.out_notouch_\[163\] cm_inst.cc_inst.out_notouch_\[171\] cm_inst.cc_inst.out_notouch_\[179\]
+ cm_inst.cc_inst.out_notouch_\[187\] _077_ _078_ _129_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
Xro_inst.gcount\[26\].div_flop_inv ro_inst.counter\[26\] ro_inst.counter_n\[26\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_31_294 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_48_Left_100 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_8_173 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nand3_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
X_489_ in[7] cm_inst.cc_inst.in\[5\] _238_ _011_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_14_228 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_1_166 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_1_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_423 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_445 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_49_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_45_320 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_33_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_9_233 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_255 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_412_ _082_ _179_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA_cm_inst.cc_inst.aoi21_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_343_ cm_inst.cc_inst.out_notouch_\[98\] cm_inst.cc_inst.out_notouch_\[106\] cm_inst.cc_inst.out_notouch_\[114\]
+ cm_inst.cc_inst.out_notouch_\[122\] _087_ _112_ _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA__472__I in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_274_ _032_ _046_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XANTENNA_cm_inst.cc_inst.addf_4_inst_A cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_11_189 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__494__I0 in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_19_245 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_342 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__382__I _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_364 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__485__I0 in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_10_275 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_37_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__292__I _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.mux2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[119\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_4
XANTENNA__476__I0 in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_3_inst_I cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_326_ cm_inst.cc_inst.out_notouch_\[130\] cm_inst.cc_inst.out_notouch_\[138\] cm_inst.cc_inst.out_notouch_\[146\]
+ cm_inst.cc_inst.out_notouch_\[154\] _077_ _095_ _096_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XTAP_TAPCELL_ROW_16_226 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_24_312 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_24_281 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_24_Left_76 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
X_257_ cm_inst.cc_inst.out_notouch_\[64\] cm_inst.cc_inst.out_notouch_\[72\] cm_inst.cc_inst.out_notouch_\[80\]
+ cm_inst.cc_inst.out_notouch_\[88\] _028_ _024_ _029_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_29_8 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.and4_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_304 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[19\].div_flop_inv ro_inst.counter\[19\] ro_inst.counter_n\[19\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XTAP_TAPCELL_ROW_13_207 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_131 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_183 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_21_262 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.and2_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_348 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_309_ _076_ _079_ _033_ _080_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA_cm_inst.cc_inst.aoi211_2_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_30_112 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xcm_inst.cc_inst.dlya_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[178\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlya_4
XANTENNA_cm_inst.cc_inst.nand4_4_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_156 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_256 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_38_234 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.inv_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_418 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_440 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.or2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[46\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or2_2
XFILLER_0_21_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_457 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_234 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_32_335 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_484 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_12_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.oai211_2_inst_C cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_11_Left_63 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.nor2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[36\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
Xcm_inst.cc_inst.addf_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[107\] cm_inst.cc_inst.out_notouch_\[108\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu9t5v0__addf_2
XFILLER_0_16_484 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.nand2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XTAP_TAPCELL_ROW_46_438 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_26_259 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_454 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_8_inst_EN cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_40_240 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_32_207 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_51_474 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.latsnq_2_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_290_ cm_inst.page\[1\] _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_23_218 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_39_395 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_488_ in[6] cm_inst.cc_inst.in\[4\] _240_ _010_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_42_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_22_251 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.mux2_2_inst_S cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_201 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_267 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_273 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_342_ _022_ _112_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_411_ cm_inst.cc_inst.out_notouch_\[101\] cm_inst.cc_inst.out_notouch_\[109\] cm_inst.cc_inst.out_notouch_\[117\]
+ cm_inst.cc_inst.out_notouch_\[125\] _137_ _138_ _178_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.addf_4_inst_B cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_273_ cm_inst.cc_inst.out_notouch_\[208\] _043_ _044_ _040_ _045_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XTAP_TAPCELL_ROW_19_246 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_39_170 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_6_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_335 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_30_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.sdffq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[161\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffq_4
XANTENNA__485__I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_2_125 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_10_265 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_21_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.aoi222_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[79\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi222_2
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_282 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_16_227 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_325_ _061_ _095_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_256_ _027_ _028_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_12_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_19_76 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_47_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_35_64 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffq_4_inst_SI cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.oai32_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[92\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai32_4
XANTENNA_cm_inst.cc_inst.and4_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi211_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_41_Left_93 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_13_208 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_154 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_316 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_21_263 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.oai21_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[81\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XANTENNA__478__I in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_4_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_308_ cm_inst.cc_inst.out_notouch_\[129\] cm_inst.cc_inst.out_notouch_\[137\] cm_inst.cc_inst.out_notouch_\[145\]
+ cm_inst.cc_inst.out_notouch_\[153\] _077_ _078_ _079_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_21_88 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xro_inst.gcount\[4\].div_flop_inv ro_inst.counter\[4\] ro_inst.counter_n\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_12_327 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi211_2_inst_C cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_124 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_376 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.icgtn_1_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_268 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_452 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_430 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_19_471 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_1_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_49_458 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_32_336 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_40_444 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_391 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_441 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.invz_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[174\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__invz_2
XANTENNA_cm_inst.cc_inst.bufz_4_inst_EN cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.sdffrsnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[165\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1
XANTENNA_cm_inst.cc_inst.addh_2_inst_A cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_439 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_34_293 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_27_43 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_9_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.icgtp_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[207\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__icgtp_1
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[6\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_51_506 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_51_475 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.latsnq_2_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_293 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.or2_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_487_ in[5] cm_inst.cc_inst.in\[3\] _240_ _009_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_22_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.bufz_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[171\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_1
XFILLER_0_10_403 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_45_399 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_45_344 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_410_ _172_ _175_ _176_ _154_ _177_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
X_341_ _110_ _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
X_272_ cm_inst.cc_inst.out_notouch_\[192\] cm_inst.cc_inst.out_notouch_\[200\] _028_
+ _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_36_377 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_8_290 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[22\].div_flop_inv ro_inst.counter\[22\] ro_inst.counter_n\[22\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
Xcm_inst.cc_inst.and2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
XTAP_TAPCELL_ROW_19_247 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_6_249 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xro_inst.gcount\[6\].div_flop ro_inst.counter_n\[6\] in[0] ro_inst.counter_n\[5\]
+ ro_inst.counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XTAP_TAPCELL_ROW_2_126 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_37_119 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_33_336 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_18_355 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_16_228 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_36_196 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_36_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_24_283 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_324_ cm_inst.cc_inst.out_notouch_\[162\] cm_inst.cc_inst.out_notouch_\[170\] cm_inst.cc_inst.out_notouch_\[178\]
+ cm_inst.cc_inst.out_notouch_\[186\] _077_ _078_ _094_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_255_ _026_ _027_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA_cm_inst.cc_inst.buf_20_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.and4_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_27_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai21_4_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SI cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi211_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_428 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.clkbuf_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_163 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_21_264 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_380 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.nor4_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor4_2
XTAP_TAPCELL_ROW_29_320 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_406 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_450 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_166 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_307_ _022_ _078_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XANTENNA_cm_inst.cc_inst.clkbuf_16_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.nand4_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand4_2
XFILLER_0_20_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_35_356 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_28_450 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_7_333 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_43_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_30_158 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_15_199 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.oai211_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[97\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_2
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.xnor2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[54\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor2_1
Xro_inst.gcount\[15\].div_flop_inv ro_inst.counter\[15\] ro_inst.counter_n\[15\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.xnor2_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_49_459 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.latrnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_32_337 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_32_88 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_32_22 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_40_412 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_40_392 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_40_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.addh_2_inst_B cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_22_412 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_1_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_19_291 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_65 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_43_10 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_40_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.or4_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_4_188 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_155 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_51_476 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.or2_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_42_410 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_342 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
X_486_ in[4] cm_inst.cc_inst.in\[2\] _240_ _008_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_22_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_1_158 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_1_169 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_415 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_10_437 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_65 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_9_203 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_9_214 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_9_225 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_45_367 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_45_356 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_5_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_13_220 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__488__I0 in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_5_146 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_36_312 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_340_ cm_inst.page\[2\] _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
X_271_ _040_ _042_ _043_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
XANTENNA_cm_inst.cc_inst.inv_8_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_19_248 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_469_ _232_ ro_inst.signal vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_50_381 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_2_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_181 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_10_234 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_10_278 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_289 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_2_127 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_SI cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_18_301 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_367 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[23\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.aoi22_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[69\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XFILLER_0_49_470 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.nor3_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_16_229 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_323_ _093_ ro_inst.counter\[1\] _016_ out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XTAP_TAPCELL_ROW_24_284 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_24_359 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_24_304 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_254_ _019_ _026_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.and4_2_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_304 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.nor2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[38\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_4
XFILLER_0_38_407 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[11\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_46_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_33_123 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xcm_inst.cc_inst.nand2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_4
XFILLER_0_37_440 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_306_ _026_ _077_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_24_189 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.buf_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_8 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_35_357 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_440 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_465 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_454 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.clkinv_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[197\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_2
XANTENNA_cm_inst.cc_inst.xnor2_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_159 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_338 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nor2_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_40_393 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai32_2_inst_B1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_476 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_186 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_476 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.latsnq_1_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.icgtp_1_inst_TE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[29\].div_flop ro_inst.counter_n\[29\] in[0] ro_inst.counter_n\[28\]
+ ro_inst.counter\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_27_67 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_45_430 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_273 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_25_262 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai222_1_inst_C1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_4_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_17_207 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.buf_3_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_3
XANTENNA_cm_inst.cc_inst.or4_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_15_Left_67 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.and4_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and4_2
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_51_477 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_51_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_42_411 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_485_ in[3] cm_inst.cc_inst.in\[1\] _240_ _007_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA_cm_inst.cc_inst.bufz_16_inst_EN cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.aoi211_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[73\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_2
XFILLER_0_9_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_259 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_18_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__497__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_265 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA__488__I1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_5_147 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_13_298 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.latq_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[124\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latq_2
XANTENNA__309__S _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_270_ _041_ _042_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
Xcm_inst.cc_inst.oai21_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[83\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_4
XANTENNA_cm_inst.cc_inst.dffsnq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_468_ _228_ _229_ _230_ _231_ ro_sel\[2\] ro_sel\[1\] _232_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.oai33_1_inst_B1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_19_249 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_42_338 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.inv_8_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_8
XFILLER_0_27_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_399_ cm_inst.cc_inst.out_notouch_\[36\] cm_inst.cc_inst.out_notouch_\[44\] cm_inst.cc_inst.out_notouch_\[52\]
+ cm_inst.cc_inst.out_notouch_\[60\] _083_ _122_ _167_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_10_182 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_15_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.latrnq_2_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_2_128 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_18_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_379 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_18_Left_70 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SETN cm_inst.cc_inst.in\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nor3_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_322_ _058_ _073_ _092_ _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor3_1
XFILLER_0_36_143 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_32_360 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_24_285 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.dlyb_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[179\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyb_1
X_253_ cm_inst.cc_inst.out_notouch_\[96\] cm_inst.cc_inst.out_notouch_\[104\] cm_inst.cc_inst.out_notouch_\[112\]
+ cm_inst.cc_inst.out_notouch_\[120\] _021_ _024_ _025_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_35_56 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_27_187 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_30_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_23_393 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_23_360 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.sdffrsnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[167\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4
XANTENNA_cm_inst.cc_inst.oai221_2_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_38_377 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_146 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_135 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_143 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_187 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_3_Left_55 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.oai221_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[99\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai221_1
X_305_ cm_inst.cc_inst.out_notouch_\[161\] cm_inst.cc_inst.out_notouch_\[169\] cm_inst.cc_inst.out_notouch_\[177\]
+ cm_inst.cc_inst.out_notouch_\[185\] _027_ _023_ _076_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XTAP_TAPCELL_ROW_12_200 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_24_168 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_35_358 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.xor3_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_452 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_7_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_7_368 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_7_379 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_168 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.icgtp_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[209\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__icgtp_4
XPHY_EDGE_ROW_45_Left_97 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_238 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_38_227 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.latrnq_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[127\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latrnq_2
XFILLER_0_34_444 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[19\].div_flop ro_inst.counter_n\[19\] in[0] ro_inst.counter_n\[18\]
+ ro_inst.counter\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XTAP_TAPCELL_ROW_40_394 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_32_339 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_400 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nor2_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.bufz_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[172\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_4
XANTENNA_cm_inst.cc_inst.oai32_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai32_2_inst_B2 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_48_450 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_16_400 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_271 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_3_360 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_252 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_34_274 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai221_4_inst_C cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.and2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_4
XTAP_TAPCELL_ROW_45_431 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai222_1_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai222_1_inst_C2 cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnq_2_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffsnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[11\].div_flop_inv ro_inst.counter\[11\] ro_inst.counter_n\[11\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.or4_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_12_inst_EN cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_40_299 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__420__S _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_48_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_51_478 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.latsnq_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[132\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latsnq_1
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_31_277 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.xor2_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_285 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_8_167 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.clkbuf_8_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
X_484_ _238_ _240_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XPHY_EDGE_ROW_32_Left_84 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA__266__S1 _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_ro_inst.gcount\[19\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_45 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__304__I _074_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_45_336 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_45_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.bufz_16_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[173\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_16
XANTENNA_cm_inst.cc_inst.latrsnq_1_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_277 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_5_148 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.oai33_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[93\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai33_1
XFILLER_0_36_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_8_271 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_1_inst_B2 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dffq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[148\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_2
X_467_ _210_ _224_ _225_ _231_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_27_358 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_398_ _081_ _165_ _120_ _166_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XFILLER_0_24_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_208 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_183 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_49_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.latrnq_2_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_2_129 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_33_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_41_361 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.xnor2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[56\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor2_4
XFILLER_0_49_483 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.nor3_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_321_ _075_ _080_ _090_ _091_ _092_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
X_252_ _023_ _024_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_339 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_68 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.buf_20_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_20
XANTENNA__473__B in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_144 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_15_306 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_15_220 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_2_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.invz_8_inst_EN cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai221_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai221_2_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_38_378 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_158 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_155 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_394 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_304_ _074_ _075_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
Xro_inst.gcount\[5\].div_flop ro_inst.counter_n\[5\] in[0] ro_inst.counter_n\[4\]
+ ro_inst.counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XTAP_TAPCELL_ROW_12_201 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__312__I _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_158 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.aoi221_4_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_20_397 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_47_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_359 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_28_431 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_28_442 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__502__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.xor3_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_7_336 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_19_442 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.aoi221_4_inst_C cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_380 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_40_395 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_32_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_25_412 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__307__I _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai32_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_161 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_20_183 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_48_451 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_31_415 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_22_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_297 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_27_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_ro_inst.gcount\[3\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_45_432 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai222_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai222_1_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_13_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or4_2_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_51_479 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_51_468 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.aoi221_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[75\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi221_1
XANTENNA_cm_inst.cc_inst.xor2_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_453 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_253 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_8_168 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.aoi22_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[71\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_4
XFILLER_0_16_297 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.clkinv_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_483_ in[2] cm_inst.cc_inst.in\[0\] _239_ _006_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_22_234 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_10_407 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_429 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dlyb_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SE cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_45_359 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_45_348 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dlyd_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[186\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyd_2
XFILLER_0_9_217 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_5_149 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__405__I _074_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_294 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai33_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_1_inst_B3 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_120 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_397_ cm_inst.cc_inst.out_notouch_\[4\] cm_inst.cc_inst.out_notouch_\[12\] _118_
+ _165_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_466_ _128_ _146_ ro_sel\[0\] _230_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_10_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_10_184 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__426__S _132_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_18_240 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.invz_4_inst_EN cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_359 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_51_104 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_320_ cm_inst.page\[4\] _091_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
X_251_ _022_ _023_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_36_189 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_32_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_24_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_20_502 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nand3_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_15_221 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_449_ cm_inst.cc_inst.out_notouch_\[199\] cm_inst.cc_inst.out_notouch_\[207\] _042_
+ _214_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_27_134 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_379 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai221_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_137 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_14_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.icgtp_4_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_303_ _035_ _074_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_24_126 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.aoi221_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.aoi221_4_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_7_348 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.xor3_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.addf_4_inst_CI cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_432 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_181 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_218 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_396 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_37_262 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_25_435 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_0_502 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai32_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_48_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_452 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nand2_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_4_inst_I cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_31_330 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_298 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.clkinv_12_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[201\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_12
XFILLER_0_34_243 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_295 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_471 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_14 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_27_59 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xcm_inst.cc_inst.dffnrnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[139\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2
XFILLER_0_45_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_43_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.oai222_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_4_159 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_36_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_51_469 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_210 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_16_221 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_8_169 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_12_482 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_482_ _235_ _239_ _055_ _237_ _005_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XFILLER_0_27_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.oai22_2_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_ro_inst.gcount\[32\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dlyb_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[181\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyb_4
XFILLER_0_38_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_229 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.invz_8_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[175\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__invz_8
XANTENNA_cm_inst.cc_inst.inv_3_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_202 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_224 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.or3_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or3_2
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_28_91 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xro_inst.gcount\[28\].div_flop ro_inst.counter_n\[28\] in[0] ro_inst.counter_n\[27\]
+ ro_inst.counter\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_51_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_465_ _171_ _189_ _225_ _229_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
Xcm_inst.cc_inst.oai221_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[101\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai221_4
XANTENNA_cm_inst.cc_inst.oai33_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.nor3_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor3_1
XANTENNA_ro_inst.gcount\[20\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_396_ _084_ cm_inst.cc_inst.out_notouch_\[20\] _163_ _105_ _164_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi211_1
Xcm_inst.cc_inst.dffnsnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[144\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1
XTAP_TAPCELL_ROW_10_185 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.nand3_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand3_1
XFILLER_0_18_305 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_18_241 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.mux2_4_inst_I0 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[29\].div_flop_inv ro_inst.counter\[29\] ro_inst.counter_n\[29\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XTAP_TAPCELL_ROW_1_120 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_51_138 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_36_135 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_250_ cm_inst.page\[1\] _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_24_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_360 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nand3_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_51_36 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_448_ _211_ _212_ _120_ _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_7_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_15_222 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_379_ _146_ ro_inst.counter\[3\] _147_ out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_23_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_50_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_50_Left_102 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.mux4_1_inst_S0 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_21_258 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_341 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_29_314 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_302_ _059_ _072_ _073_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
XFILLER_0_37_444 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_9_390 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_32_193 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.aoi221_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.dffrnq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_34_350 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_46_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.latsnq_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[134\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latsnq_4
XFILLER_0_34_436 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_414 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XPHY_EDGE_ROW_7_Left_59 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_40_397 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_48_453 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nand2_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_31_417 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_31_331 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_28_296 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_263 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_3_396 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_3_341 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_152 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.oai33_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[95\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai33_4
XANTENNA_cm_inst.cc_inst.aoi22_2_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_25_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_21_450 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_428 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_23_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xcm_inst.cc_inst.oai22_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[84\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai22_1
Xro_inst.gcount\[18\].div_flop ro_inst.counter_n\[18\] in[0] ro_inst.counter_n\[17\]
+ ro_inst.counter\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_16_233 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_299 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_481_ _234_ _239_ _091_ _237_ _004_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XANTENNA_cm_inst.cc_inst.oai22_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai22_2_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_38_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_196 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_44_350 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dlyc_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_263 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XPHY_EDGE_ROW_36_Left_88 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.dffrnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_4_140 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_464_ _225_ _056_ _227_ _228_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XFILLER_0_35_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.mux4_2_inst_I0 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_23_501 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_395_ _100_ cm_inst.cc_inst.out_notouch_\[28\] _163_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
Xcm_inst.cc_inst.dffrsnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[153\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1
XTAP_TAPCELL_ROW_10_186 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_18_242 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_45_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__505__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.mux2_4_inst_I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_1_121 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_32_364 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.sdffrnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[163\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2
XANTENNA_cm_inst.cc_inst.nand3_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_447_ cm_inst.cc_inst.out_notouch_\[135\] cm_inst.cc_inst.out_notouch_\[143\] cm_inst.cc_inst.out_notouch_\[151\]
+ cm_inst.cc_inst.out_notouch_\[159\] _118_ _098_ _212_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_378_ ro_inst.enable _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
X_516_ out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tiel
XANTENNA__342__I _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_23_397 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_23_342 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_60 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_46_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.mux4_1_inst_S1 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_147 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_259 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_29_315 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_37_370 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_301_ _068_ _071_ _036_ _072_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA_cm_inst.cc_inst.dffq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_37_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_39_Left_91 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA__337__I _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_415 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_23_Left_75 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.and3_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and3_1
XTAP_TAPCELL_ROW_34_351 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_34_448 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.aoi221_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[77\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi221_4
XFILLER_0_6_372 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_14_172 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_220 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.oai211_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_404 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_4_309 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.sdffsnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[168\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.clkbuf_3_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[190\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_3
XFILLER_0_28_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.icgtn_1_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_ro_inst.gcount\[28\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_31_407 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_332 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_16_404 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_437 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.invz_1_inst_I cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[4\].div_flop ro_inst.counter_n\[4\] in[0] ro_inst.counter_n\[3\]
+ ro_inst.counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_3_364 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.aoi22_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi22_2_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_481 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_43_49 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xro_inst.gcount\[7\].div_flop_inv ro_inst.counter\[7\] ro_inst.counter_n\[7\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.clkbuf_3_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_4_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_ro_inst.gcount\[16\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_8_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_16_289 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_10_Left_62 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_42_405 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_304 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_480_ _233_ _239_ _172_ _237_ _003_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XANTENNA_cm_inst.cc_inst.oai22_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_22_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.clkinv_8_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[200\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_8
XFILLER_0_38_49 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xcm_inst.cc_inst.xnor3_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor3_1
Xro_inst.gcount\[32\].div_flop_inv ro_inst.counter\[32\] ro_inst.counter_n\[32\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XTAP_TAPCELL_ROW_7_160 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_5_415 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_44_362 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_44_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_8_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_286 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.and3_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_4_141 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.dffrnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[151\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_2
X_463_ _127_ _226_ _073_ _092_ _227_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or4_1
X_394_ _157_ _159_ _047_ _161_ _162_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
XANTENNA_cm_inst.cc_inst.mux4_2_inst_I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_10_187 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_18_243 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__399__S1 _122_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_201 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_41_354 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_30_61 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_1_122 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_49_487 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_49_454 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_24_279 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_17_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_515_ out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tiel
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
X_446_ cm_inst.cc_inst.out_notouch_\[167\] cm_inst.cc_inst.out_notouch_\[175\] cm_inst.cc_inst.out_notouch_\[183\]
+ cm_inst.cc_inst.out_notouch_\[191\] _149_ _150_ _211_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_377_ _049_ _135_ _145_ _127_ _146_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
XANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_23_310 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_18_159 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.tiel_inst cm_inst.cc_inst.out_notouch_\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tiel
XANTENNA_cm_inst.cc_inst.dffnsnq_2_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_398 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_316 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_37_371 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_300_ _069_ _070_ _067_ _071_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
Xcm_inst.cc_inst.dffsnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[156\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffsnq_1
Xro_inst.gcount\[25\].div_flop_inv ro_inst.counter\[25\] ro_inst.counter_n\[25\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_32_162 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__299__S0 _063_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_379 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_446 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_7_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_429_ _021_ cm_inst.cc_inst.out_notouch_\[94\] _195_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
XFILLER_0_23_195 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_11_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.and4_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_34_352 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_6_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_40_Left_92 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.dffnrsnq_1_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_32_18 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_37_254 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai211_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_482 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.inv_12_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dffnrsnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[141\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1
XTAP_TAPCELL_ROW_31_333 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_3_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.latrsnq_1_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_11_187 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_39_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.aoi211_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi22_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_463 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.nor3_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor3_4
Xcm_inst.cc_inst.dffnsnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[146\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4
XFILLER_0_21_430 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_13_408 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_452 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.nand3_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand3_4
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_16_202 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.inv_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XTAP_TAPCELL_ROW_42_406 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_50_461 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_35_500 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xro_inst.gcount\[18\].div_flop_inv ro_inst.counter\[18\] ro_inst.counter_n\[18\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XTAP_TAPCELL_ROW_7_161 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SI cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_382 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_13_216 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_360 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_298 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_17_500 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.and3_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.xor2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[61\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor2_2
XTAP_TAPCELL_ROW_4_142 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_393_ _111_ _160_ _161_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
X_462_ ro_sel\[0\] _226_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
XFILLER_0_50_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.mux4_2_inst_I2 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_82 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_1_123 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_36_127 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_32_366 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_32_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_374 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_506 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_514_ out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tiel
X_445_ _210_ ro_inst.counter\[34\] _147_ out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_376_ _059_ _144_ _145_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
XANTENNA__458__A2 _222_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dlya_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[27\].div_flop ro_inst.counter_n\[27\] in[0] ro_inst.counter_n\[26\]
+ ro_inst.counter\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XANTENNA_cm_inst.cc_inst.oai31_1_inst_B cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_94 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.mux4_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[120\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_333 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_37_372 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_29_317 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_20_303 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_428_ _172_ _192_ _193_ _154_ _194_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
X_359_ _128_ ro_inst.counter\[2\] _016_ out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_51_494 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xcm_inst.cc_inst.oai22_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[86\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai22_4
XFILLER_0_36_61 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.and4_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_34_353 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_436 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_469 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_14_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_200 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_0_506 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_334 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_28_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_22_41 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.latrsnq_1_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dlyc_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[182\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyc_1
XANTENNA__380__S0 _130_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi211_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_258 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__274__I _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_299 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_426 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_21_442 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_303 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dffrsnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[155\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4
XFILLER_0_21_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__362__S0 _130_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.oai222_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[102\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai222_1
XANTENNA__508__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_3_inst_EN cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_214 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_16_225 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_12_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_407 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_50_462 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_7_162 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_372 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_13_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.bufz_16_inst_I cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[3\].div_flop_inv ro_inst.counter\[3\] ro_inst.counter_n\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_0_188 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.dffsnq_2_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.and3_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_461_ ro_sel\[0\] _225_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XTAP_TAPCELL_ROW_4_143 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.mux4_2_inst_I3 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_392_ cm_inst.cc_inst.out_notouch_\[100\] cm_inst.cc_inst.out_notouch_\[108\] cm_inst.cc_inst.out_notouch_\[116\]
+ cm_inst.cc_inst.out_notouch_\[124\] _087_ _112_ _160_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
Xro_inst.gcount\[17\].div_flop ro_inst.counter_n\[17\] in[0] ro_inst.counter_n\[16\]
+ ro_inst.counter\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XANTENNA__493__I0 in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_309 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_63 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_30_41 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_26_375 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_203 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_1_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_124 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xcm_inst.cc_inst.and3_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and3_4
XFILLER_0_49_478 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_49_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.dffsnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffrnq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_331 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_364 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_32_389 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__475__I0 in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_ro_inst.gcount\[8\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_444_ _018_ _194_ _209_ _058_ _210_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
Xcm_inst.cc_inst.sdffsnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[170\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4
X_513_ out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tiel
X_375_ _140_ _143_ _036_ _144_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA_cm_inst.cc_inst.icgtn_4_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_23_356 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_23_334 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_23_389 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_84 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_25_74 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_172 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_345 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_29_318 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_37_373 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_37_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_9_394 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_20_251 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__376__A2 _144_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_358_ _049_ _103_ _126_ _127_ _128_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
X_427_ cm_inst.cc_inst.out_notouch_\[198\] cm_inst.cc_inst.out_notouch_\[206\] _101_
+ _193_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_36_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_289_ _019_ _060_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.and4_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_34_354 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_131 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_42_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or3_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA__470__I in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.xnor3_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor3_4
XPHY_EDGE_ROW_27_Left_79 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_20_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[21\].div_flop_inv ro_inst.counter\[21\] ro_inst.counter_n\[21\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_43_248 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_ro_inst.slow_clock_inv_I in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.or2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[45\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or2_1
XFILLER_0_3_345 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_356 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_189 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__290__I cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_45_427 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.addf_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[105\] cm_inst.cc_inst.out_notouch_\[106\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu9t5v0__addf_1
XANTENNA_cm_inst.cc_inst.latrnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_410 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_8_437 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_16_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA__353__S1 _122_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_50_463 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_42_408 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_50_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_163 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.buf_16_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_16
XFILLER_0_38_340 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_38_395 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.nor2_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[3\].div_flop ro_inst.counter_n\[3\] in[0] ro_inst.counter_n\[2\]
+ ro_inst.counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XANTENNA_cm_inst.cc_inst.clkinv_20_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_240 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.icgtn_2_inst_TE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_85 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_28_96 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or4_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_340 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_234 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_14_Left_66 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_44_354 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_144 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_460_ _224_ ro_inst.saved_signal ro_inst.enable out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_391_ _107_ _158_ _034_ _159_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
Xcm_inst.cc_inst.dffsnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[158\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffsnq_4
XANTENNA_cm_inst.cc_inst.dffq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_23_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.icgtp_4_inst_TE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[14\].div_flop_inv ro_inst.counter\[14\] ro_inst.counter_n\[14\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_38_181 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_41_357 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai222_4_inst_C1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_343 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.xnor3_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_374_ _141_ _142_ _067_ _143_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_512_ _243_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tiel
X_443_ _201_ _208_ _017_ _209_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_1
XTAP_TAPCELL_ROW_15_216 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.aoi222_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[78\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi222_1
XFILLER_0_31_390 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.dffnrsnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[143\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4
XANTENNA_cm_inst.cc_inst.clkinv_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_29_319 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_49_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_374 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__293__I cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_162 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_20_252 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_43_419 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_357_ cm_inst.page\[5\] _127_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
X_426_ _190_ _191_ _132_ _192_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA_cm_inst.cc_inst.oai33_4_inst_B1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_288_ cm_inst.page\[4\] _059_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai211_4_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__447__S0 _118_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_34_355 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.and4_1_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_332 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.inv_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_4
XANTENNA_cm_inst.cc_inst.or3_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_ro_inst.gcount\[25\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_181 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_430 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_2_Left_54 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_0_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_20_157 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_48_447 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_409_ cm_inst.cc_inst.out_notouch_\[197\] cm_inst.cc_inst.out_notouch_\[205\] _042_
+ _176_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_3_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_408 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_44_Left_96 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_19_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.invz_1_inst cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[173\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__invz_1
XFILLER_0_34_249 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.clkbuf_12_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_485 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_ro_inst.gcount\[13\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_45_428 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_21_455 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_0_305 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.sdffq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai32_1_inst_B1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_271 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_42_409 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_50_464 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.nor4_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_296 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_7_164 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__421__A2 _187_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nor2_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_5_419 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.or4_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.mux4_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[122\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_4
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_4_145 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__296__I _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_390_ cm_inst.cc_inst.out_notouch_\[68\] cm_inst.cc_inst.out_notouch_\[76\] _041_
+ _158_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XPHY_EDGE_ROW_31_Left_83 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_26_300 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_216 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai222_4_inst_C2 cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai222_4_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_303 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_249 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_32_303 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_4_260 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi21_1_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.xor2_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.xnor3_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_511_ _015_ in[0] ro_sel\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
X_373_ cm_inst.cc_inst.out_notouch_\[3\] cm_inst.cc_inst.out_notouch_\[11\] cm_inst.cc_inst.out_notouch_\[19\]
+ cm_inst.cc_inst.out_notouch_\[27\] _137_ _138_ _142_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_27_119 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_442_ _203_ _205_ _037_ _207_ _208_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
XTAP_TAPCELL_ROW_23_272 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_15_217 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.aoi211_4_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_26_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_26_141 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.dlyc_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[184\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyc_4
XFILLER_0_14_303 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_22_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai31_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_37_375 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_9_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.inv_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_32_166 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_32_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_253 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_20_339 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.or4_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or4_2
Xcm_inst.cc_inst.bufz_12_inst cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[172\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_12
XANTENNA_cm_inst.cc_inst.oai33_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_4_inst_B2 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.latsnq_4_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_425_ cm_inst.cc_inst.out_notouch_\[134\] cm_inst.cc_inst.out_notouch_\[142\] cm_inst.cc_inst.out_notouch_\[150\]
+ cm_inst.cc_inst.out_notouch_\[158\] _149_ _150_ _191_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_287_ cm_inst.page\[5\] _058_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_28_439 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_356_ _115_ _125_ _017_ _126_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_1
XFILLER_0_23_199 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.addh_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[113\]
+ cm_inst.cc_inst.out_notouch_\[114\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__addh_2
XANTENNA_cm_inst.cc_inst.oai211_4_inst_C cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.oai222_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[104\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai222_4
Xcm_inst.cc_inst.nor4_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor4_1
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__447__S1 _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_417 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnq_1_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai221_1_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_450 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.nand4_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand4_1
XANTENNA_cm_inst.cc_inst.or3_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[26\].div_flop ro_inst.counter_n\[26\] in[0] ro_inst.counter_n\[25\]
+ ro_inst.counter\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_37_258 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_160 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_9_193 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_461 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_442 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_48_448 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.oai211_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[96\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
X_408_ _173_ _174_ _132_ _175_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_43_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_3_347 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_339_ _107_ _108_ _034_ _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XFILLER_0_11_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_37_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_2_32 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.latsnq_4_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_217 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_30_467 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_45_429 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_434 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.latrsnq_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[130\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latrsnq_2
XFILLER_0_33_10 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.mux2_4_inst_S cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai32_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_217 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai32_1_inst_B2 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.icgtn_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[205\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__icgtn_2
XANTENNA_cm_inst.cc_inst.nor4_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_50_465 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_7_165 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.dlyd_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.buf_16_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.or4_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_320 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_44_312 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_364 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_12_286 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__487__I0 in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_2_inst_C1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_18_237 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai222_4_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai222_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_507 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_161 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_17_301 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.xor2_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_356 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_378 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__301__S _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__321__A2 _080_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.xnor3_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_510_ _014_ in[0] ro_sel\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
X_441_ _110_ _206_ _207_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XFILLER_0_35_131 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_372_ cm_inst.cc_inst.out_notouch_\[35\] cm_inst.cc_inst.out_notouch_\[43\] cm_inst.cc_inst.out_notouch_\[51\]
+ cm_inst.cc_inst.out_notouch_\[59\] _137_ _065_ _141_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.latq_1_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_23_273 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_15_218 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_35_197 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_23_326 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.aoi211_4_inst_C cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_134 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_41_65 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_41_76 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xro_inst.gcount\[10\].div_flop_inv ro_inst.counter\[10\] ro_inst.counter_n\[10\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_14_337 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_1_231 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai31_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.or2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[47\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or2_4
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_37_376 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[16\].div_flop ro_inst.counter_n\[16\] in[0] ro_inst.counter_n\[15\]
+ ro_inst.counter\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_9_397 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_17_164 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_20_254 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_20_307 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_28_310 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.addf_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[109\] cm_inst.cc_inst.out_notouch_\[110\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu9t5v0__addf_4
XANTENNA_cm_inst.cc_inst.oai33_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_424_ cm_inst.cc_inst.out_notouch_\[166\] cm_inst.cc_inst.out_notouch_\[174\] cm_inst.cc_inst.out_notouch_\[182\]
+ cm_inst.cc_inst.out_notouch_\[190\] _130_ _095_ _190_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.oai33_4_inst_B3 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_51_410 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_286_ _016_ _056_ _057_ out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
X_355_ _117_ _121_ _074_ _124_ _125_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
XANTENNA_cm_inst.cc_inst.dffrnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.addh_4_inst_A cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai221_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai221_1_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_484 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_123 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_14_189 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_395 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_48_449 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_407_ cm_inst.cc_inst.out_notouch_\[133\] cm_inst.cc_inst.out_notouch_\[141\] cm_inst.cc_inst.out_notouch_\[149\]
+ cm_inst.cc_inst.out_notouch_\[157\] _149_ _098_ _174_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_338_ cm_inst.cc_inst.out_notouch_\[66\] cm_inst.cc_inst.out_notouch_\[74\] _041_
+ _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_51_240 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_269_ _026_ _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.clkinv_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[196\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.latsnq_4_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_2_22 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_131 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_42_251 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.latrsnq_4_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_446 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_281 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_44_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_33_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_33_88 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_16_229 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai32_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffsnq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_273 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.clkinv_8_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nor4_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_50_466 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_30_221 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_15_240 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.buf_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_2
XFILLER_0_30_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_166 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.and4_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and4_1
XTAP_TAPCELL_ROW_41_400 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_38_310 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.aoi222_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[80\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi222_4
XFILLER_0_41_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.or4_1_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nand2_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__487__I1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.aoi211_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[72\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
XANTENNA_cm_inst.cc_inst.icgtn_2_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__496__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.invz_2_inst_I cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_2_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_2_inst_C2 cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.latq_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[123\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latq_1
XTAP_TAPCELL_ROW_18_238 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_41_349 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_26_379 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_302 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_26_293 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_ro_inst.gcount\[5\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai222_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SE cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_49_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.clkbuf_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_335 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_251 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_40_393 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[2\].div_flop ro_inst.counter_n\[2\] in[0] ro_inst.counter_n\[1\]
+ ro_inst.counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
X_371_ _136_ _139_ _067_ _140_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_440_ cm_inst.cc_inst.out_notouch_\[38\] cm_inst.cc_inst.out_notouch_\[46\] cm_inst.cc_inst.out_notouch_\[54\]
+ cm_inst.cc_inst.out_notouch_\[62\] _083_ _112_ _206_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XTAP_TAPCELL_ROW_15_219 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.latq_1_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_23_338 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_23_274 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_31_382 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__511__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_22 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_41_88 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_1_221 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_393 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_22_382 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai31_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.invz_3_inst_EN cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.invz_4_inst cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[174\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__invz_4
XTAP_TAPCELL_ROW_20_255 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_13_382 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_28_311 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_423_ _189_ ro_inst.counter\[5\] _147_ out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_354_ _110_ _123_ _124_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XANTENNA_cm_inst.cc_inst.oai33_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_51_444 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_285_ ro_inst.counter\[0\] ro_inst.enable _057_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XFILLER_0_3_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.addh_4_inst_B cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai221_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_419 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_22_190 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_135 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_14_168 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_173 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_406_ cm_inst.cc_inst.out_notouch_\[165\] cm_inst.cc_inst.out_notouch_\[173\] cm_inst.cc_inst.out_notouch_\[181\]
+ cm_inst.cc_inst.out_notouch_\[189\] _130_ _150_ _173_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XTAP_TAPCELL_ROW_31_328 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_337_ _098_ _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_28_238 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.latrnq_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[126\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latrnq_1
XFILLER_0_51_274 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
X_268_ _039_ _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_47_43 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.mux4_4_inst_S0 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffq_2_inst_SE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.bufz_3_inst cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[171\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_3
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_425 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_6_Left_58 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_18_271 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_18_293 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_420 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai32_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_50_467 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nor4_2_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_15_274 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nand4_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_41_401 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_399 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_506 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_21_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_89 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_344 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_29_333 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_322 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_8_238 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.nand2_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_44_358 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_7_260 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.inv_20_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_20
XANTENNA_cm_inst.cc_inst.latrsnq_2_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_2_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai22_1_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_26_294 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_9_Left_61 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_18_239 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_30_57 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.nor4_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor4_4
XTAP_TAPCELL_ROW_1_118 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.dffq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[147\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XFILLER_0_17_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_17_347 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.nand4_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand4_4
X_370_ cm_inst.cc_inst.out_notouch_\[67\] cm_inst.cc_inst.out_notouch_\[75\] cm_inst.cc_inst.out_notouch_\[83\]
+ cm_inst.cc_inst.out_notouch_\[91\] _137_ _138_ _139_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_35_133 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_35_Left_87 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_23_275 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_16_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_394 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.oai211_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[98\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_4
XANTENNA_ro_inst.gcount\[34\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_499_ _003_ in[0] cm_inst.page\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_22_361 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_45_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_256 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.sig_cmp ro_inst.signal ro_inst.saved_signal ro_inst.running vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__xnor2_1
XTAP_TAPCELL_ROW_28_312 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_36_453 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_422_ _018_ _177_ _188_ _058_ _189_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
X_284_ _018_ _038_ _054_ _055_ _056_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
X_353_ cm_inst.cc_inst.out_notouch_\[34\] cm_inst.cc_inst.out_notouch_\[42\] cm_inst.cc_inst.out_notouch_\[50\]
+ cm_inst.cc_inst.out_notouch_\[58\] _083_ _122_ _123_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_51_478 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_ro_inst.gcount\[22\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_45 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xcm_inst.cc_inst.xor3_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[64\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor3_2
XFILLER_0_27_442 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_6_336 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_10_364 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_163 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_33_434 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__501__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_31_329 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_405_ _074_ _172_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA_ro_inst.gcount\[10\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_267_ cm_inst.page\[1\] _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
XFILLER_0_3_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai21_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_336_ _085_ cm_inst.cc_inst.out_notouch_\[82\] _104_ _105_ _106_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi211_1
XPHY_EDGE_ROW_38_Left_90 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_47_440 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_22_Left_74 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA__408__S _132_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_228 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.mux4_4_inst_S1 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dlya_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_401 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_10_161 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xro_inst.gcount\[28\].div_flop_inv ro_inst.counter\[28\] ro_inst.counter_n\[28\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
Xro_inst.slow_clock_inv in[0] ro_inst.slow_clk_n vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SE cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai31_2_inst_B cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.addf_1_inst_A cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_459 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_44_421 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_3_158 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.clkbuf_20_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[195\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_20
X_319_ _086_ _089_ _048_ _090_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_1
Xro_inst.gcount\[25\].div_flop ro_inst.counter_n\[25\] in[0] ro_inst.counter_n\[24\]
+ ro_inst.counter\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_35_6 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.aoi22_1_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_7_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.nand4_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_41_402 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_301 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.latrnq_4_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_234 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_356 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__333__A2 _097_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_4_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_12_278 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.oai31_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[88\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai31_2
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_35_348 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_315 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_250 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xcm_inst.cc_inst.dlyd_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[185\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyd_1
XANTENNA_cm_inst.cc_inst.latrsnq_2_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai22_1_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai22_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.latrsnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_26_295 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_26_348 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_1_119 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_32_307 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_4_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_253 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_48_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_276 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.dffnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[136\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnq_2
XANTENNA_cm_inst.cc_inst.mux4_1_inst_I0 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_24 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_39_484 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_498_ _002_ in[0] cm_inst.page\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XFILLER_0_26_189 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_14_210 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_14_307 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_41_126 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xcm_inst.cc_inst.clkinv_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[199\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_4
XFILLER_0_22_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_334 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_20_257 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_40_192 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_373 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_28_313 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_421_ _059_ _187_ _188_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
XFILLER_0_36_410 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.aoi21_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_283_ cm_inst.page\[5\] _055_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
X_352_ _064_ _122_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_23_137 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_34_349 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_27_454 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_376 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_SE cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_9_197 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_18_465 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_33_446 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.and4_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and4_4
XANTENNA_cm_inst.cc_inst.invz_8_inst_I cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__295__S0 _063_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.ring_osc_0 ro_inst.ring\[0\] ro_inst.enable ro_inst.ring\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
X_404_ _171_ ro_inst.counter\[4\] _147_ out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_335_ _039_ _105_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_266_ _025_ _029_ _030_ _031_ _034_ _037_ _038_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.oai21_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_47_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xro_inst.gcount\[15\].div_flop ro_inst.counter_n\[15\] in[0] ro_inst.counter_n\[14\]
+ ro_inst.counter\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XTAP_TAPCELL_ROW_47_441 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_47_67 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_6_123 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_42_221 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.aoi211_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[74\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_4
XANTENNA__499__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.addf_1_inst_B cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.and2_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.latq_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[125\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latq_4
XANTENNA_cm_inst.cc_inst.oai211_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.tieh_inst cm_inst.cc_inst.out_notouch_\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__tieh
XTAP_TAPCELL_ROW_44_422 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_58 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_33_14 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_232 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_249_ _020_ _021_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
X_318_ _040_ _088_ _089_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XANTENNA_cm_inst.cc_inst.dffnrnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dffnrnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[138\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1
XFILLER_0_47_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_35_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.and4_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi22_1_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi22_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nand4_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_41_403 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_26_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_28_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.latrnq_4_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_368 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_17_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_139 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_31_500 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.or3_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or3_1
XANTENNA_cm_inst.cc_inst.oai22_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_26_296 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_390 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_382 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_1_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_17_230 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_4_243 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_349 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_ro_inst.gcount\[18\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_23_277 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.and3_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_393 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xcm_inst.cc_inst.latrnq_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[128\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latrnq_4
XANTENNA_cm_inst.cc_inst.mux4_1_inst_I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_14_211 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_41_138 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_41_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_497_ _001_ in[0] cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XANTENNA__316__I _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_168 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_26_135 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xro_inst.gcount\[6\].div_flop_inv ro_inst.counter\[6\] ro_inst.counter_n\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_22_396 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_1_235 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_40_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_25_190 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi21_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_351_ _081_ _119_ _120_ _121_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
X_420_ _183_ _186_ _036_ _187_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_282_ _045_ _048_ _049_ _053_ _054_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
XFILLER_0_23_105 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_16_190 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[31\].div_flop_inv ro_inst.counter\[31\] ro_inst.counter_n\[31\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_36_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xro_inst.gcount\[1\].div_flop ro_inst.counter_n\[1\] in[0] ro_inst.counter_n\[0\]
+ ro_inst.counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XANTENNA_cm_inst.cc_inst.dffsnq_4_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_138 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_399 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_208 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.ring_osc_1 ro_inst.ring\[1\] ro_inst.ring\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
X_403_ _049_ _155_ _170_ _127_ _171_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
X_334_ _021_ cm_inst.cc_inst.out_notouch_\[90\] _104_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
XFILLER_0_36_252 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_265_ _036_ _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XTAP_TAPCELL_ROW_47_442 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_6_168 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_42_255 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_42_233 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.clkinv_3_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_506 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_277 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_33_200 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_18_285 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dlyb_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_44_423 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.and2_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai211_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_317_ cm_inst.cc_inst.out_notouch_\[193\] cm_inst.cc_inst.out_notouch_\[201\] _087_
+ _088_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA_cm_inst.cc_inst.dffq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.sdffq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_248_ _019_ _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
Xcm_inst.cc_inst.dffq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[149\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_4
XANTENNA_cm_inst.cc_inst.and4_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_15_222 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_225 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.aoi22_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.nand4_2_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_41_404 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_38_336 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_38_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xro_inst.gcount\[24\].div_flop_inv ro_inst.counter\[24\] ro_inst.counter_n\[24\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_29_336 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.icgtp_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_236 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[2\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai21_1_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_328 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_43_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_380 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_26_297 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SI cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_17_231 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_17_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_17_339 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_0_494 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_110 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__504__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_23_278 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_16_350 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.and3_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_31_397 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_31_386 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_320 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_496_ _000_ in[0] cm_inst.page\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XANTENNA_cm_inst.cc_inst.mux4_1_inst_I2 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_14_212 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_59 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[34\].div_flop ro_inst.counter_n\[34\] in[0] ro_inst.counter_n\[33\]
+ ro_inst.counter\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_1_225 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_49_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.sdffrnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[162\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_17_158 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_375 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_0_291 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
X_350_ _046_ _120_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
Xro_inst.gcount\[17\].div_flop_inv ro_inst.counter\[17\] ro_inst.counter_n\[17\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_281_ _037_ _052_ _053_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
XFILLER_0_8_391 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_39_272 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_479_ _238_ _239_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_22_194 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_10_345 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_378 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__438__S _118_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_33_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_33_415 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_9_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_434 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_13_194 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_36_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.ring_osc_2 ro_inst.ring\[2\] ro_inst.ring\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.aoi21_2_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_264_ _035_ _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
X_402_ _162_ _169_ _017_ _170_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_1
X_333_ _075_ _097_ _099_ _102_ _103_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XFILLER_0_47_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_47_443 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_30_321 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffq_2_inst_SI cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.clkbuf_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[189\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_2
XFILLER_0_37_80 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.dffsnq_1_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dlyd_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[187\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyd_4
XFILLER_0_18_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_33_245 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_33_234 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_21_418 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_191 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_424 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_247_ cm_inst.page\[0\] _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_316_ _082_ _087_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XPHY_EDGE_ROW_26_Left_78 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_24_201 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__281__A1 _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.and4_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_215 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_278 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__250__I cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_11_440 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_46_381 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_21_248 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_195 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.bufz_2_inst_EN cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_7_242 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_220 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xro_inst.gcount\[24\].div_flop ro_inst.counter_n\[24\] in[0] ro_inst.counter_n\[23\]
+ ro_inst.counter\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_38_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_34_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_26_298 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_26_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.buf_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.latrnq_4_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.dffrnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[150\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XTAP_TAPCELL_ROW_17_232 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XPHY_EDGE_ROW_29_Left_81 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_4_256 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[31\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_13_Left_65 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_0_111 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_35_115 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xcm_inst.cc_inst.buf_8_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_8
XFILLER_0_31_310 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.and3_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.or2_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.mux4_1_inst_I3 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_39_390 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_495_ in[4] ro_sel\[2\] _242_ _015_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XTAP_TAPCELL_ROW_14_213 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_22_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.buf_12_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_12
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.or4_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dlyd_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_354 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_280_ _050_ _051_ _033_ _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_31_173 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__298__S0 _063_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_478_ in[1] _238_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_27_446 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_10_368 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xcm_inst.cc_inst.dffnrnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[140\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4
Xro_inst.gcount\[2\].div_flop_inv ro_inst.counter\[2\] ro_inst.counter_n\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_45_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_33_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_490 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_9_189 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_401_ _164_ _166_ _037_ _168_ _169_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
X_263_ cm_inst.page\[3\] _035_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
X_332_ cm_inst.cc_inst.out_notouch_\[194\] cm_inst.cc_inst.out_notouch_\[202\] _101_
+ _102_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA__452__S0 _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__364__S _132_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_47_59 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_47_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_47_444 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.latq_2_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_30_322 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_265 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_27_243 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__248__I _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SI cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.or3_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.or3_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or3_4
XTAP_TAPCELL_ROW_44_425 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_1_Left_53 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_24_224 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_246_ _017_ _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
X_315_ _081_ _085_ cm_inst.cc_inst.out_notouch_\[209\] _086_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand3_1
XTAP_TAPCELL_ROW_9_180 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.and4_4_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_11_430 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_43_Left_95 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_38_305 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[14\].div_flop ro_inst.counter_n\[14\] in[0] ro_inst.counter_n\[13\]
+ ro_inst.counter\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XANTENNA_cm_inst.cc_inst.xnor2_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_44_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_44_319 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_37_360 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_29_316 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_12_196 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_12_238 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_12_227 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_35_319 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_93 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_28_393 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__261__I _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_135 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_26_299 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_34_374 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_34_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_503 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_9_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_17_233 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.xor2_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[60\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor2_1
Xro_inst.gcount\[20\].div_flop_inv ro_inst.counter\[20\] ro_inst.counter_n\[20\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_29_179 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_146 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_124 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai32_4_inst_B1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_40_322 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_396 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.icgtn_1_inst_TE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_0_112 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__457__S _074_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_396 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.or2_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_12_inst_I cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_488 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
X_494_ in[3] ro_sel\[1\] _242_ _014_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XTAP_TAPCELL_ROW_14_214 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_30_Left_82 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_1_216 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_9_338 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.or4_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_40_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_48_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.xnor3_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai221_1_inst_C cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_39_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__298__S1 _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_477_ in[4] _111_ _236_ _002_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_27_414 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.invz_3_inst_I cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_61 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_42_93 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_342 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_SI cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_33_417 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_400_ _110_ _167_ _168_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
X_331_ _100_ _101_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_36_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.nor3_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_262_ _033_ _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
Xcm_inst.cc_inst.aoi21_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[67\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_2
XTAP_TAPCELL_ROW_47_445 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_47_38 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xro_inst.gcount\[13\].div_flop_inv ro_inst.counter\[13\] ro_inst.counter_n\[13\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_2_18 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.latq_2_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_42_236 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_42_225 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_323 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_23_483 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_SETN cm_inst.cc_inst.in\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.or3_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_461 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__375__S _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_314_ _084_ _085_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
X_245_ cm_inst.page\[4\] _017_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_236 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_15_236 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_239 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai221_4_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_11_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_38_328 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__507__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__407__S1 _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_501 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_ro_inst.gcount\[27\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_18 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.xnor2_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_12_197 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.sdffrnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[164\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4
XFILLER_0_47_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_31_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_28_372 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_233 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_222 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_3_132 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nor4_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_ro_inst.gcount\[15\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_372 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_19_394 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__401__B _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_234 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_40_312 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_37_180 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_342 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai32_4_inst_B2 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai32_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__483__I0 in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_113 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_48_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_31_323 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi221_1_inst_C cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_493_ in[2] _225_ _242_ _013_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
Xcm_inst.cc_inst.hold_inst cm_inst.cc_inst.out_notouch_\[173\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__hold
XFILLER_0_26_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_22_270 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_14_215 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_34_183 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_378 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_1_239 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_45_415 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_31_62 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_13_323 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.or4_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.mux2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[118\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_2
XFILLER_0_0_283 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_378 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_28_307 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__267__I cm_inst.page\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.xnor3_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_31_120 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_16_194 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_476_ in[3] _107_ _236_ _001_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_50_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_33_343 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_9_158 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_470 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai31_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[33\].div_flop ro_inst.counter_n\[33\] in[0] ro_inst.counter_n\[32\]
+ ro_inst.counter\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
X_330_ _026_ _100_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_36_256 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nor3_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_261_ _032_ _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrnq_2_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_47_446 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_30_324 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_459_ _018_ _215_ _223_ _058_ _224_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi211_1
Xcm_inst.cc_inst.dlya_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[177\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlya_2
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_10_123 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_10_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.inv_16_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_16
XFILLER_0_5_150 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or3_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_289 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_244_ ro_inst.enable _016_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
X_313_ _083_ _084_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
XFILLER_0_20_432 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dffrnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[152\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_4
XFILLER_0_23_52 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_15_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_207 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.oai221_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai221_4_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.xor3_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_11_410 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_443 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_307 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_40_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xro_inst.clock_gate ro_inst.ring\[0\] ro_inst.running _243_ ro_inst.counter\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__icgtp_1
XTAP_TAPCELL_ROW_12_198 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_12_229 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_43_354 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_43_310 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.nor4_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.icgtp_1_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_3_133 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_17_235 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.addf_2_inst_A cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_25_290 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_25_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai32_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_40_368 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__483__I1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_0_114 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_48_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_16_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_31_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_302 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnq_4_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_413 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_492_ in[5] in[6] in[7] in[1] _242_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand4_1
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_22_271 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.aoi222_1_inst_C1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.sdffq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[160\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffq_2
XFILLER_0_1_218 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.bufz_1_inst_I cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_17_Left_69 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.or4_4_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.invz_12_inst cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[175\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__invz_12
XFILLER_0_13_302 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xro_inst.gcount\[23\].div_flop ro_inst.counter_n\[23\] in[0] ro_inst.counter_n\[22\]
+ ro_inst.counter\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_36_363 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_28_308 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.xnor3_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_31_187 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.clkbuf_16_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[194\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_16
Xcm_inst.cc_inst.oai32_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[91\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai32_2
X_475_ in[2] _042_ _237_ _000_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_27_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__455__S0 _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_22_143 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_2_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffrsnq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SE cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.inv_20_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__368__I _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_33_344 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_26_482 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai31_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_260_ cm_inst.page\[2\] _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
Xcm_inst.cc_inst.inv_3_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_3
XFILLER_0_8_181 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nor3_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_30_325 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_458_ _059_ _222_ _223_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_389_ _085_ cm_inst.cc_inst.out_notouch_\[84\] _156_ _105_ _157_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi211_1
XFILLER_0_2_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.clkinv_16_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_33_238 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_312_ _082_ _083_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_32_260 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__471__I in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_249 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_17_290 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.xor2_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[62\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor2_4
XANTENNA_cm_inst.cc_inst.aoi221_2_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_15_216 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_15_205 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai221_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.xor3_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_500 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_5_Left_57 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_6_153 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_37_374 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_341 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_12_199 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.dffsnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_85 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_7_246 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_235 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_47_Left_99 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_3_134 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nor4_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_127 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_34_322 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_399 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__397__S _118_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_25_291 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_17_236 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_40_303 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.addf_2_inst_B cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_333 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai32_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[13\].div_flop ro_inst.counter_n\[13\] in[0] ro_inst.counter_n\[12\]
+ ro_inst.counter\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_115 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_0_104 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_31_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_260 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.sig_latch ro_inst.signal ro_inst.slow_clk_n ro_inst.saved_signal vdd vdd
+ vss vss gf180mcu_fd_sc_mcu9t5v0__latq_1
XANTENNA_cm_inst.cc_inst.buf_12_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_491_ _241_ _012_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.aoi222_1_inst_C2 cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_1_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_34_141 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_30_380 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_8_Left_60 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_40_188 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_174 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_13_369 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_28_309 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_36_364 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_8_330 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_34_Left_86 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.oai22_4_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_233 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_474_ _236_ _237_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XANTENNA__455__S1 _122_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.or4_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or4_1
XFILLER_0_42_41 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_33_345 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_ro_inst.gcount\[7\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_5_300 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai31_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_41_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.invz_2_inst_EN cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.addh_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[111\]
+ cm_inst.cc_inst.out_notouch_\[112\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__addh_1
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_51_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_8_193 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XANTENNA_cm_inst.cc_inst.nand3_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_30_326 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_388_ _021_ cm_inst.cc_inst.out_notouch_\[92\] _156_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
X_457_ _218_ _221_ _074_ _222_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XANTENNA_cm_inst.cc_inst.dlyc_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_41_294 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_152 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__289__I _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_311_ cm_inst.page\[0\] _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XFILLER_0_32_272 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi221_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi221_2_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_501 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_509_ _013_ in[0] ro_sel\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XPHY_EDGE_ROW_21_Left_73 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xcm_inst.cc_inst.latrsnq_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[129\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latrsnq_1
XANTENNA_cm_inst.cc_inst.xor3_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_11_434 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_478 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.sdffq_1_inst_SE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.addf_2_inst_CI cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.icgtn_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[204\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__icgtn_1
XTAP_TAPCELL_ROW_6_154 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__495__I0 in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrsnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_231 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_97 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_258 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_225 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_3_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.clkbuf_8_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[192\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_8
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__486__I0 in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_3_135 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nor4_1_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_22_507 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nand4_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__477__I0 in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.clkinv_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_25_292 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_40_326 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.dffq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_0_116 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_0_105 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_3_272 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.aoi22_4_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_39_384 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_490_ _238_ _016_ _236_ _241_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XANTENNA_cm_inst.cc_inst.aoi222_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_1_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.clock_gate_inv ro_inst.counter\[0\] ro_inst.counter_n\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_38_470 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_10 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_13_326 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffrsnq_4_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__302__A2 _072_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_0_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_365 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_44_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.oai22_4_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai22_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_473_ _233_ _234_ _235_ in[1] _236_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai31_1
XFILLER_0_39_278 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_27_418 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai21_2_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_22_123 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.nor2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[37\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor2_2
XTAP_TAPCELL_ROW_33_346 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.mux2_2_inst_I0 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.nand2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_2
Xro_inst.gcount\[9\].div_flop_inv ro_inst.counter\[9\] ro_inst.counter_n\[9\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.mux4_4_inst_I0 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.nand3_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_456_ _219_ _220_ _182_ _221_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XTAP_TAPCELL_ROW_30_327 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_27_259 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_387_ _075_ _152_ _153_ _154_ _155_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_23_487 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_53 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_5_197 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_14_410 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_465 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_44_419 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_310_ _078_ _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
Xro_inst.gcount\[34\].div_flop_inv ro_inst.counter\[34\] ro_inst.counter_n\[34\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.invz_12_inst_I cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_32_295 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_174 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.aoi221_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_424 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai21_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_ro_inst.gcount\[24\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[32\].div_flop ro_inst.counter_n\[32\] in[0] ro_inst.counter_n\[31\]
+ ro_inst.counter\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
X_508_ _012_ in[0] ro_inst.enable vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
X_439_ _081_ _204_ _120_ _205_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_1
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_6_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SE cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_251 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_6_155 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_37_343 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_37_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.buf_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_20_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[12\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_302 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_28_376 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_190 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__486__I1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_3_136 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_49_Left_101 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.nand4_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai211_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_37_184 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_25_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_40_305 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_33_390 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_43 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA__442__B _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_76 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_0_117 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_0_106 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.aoi22_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi22_4_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.oai21_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[82\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai21_2
XFILLER_0_39_405 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_39_385 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[27\].div_flop_inv ro_inst.counter\[27\] ro_inst.counter_n\[27\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.aoi222_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_382 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.latrsnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_45_419 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_25_198 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_305 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_0_210 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_0_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_0_287 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA__510__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_36_366 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_8_310 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_321 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_179 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_146 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_198 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai22_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_202 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
X_472_ in[7] _235_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
XTAP_TAPCELL_ROW_27_300 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_35_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.invz_3_inst cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[174\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__invz_3
Xcm_inst.cc_inst.sdffrsnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\]
+ cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[166\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2
XTAP_TAPCELL_ROW_33_347 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.buf_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_474 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.mux2_2_inst_I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_36_249 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_8_195 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.and3_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_496 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrsnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi21_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[22\].div_flop ro_inst.counter_n\[22\] in[0] ro_inst.counter_n\[21\]
+ ro_inst.counter\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XANTENNA_cm_inst.cc_inst.mux4_4_inst_I1 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_386_ _099_ _154_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XANTENNA_cm_inst.cc_inst.nand3_2_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_455_ cm_inst.cc_inst.out_notouch_\[7\] cm_inst.cc_inst.out_notouch_\[15\] cm_inst.cc_inst.out_notouch_\[23\]
+ cm_inst.cc_inst.out_notouch_\[31\] _020_ _122_ _220_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.clkbuf_20_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_50_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.icgtp_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[208\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__icgtp_2
XFILLER_0_33_208 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_238 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_41_296 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_41_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_SE cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA__291__S1 _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_32_274 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.bufz_2_inst cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[171\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_2
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_175 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai21_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_507_ _011_ in[0] cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
X_438_ cm_inst.cc_inst.out_notouch_\[6\] cm_inst.cc_inst.out_notouch_\[14\] _118_
+ _204_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_369_ _064_ _138_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_11_414 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_46_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__355__B _074_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_14_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_14_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_6_156 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.and2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_2
XANTENNA_cm_inst.cc_inst.and2_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_34_99 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_28_300 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_238 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_216 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_191 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_11_222 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_137 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_311 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nand4_1_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrnq_1_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai211_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.or4_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__or4_4
XFILLER_0_29_99 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_0_107 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xcm_inst.cc_inst.addh_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[115\]
+ cm_inst.cc_inst.out_notouch_\[116\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__addh_4
XANTENNA_cm_inst.cc_inst.aoi22_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_39_417 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_39_386 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_14_209 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_34_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_188 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.dffrnq_4_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_461 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_200 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_233 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_244 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_299 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_367 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.xnor2_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.out_notouch_\[55\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xnor2_2
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_31_169 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.invz_12_inst_EN cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_27_301 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_471_ in[6] _234_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
Xro_inst.gcount\[12\].div_flop ro_inst.counter_n\[12\] in[0] ro_inst.counter_n\[11\]
+ ro_inst.counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_50_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SI cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_45 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_45_206 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_42_77 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_33_348 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__367__S0 _063_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.latrsnq_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[131\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latrsnq_4
Xcm_inst.cc_inst.xor3_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor3_1
XANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
Xcm_inst.cc_inst.icgtn_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[206\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__icgtn_4
XFILLER_0_8_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.and3_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.clkinv_20_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[203\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_20
XFILLER_0_12_191 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi21_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.mux4_4_inst_I2 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_27_239 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_385_ cm_inst.cc_inst.out_notouch_\[196\] cm_inst.cc_inst.out_notouch_\[204\] _101_
+ _153_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_454_ cm_inst.cc_inst.out_notouch_\[39\] cm_inst.cc_inst.out_notouch_\[47\] cm_inst.cc_inst.out_notouch_\[55\]
+ cm_inst.cc_inst.out_notouch_\[63\] _179_ _180_ _219_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA__500__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_23_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_23_401 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_41_220 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_5_155 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_41_275 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_41_286 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_32_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_176 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_506_ _010_ in[0] cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XANTENNA_cm_inst.cc_inst.dffnsnq_4_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_299_ cm_inst.cc_inst.out_notouch_\[1\] cm_inst.cc_inst.out_notouch_\[9\] cm_inst.cc_inst.out_notouch_\[17\]
+ cm_inst.cc_inst.out_notouch_\[25\] _063_ _065_ _070_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_368_ _082_ _137_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
Xro_inst.gcount\[5\].div_flop_inv ro_inst.counter\[5\] ro_inst.counter_n\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
X_437_ _084_ cm_inst.cc_inst.out_notouch_\[22\] _202_ _105_ _203_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi211_1
XFILLER_0_23_231 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_15_209 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_2_147 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_426 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai221_2_inst_C cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.icgtn_4_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_504 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.invz_4_inst_I cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__489__I0 in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_6_157 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_37_378 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.and2_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_278 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XPHY_EDGE_ROW_25_Left_77 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.dffnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[30\].div_flop_inv ro_inst.counter\[30\] ro_inst.counter_n\[30\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_28_323 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_312 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_412 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_192 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.aoi22_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[70\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_2
XTAP_TAPCELL_ROW_3_138 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.aoi211_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_34_326 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nand4_1_inst_A4 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xcm_inst.cc_inst.oai31_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[87\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai31_1
XFILLER_0_25_337 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_67 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_78 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_108 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_31_318 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_24_381 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnsnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_3_275 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_3_264 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_387 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_34_145 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[9\].div_flop ro_inst.counter_n\[9\] in[0] ro_inst.counter_n\[8\]
+ ro_inst.counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_22_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_22_265 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_19_186 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_440 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_31_46 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xcm_inst.cc_inst.dffnq_1_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[135\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnq_1
XTAP_TAPCELL_ROW_36_368 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XPHY_EDGE_ROW_28_Left_80 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_8_312 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_8_334 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_12_Left_64 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_16_167 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[4\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.clkinv_3_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[198\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_3
XTAP_TAPCELL_ROW_27_302 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_470_ in[5] _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkinv_1
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xro_inst.gcount\[23\].div_flop_inv ro_inst.counter\[23\] ro_inst.counter_n\[23\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_42_45 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_26_421 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_410 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_5_304 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_21_181 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_49_460 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.and3_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_12_170 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.mux4_4_inst_I3 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_453_ _216_ _217_ _182_ _218_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_27_207 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_384_ _148_ _151_ _132_ _152_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_23_413 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
Xcm_inst.cc_inst.buf_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_4
XANTENNA_cm_inst.cc_inst.aoi221_2_inst_C cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_46_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_26_251 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.icgtn_2_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_20_405 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_20_449 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_177 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_505_ _009_ in[0] cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XFILLER_0_28_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_23_14 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
X_436_ _100_ cm_inst.cc_inst.out_notouch_\[30\] _202_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__and2_1
XFILLER_0_43_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_298_ cm_inst.cc_inst.out_notouch_\[33\] cm_inst.cc_inst.out_notouch_\[41\] cm_inst.cc_inst.out_notouch_\[49\]
+ cm_inst.cc_inst.out_notouch_\[57\] _063_ _061_ _069_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_367_ cm_inst.cc_inst.out_notouch_\[99\] cm_inst.cc_inst.out_notouch_\[107\] cm_inst.cc_inst.out_notouch_\[115\]
+ cm_inst.cc_inst.out_notouch_\[123\] _063_ _065_ _136_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA__498__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_23_298 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_438 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffq_1_inst_SI cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.latrsnq_4_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__489__I1 cm_inst.cc_inst.in\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_6_158 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_37_313 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_368 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_37_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xro_inst.gcount\[16\].div_flop_inv ro_inst.counter\[16\] ro_inst.counter_n\[16\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XPHY_EDGE_ROW_0_Left_52 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_20_235 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_28_335 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_7_207 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_419_ _184_ _185_ _182_ _186_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XTAP_TAPCELL_ROW_11_193 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.buf_8_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi211_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_368 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_42_Left_94 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
Xro_inst.gcount\[31\].div_flop ro_inst.counter_n\[31\] in[0] ro_inst.counter_n\[30\]
+ ro_inst.counter\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
Xcm_inst.cc_inst.dlyb_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[180\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dlyb_2
XANTENNA_cm_inst.cc_inst.or3_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffsnq_4_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_40_319 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_40_308 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_21_500 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_109 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.oai211_1_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_28_187 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_28_132 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_8_505 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_24_393 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.bufz_1_inst_EN cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_39_388 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.oai221_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[100\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai221_2
XFILLER_0_19_154 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_22_266 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_474 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_38_463 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_5_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_0_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_36_369 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_441 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_27_303 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA__327__S _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffsnq_4_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_22_127 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or2_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.icgtp_2_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.sdffq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dlya_4_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.icgtn_4_inst_TE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai31_4_inst_B cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_44_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.sdffq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_271 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_143 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_ro_inst.gcount\[33\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_32_403 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_198 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
X_383_ cm_inst.cc_inst.out_notouch_\[132\] cm_inst.cc_inst.out_notouch_\[140\] cm_inst.cc_inst.out_notouch_\[148\]
+ cm_inst.cc_inst.out_notouch_\[156\] _149_ _150_ _151_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
X_452_ cm_inst.cc_inst.out_notouch_\[71\] cm_inst.cc_inst.out_notouch_\[79\] cm_inst.cc_inst.out_notouch_\[87\]
+ cm_inst.cc_inst.out_notouch_\[95\] _020_ _180_ _217_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_41_299 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.latsnq_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[133\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__latsnq_2
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_14_414 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_RN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.icgtp_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_ro_inst.gcount\[21\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.bufz_2_inst_I cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_32_211 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_17_230 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.xnor3_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_4_190 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_9_178 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_20_428 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_43_412 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_504_ _008_ in[0] cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
X_435_ _196_ _198_ _047_ _200_ _201_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai211_1
X_366_ _075_ _133_ _134_ _099_ _135_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
X_297_ _062_ _066_ _067_ _068_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_23_277 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
Xcm_inst.cc_inst.oai33_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.in\[5\] cm_inst.cc_inst.out_notouch_\[94\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai33_2
XANTENNA_cm_inst.cc_inst.latrsnq_4_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[21\].div_flop ro_inst.counter_n\[21\] in[0] ro_inst.counter_n\[20\]
+ ro_inst.counter\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_10_461 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_14_233 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.sdffsnq_1_inst_SI cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_6_159 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_37_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_271 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.aoi211_1_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_306 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_314 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_349_ cm_inst.cc_inst.out_notouch_\[2\] cm_inst.cc_inst.out_notouch_\[10\] _118_
+ _119_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
X_418_ cm_inst.cc_inst.out_notouch_\[5\] cm_inst.cc_inst.out_notouch_\[13\] cm_inst.cc_inst.out_notouch_\[21\]
+ cm_inst.cc_inst.out_notouch_\[29\] _020_ _122_ _185_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XTAP_TAPCELL_ROW_11_194 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[1\].div_flop_inv ro_inst.counter\[1\] ro_inst.counter_n\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XTAP_TAPCELL_ROW_19_250 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.inv_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.or3_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_10_291 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_25_339 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_25_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_25_286 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_33_394 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_33_383 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.xnor2_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_28_111 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai211_1_inst_C cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_43_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.xor3_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[65\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__xor3_4
XTAP_TAPCELL_ROW_39_389 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_39_409 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_47_486 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_267 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_188 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA__412__I _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_420 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__503__CLK in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_0_214 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.nor2_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_320 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.latsnq_1_inst_D cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_44_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SETN cm_inst.cc_inst.in\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_12_331 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_147 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_39_228 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_27_304 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nor4_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_35_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.or2_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.icgtp_2_inst_TE cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.mux2_1_inst_S cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_478 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai222_2_inst_C1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_32_340 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_32_459 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_382_ _061_ _150_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XFILLER_0_27_209 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_451_ cm_inst.cc_inst.out_notouch_\[103\] cm_inst.cc_inst.out_notouch_\[111\] cm_inst.cc_inst.out_notouch_\[119\]
+ cm_inst.cc_inst.out_notouch_\[127\] _179_ _138_ _216_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_2_309 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_37_14 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_14_404 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
Xcm_inst.cc_inst.aoi221_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.in\[4\] cm_inst.cc_inst.out_notouch_\[76\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi221_2
XFILLER_0_41_234 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
Xro_inst.gcount\[11\].div_flop ro_inst.counter_n\[11\] in[0] ro_inst.counter_n\[10\]
+ ro_inst.counter\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XFILLER_0_27_80 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.sdffrnq_1_inst_SI cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_442 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.xnor3_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_17_297 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.clkbuf_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[188\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
XTAP_TAPCELL_ROW_9_179 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
X_503_ _007_ in[0] cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XANTENNA_cm_inst.cc_inst.nor3_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_43_413 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.oai31_4_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[89\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai31_4
X_296_ _032_ _067_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_434_ _111_ _199_ _200_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand2_1
X_365_ cm_inst.cc_inst.out_notouch_\[195\] cm_inst.cc_inst.out_notouch_\[203\] _101_
+ _134_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_2_139 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_11_418 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai33_2_inst_B1 cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_489 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.oai31_4_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_10_451 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.latsnq_2_inst_SETN cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_37_337 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_34_26 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_28_304 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi211_1_inst_C cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
X_348_ _060_ _118_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
X_279_ cm_inst.cc_inst.out_notouch_\[128\] cm_inst.cc_inst.out_notouch_\[136\] cm_inst.cc_inst.out_notouch_\[144\]
+ cm_inst.cc_inst.out_notouch_\[152\] _027_ _023_ _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
Xcm_inst.cc_inst.dffnq_4_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[137\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnq_4
XANTENNA__325__I _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_417_ cm_inst.cc_inst.out_notouch_\[37\] cm_inst.cc_inst.out_notouch_\[45\] cm_inst.cc_inst.out_notouch_\[53\]
+ cm_inst.cc_inst.out_notouch_\[61\] _179_ _180_ _184_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_11_226 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_19_315 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA_cm_inst.cc_inst.or3_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__492__A1 in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_2_130 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.inv_12_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_12
XANTENNA_cm_inst.cc_inst.dlyc_2_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_33_340 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_329 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_25_287 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_29_59 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.xnor2_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xro_inst.gcount\[12\].div_flop_inv ro_inst.counter\[12\] ro_inst.counter_n\[12\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu9t5v0__inv_1
XANTENNA_cm_inst.cc_inst.addh_1_inst_A cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_24_395 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_3_256 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_502 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_35_80 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_34_137 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_22_268 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_38_443 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_38_432 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_202 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_ro_inst.gcount\[29\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_33_192 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_0_248 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_cm_inst.cc_inst.nor2_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_CLKN cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.latsnq_1_inst_E cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_29_443 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_410 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_12_310 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.nor4_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffrsnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XTAP_TAPCELL_ROW_35_360 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XTAP_TAPCELL_ROW_27_305 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_35_468 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_22_129 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XANTENNA_ro_inst.gcount\[17\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.dffnrnq_1_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_251 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_26_402 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XANTENNA_cm_inst.cc_inst.oai222_2_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai222_2_inst_C2 cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_173 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xro_inst.gcount\[8\].div_flop ro_inst.counter_n\[8\] in[0] ro_inst.counter_n\[7\]
+ ro_inst.counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XPHY_EDGE_ROW_16_Left_68 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_44_265 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_32_341 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_32_427 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_29_273 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_17_413 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_4_384 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_12_195 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.xor2_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_381_ _060_ _149_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__buf_1
X_450_ _172_ _213_ _214_ _154_ _215_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi22_1
XFILLER_0_23_416 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.aoi222_4_inst_C1 cm_inst.cc_inst.in\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_46_433 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA__328__I _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_276 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_41_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_49_346 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_37_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.xnor3_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_9_487 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_13_460 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_43_414 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_502_ _006_ in[0] cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffq_1
XANTENNA__349__S _118_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_433_ cm_inst.cc_inst.out_notouch_\[102\] cm_inst.cc_inst.out_notouch_\[110\] cm_inst.cc_inst.out_notouch_\[118\]
+ cm_inst.cc_inst.out_notouch_\[126\] _087_ _112_ _199_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA_cm_inst.cc_inst.nor3_1_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_51_480 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
X_295_ cm_inst.cc_inst.out_notouch_\[65\] cm_inst.cc_inst.out_notouch_\[73\] cm_inst.cc_inst.out_notouch_\[81\]
+ cm_inst.cc_inst.out_notouch_\[89\] _063_ _065_ _066_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XANTENNA__424__S0 _130_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_2_inst_B2 cm_inst.cc_inst.in\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai33_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
X_364_ _129_ _131_ _132_ _133_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_31_290 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_23_235 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
Xcm_inst.cc_inst.clkbuf_12_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.out_notouch_\[193\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__clkbuf_12
XANTENNA_cm_inst.cc_inst.clkbuf_1_inst_I cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_19_508 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.oai31_4_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_32
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XFILLER_0_1_173 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_10_441 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.nor3_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nor3_2
XPHY_EDGE_ROW_19_Left_71 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XANTENNA__406__S0 _130_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_33_500 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.dffnsnq_2_inst cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[0\]
+ cm_inst.cc_inst.out_notouch_\[145\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2
XFILLER_0_9_251 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_9_273 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XTAP_TAPCELL_ROW_5_150 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.nand3_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__nand3_2
X_416_ _178_ _181_ _182_ _183_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux2_1
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
X_347_ _084_ cm_inst.cc_inst.out_notouch_\[18\] _116_ _039_ _117_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__aoi211_1
X_278_ cm_inst.cc_inst.out_notouch_\[160\] cm_inst.cc_inst.out_notouch_\[168\] cm_inst.cc_inst.out_notouch_\[176\]
+ cm_inst.cc_inst.out_notouch_\[184\] _027_ _023_ _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_34_319 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XANTENNA_cm_inst.cc_inst.xor3_1_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__251__I _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA__492__A2 in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_2_131 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_10_282 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XPHY_EDGE_ROW_4_Left_56 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_37_135 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_288 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xcm_inst.cc_inst.bufz_8_inst cm_inst.cc_inst.in\[2\] cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[172\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__bufz_8
XFILLER_0_18_371 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XANTENNA_cm_inst.cc_inst.addh_1_inst_B cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.latrsnq_2_inst_SETN cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_3_268 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_46_Left_98 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_34_127 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_269 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XFILLER_0_19_146 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_42_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_30_300 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.bufz_8_inst_I cm_inst.cc_inst.in\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_38_466 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XTAP_TAPCELL_ROW_38_380 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_ro_inst.gcount\[1\].div_flop_RN in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_13_203 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
Xro_inst.gcount\[30\].div_flop ro_inst.counter_n\[30\] in[0] ro_inst.counter_n\[29\]
+ ro_inst.counter\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
XANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_D cm_inst.cc_inst.in\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_8_327 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XFILLER_0_24_193 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_8
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_16
XTAP_TAPCELL_ROW_27_306 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.nor4_4_inst_A3 cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XTAP_TAPCELL_ROW_35_361 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.aoi21_4_inst_B cm_inst.cc_inst.in\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_30_174 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_30_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_26_425 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA_cm_inst.cc_inst.oai222_2_inst_A1 cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.oai222_2_inst_B2 cm_inst.cc_inst.in\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_21_185 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_21_196 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_1
XFILLER_0_29_241 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_25_480 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_12_163 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XANTENNA_cm_inst.cc_inst.xor2_2_inst_A2 cm_inst.cc_inst.in\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_4_inst_B1 cm_inst.cc_inst.in\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XANTENNA_cm_inst.cc_inst.aoi222_4_inst_C2 cm_inst.cc_inst.in\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
X_380_ cm_inst.cc_inst.out_notouch_\[164\] cm_inst.cc_inst.out_notouch_\[172\] cm_inst.cc_inst.out_notouch_\[180\]
+ cm_inst.cc_inst.out_notouch_\[188\] _130_ _095_ _148_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__mux4_1
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_64
XPHY_EDGE_ROW_33_Left_85 vdd vss gf180mcu_fd_sc_mcu9t5v0__endcap
XFILLER_0_7_190 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XFILLER_0_16_480 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
Xcm_inst.cc_inst.oai22_2_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.in\[3\] cm_inst.cc_inst.out_notouch_\[85\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__oai22_2
XTAP_TAPCELL_ROW_46_434 vdd vss gf180mcu_fd_sc_mcu9t5v0__filltie
XANTENNA_cm_inst.cc_inst.dffrnq_2_inst_CLK cm_inst.cc_inst.in\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu9t5v0__antenna
XFILLER_0_26_255 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fillcap_4
XFILLER_0_22_461 vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__fill_2
XANTENNA__280__S _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__antenna
Xcm_inst.cc_inst.aoi21_1_inst cm_inst.cc_inst.in\[0\] cm_inst.cc_inst.in\[1\] cm_inst.cc_inst.in\[2\]
+ cm_inst.cc_inst.out_notouch_\[66\] vdd vdd vss vss gf180mcu_fd_sc_mcu9t5v0__aoi21_1
.ends

