magic
tech gf180mcuD
magscale 1 5
timestamp 1702442008
<< obsm1 >>
rect 672 1538 59304 48313
<< metal2 >>
rect 26208 49600 26264 50000
rect 26544 49600 26600 50000
rect 27216 49600 27272 50000
rect 27888 49600 27944 50000
rect 28560 49600 28616 50000
rect 28896 49600 28952 50000
rect 29232 49600 29288 50000
rect 29904 49600 29960 50000
rect 30912 49600 30968 50000
rect 31248 49600 31304 50000
rect 31584 49600 31640 50000
rect 31920 49600 31976 50000
rect 32256 49600 32312 50000
rect 0 0 56 400
rect 336 0 392 400
rect 672 0 728 400
rect 1008 0 1064 400
rect 1344 0 1400 400
rect 1680 0 1736 400
rect 2016 0 2072 400
rect 2352 0 2408 400
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 26880 0 26936 400
rect 31248 0 31304 400
rect 31584 0 31640 400
rect 31920 0 31976 400
<< obsm2 >>
rect 462 49570 26178 49600
rect 26294 49570 26514 49600
rect 26630 49570 27186 49600
rect 27302 49570 27858 49600
rect 27974 49570 28530 49600
rect 28646 49570 28866 49600
rect 28982 49570 29202 49600
rect 29318 49570 29874 49600
rect 29990 49570 30882 49600
rect 30998 49570 31218 49600
rect 31334 49570 31554 49600
rect 31670 49570 31890 49600
rect 32006 49570 32226 49600
rect 32342 49570 59122 49600
rect 462 430 59122 49570
rect 462 350 642 430
rect 758 350 978 430
rect 1094 350 1314 430
rect 1430 350 1650 430
rect 1766 350 1986 430
rect 2102 350 2322 430
rect 2438 350 2658 430
rect 2774 350 2994 430
rect 3110 350 3330 430
rect 3446 350 26850 430
rect 26966 350 31218 430
rect 31334 350 31554 430
rect 31670 350 31890 430
rect 32006 350 59122 430
<< metal3 >>
rect 0 40992 400 41048
rect 59600 24864 60000 24920
rect 0 22848 400 22904
rect 0 22512 400 22568
<< obsm3 >>
rect 400 41078 59600 48230
rect 430 40962 59600 41078
rect 400 24950 59600 40962
rect 400 24834 59570 24950
rect 400 22934 59600 24834
rect 430 22818 59600 22934
rect 400 22598 59600 22818
rect 430 22482 59600 22598
rect 400 1554 59600 22482
<< metal4 >>
rect 2224 1538 2384 48246
rect 9904 1538 10064 48246
rect 17584 1538 17744 48246
rect 25264 1538 25424 48246
rect 32944 1538 33104 48246
rect 40624 1538 40784 48246
rect 48304 1538 48464 48246
rect 55984 1538 56144 48246
<< obsm4 >>
rect 1806 1801 2194 42887
rect 2414 1801 9874 42887
rect 10094 1801 17554 42887
rect 17774 1801 25234 42887
rect 25454 1801 32914 42887
rect 33134 1801 40594 42887
rect 40814 1801 48274 42887
rect 48494 1801 52850 42887
<< labels >>
rlabel metal3 s 0 40992 400 41048 6 clk
port 1 nsew signal input
rlabel metal2 s 27216 49600 27272 50000 6 in[0]
port 2 nsew signal input
rlabel metal2 s 0 0 56 400 6 in[10]
port 3 nsew signal input
rlabel metal2 s 336 0 392 400 6 in[11]
port 4 nsew signal input
rlabel metal2 s 672 0 728 400 6 in[12]
port 5 nsew signal input
rlabel metal2 s 1008 0 1064 400 6 in[13]
port 6 nsew signal input
rlabel metal2 s 1344 0 1400 400 6 in[14]
port 7 nsew signal input
rlabel metal2 s 1680 0 1736 400 6 in[15]
port 8 nsew signal input
rlabel metal2 s 2016 0 2072 400 6 in[16]
port 9 nsew signal input
rlabel metal2 s 2352 0 2408 400 6 in[17]
port 10 nsew signal input
rlabel metal2 s 26544 49600 26600 50000 6 in[1]
port 11 nsew signal input
rlabel metal2 s 26208 49600 26264 50000 6 in[2]
port 12 nsew signal input
rlabel metal3 s 0 22512 400 22568 6 in[3]
port 13 nsew signal input
rlabel metal3 s 0 22848 400 22904 6 in[4]
port 14 nsew signal input
rlabel metal2 s 26880 0 26936 400 6 in[5]
port 15 nsew signal input
rlabel metal2 s 28896 49600 28952 50000 6 in[6]
port 16 nsew signal input
rlabel metal2 s 2688 0 2744 400 6 in[7]
port 17 nsew signal input
rlabel metal2 s 3024 0 3080 400 6 in[8]
port 18 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 in[9]
port 19 nsew signal input
rlabel metal2 s 31248 0 31304 400 6 out[0]
port 20 nsew signal output
rlabel metal2 s 28560 49600 28616 50000 6 out[10]
port 21 nsew signal output
rlabel metal2 s 32256 49600 32312 50000 6 out[11]
port 22 nsew signal output
rlabel metal2 s 31584 0 31640 400 6 out[1]
port 23 nsew signal output
rlabel metal3 s 59600 24864 60000 24920 6 out[2]
port 24 nsew signal output
rlabel metal2 s 31920 0 31976 400 6 out[3]
port 25 nsew signal output
rlabel metal2 s 31248 49600 31304 50000 6 out[4]
port 26 nsew signal output
rlabel metal2 s 31584 49600 31640 50000 6 out[5]
port 27 nsew signal output
rlabel metal2 s 31920 49600 31976 50000 6 out[6]
port 28 nsew signal output
rlabel metal2 s 30912 49600 30968 50000 6 out[7]
port 29 nsew signal output
rlabel metal2 s 29904 49600 29960 50000 6 out[8]
port 30 nsew signal output
rlabel metal2 s 29232 49600 29288 50000 6 out[9]
port 31 nsew signal output
rlabel metal2 s 27888 49600 27944 50000 6 rst_n
port 32 nsew signal input
rlabel metal4 s 2224 1538 2384 48246 6 vdd
port 33 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 48246 6 vdd
port 33 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 48246 6 vdd
port 33 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 48246 6 vdd
port 33 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 48246 6 vss
port 34 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 48246 6 vss
port 34 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 48246 6 vss
port 34 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 48246 6 vss
port 34 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6172208
string GDS_FILE /home/htamas/progs/gfmpw1-multi.v2/openlane/totp/runs/23_12_13_05_26/results/signoff/totp.magic.gds
string GDS_START 376876
<< end >>

