magic
tech gf180mcuD
magscale 1 10
timestamp 1702441927
<< metal1 >>
rect 1344 44714 46592 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 46592 44714
rect 1344 44628 46592 44662
rect 1344 43930 46592 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 46592 43930
rect 1344 43844 46592 43878
rect 1710 43762 1762 43774
rect 28354 43710 28366 43762
rect 28418 43710 28430 43762
rect 1710 43698 1762 43710
rect 30494 43650 30546 43662
rect 13234 43598 13246 43650
rect 13298 43598 13310 43650
rect 28242 43598 28254 43650
rect 28306 43598 28318 43650
rect 30494 43586 30546 43598
rect 29486 43538 29538 43550
rect 13010 43486 13022 43538
rect 13074 43486 13086 43538
rect 19170 43486 19182 43538
rect 19234 43486 19246 43538
rect 25330 43486 25342 43538
rect 25394 43486 25406 43538
rect 26114 43486 26126 43538
rect 26178 43486 26190 43538
rect 29486 43474 29538 43486
rect 30830 43538 30882 43550
rect 30830 43474 30882 43486
rect 25790 43426 25842 43438
rect 19842 43374 19854 43426
rect 19906 43374 19918 43426
rect 22306 43374 22318 43426
rect 22370 43374 22382 43426
rect 28690 43374 28702 43426
rect 28754 43374 28766 43426
rect 25790 43362 25842 43374
rect 27246 43314 27298 43326
rect 27246 43250 27298 43262
rect 30270 43314 30322 43326
rect 30270 43250 30322 43262
rect 1344 43146 46592 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 46592 43146
rect 1344 43060 46592 43094
rect 20078 42754 20130 42766
rect 22430 42754 22482 42766
rect 13570 42702 13582 42754
rect 13634 42702 13646 42754
rect 14914 42702 14926 42754
rect 14978 42702 14990 42754
rect 21970 42702 21982 42754
rect 22034 42702 22046 42754
rect 22866 42702 22878 42754
rect 22930 42702 22942 42754
rect 23314 42702 23326 42754
rect 23378 42702 23390 42754
rect 29250 42702 29262 42754
rect 29314 42702 29326 42754
rect 30482 42702 30494 42754
rect 30546 42702 30558 42754
rect 20078 42690 20130 42702
rect 22430 42690 22482 42702
rect 19742 42642 19794 42654
rect 17938 42590 17950 42642
rect 18002 42590 18014 42642
rect 19742 42578 19794 42590
rect 20750 42642 20802 42654
rect 26686 42642 26738 42654
rect 25554 42590 25566 42642
rect 25618 42590 25630 42642
rect 20750 42578 20802 42590
rect 26686 42578 26738 42590
rect 27918 42642 27970 42654
rect 27918 42578 27970 42590
rect 28478 42642 28530 42654
rect 33506 42590 33518 42642
rect 33570 42590 33582 42642
rect 28478 42578 28530 42590
rect 1710 42530 1762 42542
rect 1710 42466 1762 42478
rect 20414 42530 20466 42542
rect 20414 42466 20466 42478
rect 28142 42530 28194 42542
rect 28142 42466 28194 42478
rect 46174 42530 46226 42542
rect 46174 42466 46226 42478
rect 1344 42362 46592 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 46592 42362
rect 1344 42276 46592 42310
rect 33506 42030 33518 42082
rect 33570 42030 33582 42082
rect 19518 41970 19570 41982
rect 30046 41970 30098 41982
rect 12786 41918 12798 41970
rect 12850 41918 12862 41970
rect 14130 41918 14142 41970
rect 14194 41918 14206 41970
rect 20178 41918 20190 41970
rect 20242 41918 20254 41970
rect 22978 41918 22990 41970
rect 23042 41918 23054 41970
rect 23426 41918 23438 41970
rect 23490 41918 23502 41970
rect 25666 41918 25678 41970
rect 25730 41918 25742 41970
rect 26450 41918 26462 41970
rect 26514 41918 26526 41970
rect 19518 41906 19570 41918
rect 30046 41906 30098 41918
rect 30606 41970 30658 41982
rect 30606 41906 30658 41918
rect 30830 41970 30882 41982
rect 30830 41906 30882 41918
rect 31726 41970 31778 41982
rect 32498 41918 32510 41970
rect 32562 41918 32574 41970
rect 31726 41906 31778 41918
rect 18510 41858 18562 41870
rect 16034 41806 16046 41858
rect 16098 41806 16110 41858
rect 18510 41794 18562 41806
rect 28926 41858 28978 41870
rect 28926 41794 28978 41806
rect 24222 41746 24274 41758
rect 24222 41682 24274 41694
rect 1344 41578 46592 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 46592 41578
rect 1344 41492 46592 41526
rect 13694 41186 13746 41198
rect 14130 41134 14142 41186
rect 14194 41134 14206 41186
rect 14578 41134 14590 41186
rect 14642 41134 14654 41186
rect 23426 41134 23438 41186
rect 23490 41134 23502 41186
rect 24098 41134 24110 41186
rect 24162 41134 24174 41186
rect 26338 41134 26350 41186
rect 26402 41134 26414 41186
rect 26898 41134 26910 41186
rect 26962 41134 26974 41186
rect 29474 41134 29486 41186
rect 29538 41134 29550 41186
rect 29922 41134 29934 41186
rect 29986 41134 29998 41186
rect 31378 41134 31390 41186
rect 31442 41134 31454 41186
rect 32274 41134 32286 41186
rect 32338 41134 32350 41186
rect 13694 41122 13746 41134
rect 19294 41074 19346 41086
rect 19294 41010 19346 41022
rect 19630 41074 19682 41086
rect 19630 41010 19682 41022
rect 22878 41074 22930 41086
rect 22878 41010 22930 41022
rect 23214 41074 23266 41086
rect 23214 41010 23266 41022
rect 27582 41074 27634 41086
rect 27582 41010 27634 41022
rect 29150 41074 29202 41086
rect 29150 41010 29202 41022
rect 30606 41074 30658 41086
rect 30606 41010 30658 41022
rect 12574 40962 12626 40974
rect 13470 40962 13522 40974
rect 18062 40962 18114 40974
rect 12898 40910 12910 40962
rect 12962 40910 12974 40962
rect 17378 40910 17390 40962
rect 17442 40910 17454 40962
rect 12574 40898 12626 40910
rect 13470 40898 13522 40910
rect 18062 40898 18114 40910
rect 19070 40962 19122 40974
rect 28254 40962 28306 40974
rect 27906 40910 27918 40962
rect 27970 40910 27982 40962
rect 30146 40910 30158 40962
rect 30210 40910 30222 40962
rect 19070 40898 19122 40910
rect 28254 40898 28306 40910
rect 1344 40794 46592 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 46592 40794
rect 1344 40708 46592 40742
rect 24110 40626 24162 40638
rect 24110 40562 24162 40574
rect 11454 40514 11506 40526
rect 11454 40450 11506 40462
rect 12126 40514 12178 40526
rect 15934 40514 15986 40526
rect 12562 40462 12574 40514
rect 12626 40462 12638 40514
rect 12126 40450 12178 40462
rect 15934 40450 15986 40462
rect 26798 40514 26850 40526
rect 30382 40514 30434 40526
rect 27794 40462 27806 40514
rect 27858 40462 27870 40514
rect 37874 40462 37886 40514
rect 37938 40462 37950 40514
rect 26798 40450 26850 40462
rect 30382 40450 30434 40462
rect 16270 40402 16322 40414
rect 28478 40402 28530 40414
rect 31278 40402 31330 40414
rect 11218 40350 11230 40402
rect 11282 40350 11294 40402
rect 11890 40350 11902 40402
rect 11954 40350 11966 40402
rect 14242 40350 14254 40402
rect 14306 40350 14318 40402
rect 15138 40350 15150 40402
rect 15202 40350 15214 40402
rect 17378 40350 17390 40402
rect 17442 40350 17454 40402
rect 19394 40350 19406 40402
rect 19458 40350 19470 40402
rect 19842 40350 19854 40402
rect 19906 40350 19918 40402
rect 22082 40350 22094 40402
rect 22146 40350 22158 40402
rect 23874 40350 23886 40402
rect 23938 40350 23950 40402
rect 27122 40350 27134 40402
rect 27186 40350 27198 40402
rect 27570 40350 27582 40402
rect 27634 40350 27646 40402
rect 28914 40350 28926 40402
rect 28978 40350 28990 40402
rect 29922 40350 29934 40402
rect 29986 40350 29998 40402
rect 30818 40350 30830 40402
rect 30882 40350 30894 40402
rect 16270 40338 16322 40350
rect 28478 40338 28530 40350
rect 31278 40338 31330 40350
rect 31838 40402 31890 40414
rect 35074 40350 35086 40402
rect 35138 40350 35150 40402
rect 35522 40350 35534 40402
rect 35586 40350 35598 40402
rect 31838 40338 31890 40350
rect 13906 40238 13918 40290
rect 13970 40238 13982 40290
rect 18274 40238 18286 40290
rect 18338 40238 18350 40290
rect 15486 40178 15538 40190
rect 38670 40178 38722 40190
rect 23090 40126 23102 40178
rect 23154 40126 23166 40178
rect 15486 40114 15538 40126
rect 38670 40114 38722 40126
rect 1344 40010 46592 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 46592 40010
rect 1344 39924 46592 39958
rect 34190 39842 34242 39854
rect 34190 39778 34242 39790
rect 22094 39730 22146 39742
rect 13682 39678 13694 39730
rect 13746 39678 13758 39730
rect 22094 39666 22146 39678
rect 22430 39730 22482 39742
rect 37650 39678 37662 39730
rect 37714 39678 37726 39730
rect 22430 39666 22482 39678
rect 15038 39618 15090 39630
rect 21310 39618 21362 39630
rect 24110 39618 24162 39630
rect 14354 39566 14366 39618
rect 14418 39566 14430 39618
rect 15586 39566 15598 39618
rect 15650 39566 15662 39618
rect 16146 39566 16158 39618
rect 16210 39566 16222 39618
rect 19394 39566 19406 39618
rect 19458 39566 19470 39618
rect 22754 39566 22766 39618
rect 22818 39566 22830 39618
rect 23202 39566 23214 39618
rect 23266 39566 23278 39618
rect 24434 39566 24446 39618
rect 24498 39566 24510 39618
rect 25554 39566 25566 39618
rect 25618 39566 25630 39618
rect 28018 39566 28030 39618
rect 28082 39566 28094 39618
rect 29810 39566 29822 39618
rect 29874 39566 29886 39618
rect 30034 39566 30046 39618
rect 30098 39566 30110 39618
rect 33618 39566 33630 39618
rect 33682 39566 33694 39618
rect 15038 39554 15090 39566
rect 21310 39554 21362 39566
rect 24110 39554 24162 39566
rect 19070 39506 19122 39518
rect 27694 39506 27746 39518
rect 9202 39454 9214 39506
rect 9266 39454 9278 39506
rect 21634 39454 21646 39506
rect 21698 39454 21710 39506
rect 19070 39442 19122 39454
rect 27694 39442 27746 39454
rect 28254 39506 28306 39518
rect 28254 39442 28306 39454
rect 29374 39506 29426 39518
rect 29374 39442 29426 39454
rect 33182 39506 33234 39518
rect 37886 39506 37938 39518
rect 37314 39454 37326 39506
rect 37378 39454 37390 39506
rect 33182 39442 33234 39454
rect 37886 39442 37938 39454
rect 38670 39506 38722 39518
rect 38670 39442 38722 39454
rect 39454 39506 39506 39518
rect 39454 39442 39506 39454
rect 14814 39394 14866 39406
rect 12786 39342 12798 39394
rect 12850 39342 12862 39394
rect 14814 39330 14866 39342
rect 15262 39394 15314 39406
rect 15262 39330 15314 39342
rect 20526 39394 20578 39406
rect 29150 39394 29202 39406
rect 23426 39342 23438 39394
rect 23490 39342 23502 39394
rect 20526 39330 20578 39342
rect 29150 39330 29202 39342
rect 34750 39394 34802 39406
rect 34750 39330 34802 39342
rect 1344 39226 46592 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 46592 39226
rect 1344 39140 46592 39174
rect 21758 39058 21810 39070
rect 39454 39058 39506 39070
rect 4834 39006 4846 39058
rect 4898 39006 4910 39058
rect 29362 39006 29374 39058
rect 29426 39006 29438 39058
rect 21758 38994 21810 39006
rect 39454 38994 39506 39006
rect 16718 38946 16770 38958
rect 20974 38946 21026 38958
rect 11666 38894 11678 38946
rect 11730 38894 11742 38946
rect 18386 38894 18398 38946
rect 18450 38894 18462 38946
rect 16718 38882 16770 38894
rect 20974 38882 21026 38894
rect 21310 38946 21362 38958
rect 32510 38946 32562 38958
rect 22418 38894 22430 38946
rect 22482 38894 22494 38946
rect 23986 38894 23998 38946
rect 24050 38894 24062 38946
rect 27570 38894 27582 38946
rect 27634 38894 27646 38946
rect 21310 38882 21362 38894
rect 32510 38882 32562 38894
rect 1934 38834 1986 38846
rect 16270 38834 16322 38846
rect 19070 38834 19122 38846
rect 23214 38834 23266 38846
rect 38558 38834 38610 38846
rect 2370 38782 2382 38834
rect 2434 38782 2446 38834
rect 14354 38782 14366 38834
rect 14418 38782 14430 38834
rect 15250 38782 15262 38834
rect 15314 38782 15326 38834
rect 17714 38782 17726 38834
rect 17778 38782 17790 38834
rect 18274 38782 18286 38834
rect 18338 38782 18350 38834
rect 19618 38782 19630 38834
rect 19682 38782 19694 38834
rect 20514 38782 20526 38834
rect 20578 38782 20590 38834
rect 22194 38782 22206 38834
rect 22258 38782 22270 38834
rect 23762 38782 23774 38834
rect 23826 38782 23838 38834
rect 32274 38782 32286 38834
rect 32338 38782 32350 38834
rect 33058 38782 33070 38834
rect 33122 38782 33134 38834
rect 33506 38782 33518 38834
rect 33570 38782 33582 38834
rect 35858 38782 35870 38834
rect 35922 38782 35934 38834
rect 36306 38782 36318 38834
rect 36370 38782 36382 38834
rect 37762 38782 37774 38834
rect 37826 38782 37838 38834
rect 1934 38770 1986 38782
rect 16270 38770 16322 38782
rect 19070 38770 19122 38782
rect 23214 38770 23266 38782
rect 38558 38770 38610 38782
rect 39118 38834 39170 38846
rect 41582 38834 41634 38846
rect 39666 38782 39678 38834
rect 39730 38782 39742 38834
rect 39118 38770 39170 38782
rect 41582 38770 41634 38782
rect 41806 38834 41858 38846
rect 41806 38770 41858 38782
rect 17390 38722 17442 38734
rect 13794 38670 13806 38722
rect 13858 38670 13870 38722
rect 17390 38658 17442 38670
rect 24558 38722 24610 38734
rect 24558 38658 24610 38670
rect 38222 38722 38274 38734
rect 38222 38658 38274 38670
rect 41134 38722 41186 38734
rect 41134 38658 41186 38670
rect 41358 38722 41410 38734
rect 41682 38670 41694 38722
rect 41746 38670 41758 38722
rect 41358 38658 41410 38670
rect 5406 38610 5458 38622
rect 5406 38546 5458 38558
rect 22878 38610 22930 38622
rect 40910 38610 40962 38622
rect 37202 38558 37214 38610
rect 37266 38558 37278 38610
rect 22878 38546 22930 38558
rect 40910 38546 40962 38558
rect 1344 38442 46592 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 46592 38442
rect 1344 38356 46592 38390
rect 14814 38162 14866 38174
rect 14814 38098 14866 38110
rect 20190 38162 20242 38174
rect 22082 38110 22094 38162
rect 22146 38110 22158 38162
rect 43138 38110 43150 38162
rect 43202 38110 43214 38162
rect 20190 38098 20242 38110
rect 16494 38050 16546 38062
rect 19182 38050 19234 38062
rect 22542 38050 22594 38062
rect 13682 37998 13694 38050
rect 13746 37998 13758 38050
rect 15138 37998 15150 38050
rect 15202 37998 15214 38050
rect 15586 37998 15598 38050
rect 15650 37998 15662 38050
rect 16818 37998 16830 38050
rect 16882 37998 16894 38050
rect 17938 37998 17950 38050
rect 18002 37998 18014 38050
rect 20626 37998 20638 38050
rect 20690 37998 20702 38050
rect 16494 37986 16546 37998
rect 19182 37986 19234 37998
rect 22542 37986 22594 37998
rect 22990 38050 23042 38062
rect 23426 37998 23438 38050
rect 23490 37998 23502 38050
rect 31714 37998 31726 38050
rect 31778 37998 31790 38050
rect 32498 37998 32510 38050
rect 32562 37998 32574 38050
rect 37314 37998 37326 38050
rect 37378 37998 37390 38050
rect 37762 37998 37774 38050
rect 37826 37998 37838 38050
rect 38994 37998 39006 38050
rect 39058 37998 39070 38050
rect 40002 37998 40014 38050
rect 40066 37998 40078 38050
rect 40898 37998 40910 38050
rect 40962 37998 40974 38050
rect 42466 37998 42478 38050
rect 42530 37998 42542 38050
rect 42690 37998 42702 38050
rect 42754 37998 42766 38050
rect 22990 37986 23042 37998
rect 13470 37938 13522 37950
rect 13470 37874 13522 37886
rect 18846 37938 18898 37950
rect 18846 37874 18898 37886
rect 21310 37938 21362 37950
rect 21310 37874 21362 37886
rect 23886 37938 23938 37950
rect 36990 37938 37042 37950
rect 34626 37886 34638 37938
rect 34690 37886 34702 37938
rect 36082 37886 36094 37938
rect 36146 37886 36158 37938
rect 23886 37874 23938 37886
rect 36990 37874 37042 37886
rect 38446 37938 38498 37950
rect 43698 37886 43710 37938
rect 43762 37886 43774 37938
rect 38446 37874 38498 37886
rect 19854 37826 19906 37838
rect 15810 37774 15822 37826
rect 15874 37774 15886 37826
rect 19506 37774 19518 37826
rect 19570 37774 19582 37826
rect 19854 37762 19906 37774
rect 21646 37826 21698 37838
rect 24558 37826 24610 37838
rect 24210 37774 24222 37826
rect 24274 37774 24286 37826
rect 21646 37762 21698 37774
rect 24558 37762 24610 37774
rect 24894 37826 24946 37838
rect 25218 37774 25230 37826
rect 25282 37774 25294 37826
rect 37986 37774 37998 37826
rect 38050 37774 38062 37826
rect 24894 37762 24946 37774
rect 1344 37658 46592 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 46592 37658
rect 1344 37572 46592 37606
rect 14702 37490 14754 37502
rect 25790 37490 25842 37502
rect 5394 37438 5406 37490
rect 5458 37438 5470 37490
rect 13458 37438 13470 37490
rect 13522 37438 13534 37490
rect 22530 37438 22542 37490
rect 22594 37438 22606 37490
rect 14702 37426 14754 37438
rect 25790 37426 25842 37438
rect 29710 37490 29762 37502
rect 29710 37426 29762 37438
rect 30046 37490 30098 37502
rect 30046 37426 30098 37438
rect 38558 37490 38610 37502
rect 38558 37426 38610 37438
rect 41694 37490 41746 37502
rect 41694 37426 41746 37438
rect 16046 37378 16098 37390
rect 21310 37378 21362 37390
rect 28366 37378 28418 37390
rect 18946 37326 18958 37378
rect 19010 37326 19022 37378
rect 19730 37326 19742 37378
rect 19794 37326 19806 37378
rect 24434 37326 24446 37378
rect 24498 37326 24510 37378
rect 16046 37314 16098 37326
rect 21310 37314 21362 37326
rect 28366 37314 28418 37326
rect 32398 37378 32450 37390
rect 32398 37314 32450 37326
rect 34638 37378 34690 37390
rect 40910 37378 40962 37390
rect 40338 37326 40350 37378
rect 40402 37326 40414 37378
rect 34638 37314 34690 37326
rect 40910 37314 40962 37326
rect 2718 37266 2770 37278
rect 10782 37266 10834 37278
rect 15038 37266 15090 37278
rect 3154 37214 3166 37266
rect 3218 37214 3230 37266
rect 11218 37214 11230 37266
rect 11282 37214 11294 37266
rect 2718 37202 2770 37214
rect 10782 37202 10834 37214
rect 15038 37202 15090 37214
rect 15710 37266 15762 37278
rect 22878 37266 22930 37278
rect 26462 37266 26514 37278
rect 17826 37214 17838 37266
rect 17890 37214 17902 37266
rect 18722 37214 18734 37266
rect 18786 37214 18798 37266
rect 23426 37214 23438 37266
rect 23490 37214 23502 37266
rect 23986 37214 23998 37266
rect 24050 37214 24062 37266
rect 24546 37214 24558 37266
rect 24610 37214 24622 37266
rect 26114 37214 26126 37266
rect 26178 37214 26190 37266
rect 15710 37202 15762 37214
rect 22878 37202 22930 37214
rect 26462 37202 26514 37214
rect 28702 37266 28754 37278
rect 28702 37202 28754 37214
rect 30382 37266 30434 37278
rect 35870 37266 35922 37278
rect 37662 37266 37714 37278
rect 31266 37214 31278 37266
rect 31330 37214 31342 37266
rect 32162 37214 32174 37266
rect 32226 37214 32238 37266
rect 34402 37214 34414 37266
rect 34466 37214 34478 37266
rect 35410 37214 35422 37266
rect 35474 37214 35486 37266
rect 36642 37214 36654 37266
rect 36706 37214 36718 37266
rect 38882 37214 38894 37266
rect 38946 37214 38958 37266
rect 40002 37214 40014 37266
rect 40066 37214 40078 37266
rect 41234 37214 41246 37266
rect 41298 37214 41310 37266
rect 43138 37214 43150 37266
rect 43202 37214 43214 37266
rect 44146 37214 44158 37266
rect 44210 37214 44222 37266
rect 30382 37202 30434 37214
rect 35870 37202 35922 37214
rect 37662 37202 37714 37214
rect 16494 37154 16546 37166
rect 14354 37102 14366 37154
rect 14418 37102 14430 37154
rect 16494 37090 16546 37102
rect 17390 37154 17442 37166
rect 33966 37154 34018 37166
rect 42030 37154 42082 37166
rect 19506 37102 19518 37154
rect 19570 37102 19582 37154
rect 21970 37102 21982 37154
rect 22034 37102 22046 37154
rect 25330 37102 25342 37154
rect 25394 37102 25406 37154
rect 29250 37102 29262 37154
rect 29314 37102 29326 37154
rect 31602 37102 31614 37154
rect 31666 37102 31678 37154
rect 35746 37102 35758 37154
rect 35810 37102 35822 37154
rect 37426 37102 37438 37154
rect 37490 37102 37502 37154
rect 38098 37102 38110 37154
rect 38162 37102 38174 37154
rect 39554 37102 39566 37154
rect 39618 37102 39630 37154
rect 17390 37090 17442 37102
rect 33966 37090 34018 37102
rect 42030 37090 42082 37102
rect 6190 37042 6242 37054
rect 26126 37042 26178 37054
rect 42814 37042 42866 37054
rect 24322 36990 24334 37042
rect 24386 36990 24398 37042
rect 36530 36990 36542 37042
rect 36594 36990 36606 37042
rect 6190 36978 6242 36990
rect 26126 36978 26178 36990
rect 42814 36978 42866 36990
rect 1344 36874 46592 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 46592 36874
rect 1344 36788 46592 36822
rect 22318 36706 22370 36718
rect 35410 36654 35422 36706
rect 35474 36654 35486 36706
rect 22318 36642 22370 36654
rect 13694 36594 13746 36606
rect 17838 36594 17890 36606
rect 43374 36594 43426 36606
rect 12898 36542 12910 36594
rect 12962 36542 12974 36594
rect 15474 36542 15486 36594
rect 15538 36542 15550 36594
rect 19618 36542 19630 36594
rect 19682 36542 19694 36594
rect 28130 36542 28142 36594
rect 28194 36542 28206 36594
rect 35970 36542 35982 36594
rect 36034 36542 36046 36594
rect 37090 36542 37102 36594
rect 37154 36542 37166 36594
rect 13694 36530 13746 36542
rect 17838 36530 17890 36542
rect 43374 36530 43426 36542
rect 14254 36482 14306 36494
rect 21646 36482 21698 36494
rect 9426 36430 9438 36482
rect 9490 36430 9502 36482
rect 10098 36430 10110 36482
rect 10162 36430 10174 36482
rect 19506 36430 19518 36482
rect 19570 36430 19582 36482
rect 14254 36418 14306 36430
rect 21646 36418 21698 36430
rect 21870 36482 21922 36494
rect 21870 36418 21922 36430
rect 22094 36482 22146 36494
rect 22094 36418 22146 36430
rect 25118 36482 25170 36494
rect 30606 36482 30658 36494
rect 39790 36482 39842 36494
rect 25442 36430 25454 36482
rect 25506 36430 25518 36482
rect 29474 36430 29486 36482
rect 29538 36430 29550 36482
rect 29922 36430 29934 36482
rect 29986 36430 29998 36482
rect 31378 36430 31390 36482
rect 31442 36430 31454 36482
rect 32274 36430 32286 36482
rect 32338 36430 32350 36482
rect 32946 36430 32958 36482
rect 33010 36430 33022 36482
rect 34290 36430 34302 36482
rect 34354 36430 34366 36482
rect 36194 36430 36206 36482
rect 36258 36430 36270 36482
rect 38546 36430 38558 36482
rect 38610 36430 38622 36482
rect 39442 36430 39454 36482
rect 39506 36430 39518 36482
rect 25118 36418 25170 36430
rect 30606 36418 30658 36430
rect 39790 36418 39842 36430
rect 43038 36482 43090 36494
rect 43038 36418 43090 36430
rect 43262 36482 43314 36494
rect 43262 36418 43314 36430
rect 43486 36482 43538 36494
rect 43486 36418 43538 36430
rect 6302 36370 6354 36382
rect 6302 36306 6354 36318
rect 6638 36370 6690 36382
rect 6638 36306 6690 36318
rect 7086 36370 7138 36382
rect 7086 36306 7138 36318
rect 9662 36370 9714 36382
rect 16494 36370 16546 36382
rect 10770 36318 10782 36370
rect 10834 36318 10846 36370
rect 15250 36318 15262 36370
rect 15314 36318 15326 36370
rect 9662 36306 9714 36318
rect 16494 36306 16546 36318
rect 19630 36370 19682 36382
rect 26574 36370 26626 36382
rect 20738 36318 20750 36370
rect 20802 36318 20814 36370
rect 23538 36318 23550 36370
rect 23602 36318 23614 36370
rect 19630 36306 19682 36318
rect 26574 36306 26626 36318
rect 29150 36370 29202 36382
rect 39230 36370 39282 36382
rect 38098 36318 38110 36370
rect 38162 36318 38174 36370
rect 29150 36306 29202 36318
rect 39230 36306 39282 36318
rect 40686 36370 40738 36382
rect 40686 36306 40738 36318
rect 41022 36370 41074 36382
rect 41022 36306 41074 36318
rect 5182 36258 5234 36270
rect 5966 36258 6018 36270
rect 5618 36206 5630 36258
rect 5682 36206 5694 36258
rect 5182 36194 5234 36206
rect 5966 36194 6018 36206
rect 6974 36258 7026 36270
rect 22766 36258 22818 36270
rect 27806 36258 27858 36270
rect 15362 36206 15374 36258
rect 15426 36206 15438 36258
rect 24882 36206 24894 36258
rect 24946 36206 24958 36258
rect 6974 36194 7026 36206
rect 22766 36194 22818 36206
rect 27806 36194 27858 36206
rect 28590 36258 28642 36270
rect 37550 36258 37602 36270
rect 40126 36258 40178 36270
rect 30146 36206 30158 36258
rect 30210 36206 30222 36258
rect 38546 36206 38558 36258
rect 38610 36206 38622 36258
rect 28590 36194 28642 36206
rect 37550 36194 37602 36206
rect 40126 36194 40178 36206
rect 1344 36090 46592 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 46592 36090
rect 1344 36004 46592 36038
rect 7534 35922 7586 35934
rect 6738 35870 6750 35922
rect 6802 35870 6814 35922
rect 7534 35858 7586 35870
rect 10110 35922 10162 35934
rect 10110 35858 10162 35870
rect 15486 35922 15538 35934
rect 19966 35922 20018 35934
rect 16482 35870 16494 35922
rect 16546 35870 16558 35922
rect 19618 35870 19630 35922
rect 19682 35870 19694 35922
rect 15486 35858 15538 35870
rect 19966 35858 20018 35870
rect 27358 35922 27410 35934
rect 39118 35922 39170 35934
rect 31826 35870 31838 35922
rect 31890 35870 31902 35922
rect 27358 35858 27410 35870
rect 39118 35858 39170 35870
rect 39902 35922 39954 35934
rect 43026 35870 43038 35922
rect 43090 35870 43102 35922
rect 39902 35858 39954 35870
rect 15822 35810 15874 35822
rect 21198 35810 21250 35822
rect 35534 35810 35586 35822
rect 41134 35810 41186 35822
rect 17602 35758 17614 35810
rect 17666 35758 17678 35810
rect 22194 35758 22206 35810
rect 22258 35758 22270 35810
rect 26674 35758 26686 35810
rect 26738 35758 26750 35810
rect 30930 35758 30942 35810
rect 30994 35758 31006 35810
rect 36530 35758 36542 35810
rect 36594 35758 36606 35810
rect 15822 35746 15874 35758
rect 21198 35746 21250 35758
rect 35534 35746 35586 35758
rect 41134 35746 41186 35758
rect 41470 35810 41522 35822
rect 41470 35746 41522 35758
rect 44830 35810 44882 35822
rect 44830 35746 44882 35758
rect 3838 35698 3890 35710
rect 20862 35698 20914 35710
rect 22878 35698 22930 35710
rect 25902 35698 25954 35710
rect 27134 35698 27186 35710
rect 34190 35698 34242 35710
rect 4498 35646 4510 35698
rect 4562 35646 4574 35698
rect 10658 35646 10670 35698
rect 10722 35646 10734 35698
rect 12898 35646 12910 35698
rect 12962 35646 12974 35698
rect 13458 35646 13470 35698
rect 13522 35646 13534 35698
rect 16706 35646 16718 35698
rect 16770 35646 16782 35698
rect 17490 35646 17502 35698
rect 17554 35646 17566 35698
rect 21522 35646 21534 35698
rect 21586 35646 21598 35698
rect 21970 35646 21982 35698
rect 22034 35646 22046 35698
rect 23314 35646 23326 35698
rect 23378 35646 23390 35698
rect 24322 35646 24334 35698
rect 24386 35646 24398 35698
rect 26338 35646 26350 35698
rect 26402 35646 26414 35698
rect 27682 35646 27694 35698
rect 27746 35646 27758 35698
rect 28242 35646 28254 35698
rect 28306 35646 28318 35698
rect 3838 35634 3890 35646
rect 20862 35634 20914 35646
rect 22878 35634 22930 35646
rect 25902 35634 25954 35646
rect 27134 35634 27186 35646
rect 34190 35634 34242 35646
rect 34750 35698 34802 35710
rect 37214 35698 37266 35710
rect 42702 35698 42754 35710
rect 35970 35646 35982 35698
rect 36034 35646 36046 35698
rect 36418 35646 36430 35698
rect 36482 35646 36494 35698
rect 37762 35646 37774 35698
rect 37826 35646 37838 35698
rect 38546 35646 38558 35698
rect 38610 35646 38622 35698
rect 39330 35646 39342 35698
rect 39394 35646 39406 35698
rect 43474 35646 43486 35698
rect 43538 35646 43550 35698
rect 34750 35634 34802 35646
rect 37214 35634 37266 35646
rect 42702 35634 42754 35646
rect 3614 35586 3666 35598
rect 3614 35522 3666 35534
rect 7870 35586 7922 35598
rect 7870 35522 7922 35534
rect 19182 35586 19234 35598
rect 42366 35586 42418 35598
rect 20402 35534 20414 35586
rect 20466 35534 20478 35586
rect 19182 35522 19234 35534
rect 42366 35522 42418 35534
rect 44718 35586 44770 35598
rect 44718 35522 44770 35534
rect 7758 35474 7810 35486
rect 7758 35410 7810 35422
rect 14590 35474 14642 35486
rect 14590 35410 14642 35422
rect 18286 35474 18338 35486
rect 18286 35410 18338 35422
rect 18622 35474 18674 35486
rect 18622 35410 18674 35422
rect 25566 35474 25618 35486
rect 25566 35410 25618 35422
rect 1344 35306 46592 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 46592 35306
rect 1344 35220 46592 35254
rect 2942 35138 2994 35150
rect 2942 35074 2994 35086
rect 9214 35138 9266 35150
rect 33182 35138 33234 35150
rect 28466 35086 28478 35138
rect 28530 35086 28542 35138
rect 9214 35074 9266 35086
rect 33182 35074 33234 35086
rect 3054 35026 3106 35038
rect 3054 34962 3106 34974
rect 22878 35026 22930 35038
rect 22878 34962 22930 34974
rect 26574 35026 26626 35038
rect 26574 34962 26626 34974
rect 27134 35026 27186 35038
rect 27134 34962 27186 34974
rect 37998 35026 38050 35038
rect 37998 34962 38050 34974
rect 38222 35026 38274 35038
rect 38222 34962 38274 34974
rect 41470 35026 41522 35038
rect 41470 34962 41522 34974
rect 5518 34914 5570 34926
rect 14590 34914 14642 34926
rect 24334 34914 24386 34926
rect 29150 34914 29202 34926
rect 3490 34862 3502 34914
rect 3554 34862 3566 34914
rect 6178 34862 6190 34914
rect 6242 34862 6254 34914
rect 14914 34862 14926 34914
rect 14978 34862 14990 34914
rect 15362 34862 15374 34914
rect 15426 34862 15438 34914
rect 16594 34862 16606 34914
rect 16658 34862 16670 34914
rect 17714 34862 17726 34914
rect 17778 34862 17790 34914
rect 23202 34862 23214 34914
rect 23266 34862 23278 34914
rect 23762 34862 23774 34914
rect 23826 34862 23838 34914
rect 24882 34862 24894 34914
rect 24946 34862 24958 34914
rect 26002 34862 26014 34914
rect 26066 34862 26078 34914
rect 5518 34850 5570 34862
rect 14590 34850 14642 34862
rect 24334 34850 24386 34862
rect 29150 34850 29202 34862
rect 29374 34914 29426 34926
rect 39118 34914 39170 34926
rect 29698 34862 29710 34914
rect 29762 34862 29774 34914
rect 30146 34862 30158 34914
rect 30210 34862 30222 34914
rect 37426 34862 37438 34914
rect 37490 34862 37502 34914
rect 38658 34862 38670 34914
rect 38722 34862 38734 34914
rect 29374 34850 29426 34862
rect 39118 34850 39170 34862
rect 39454 34914 39506 34926
rect 39454 34850 39506 34862
rect 40126 34914 40178 34926
rect 41010 34862 41022 34914
rect 41074 34862 41086 34914
rect 41906 34862 41918 34914
rect 41970 34862 41982 34914
rect 42690 34862 42702 34914
rect 42754 34862 42766 34914
rect 40126 34850 40178 34862
rect 1710 34802 1762 34814
rect 1710 34738 1762 34750
rect 2046 34802 2098 34814
rect 11118 34802 11170 34814
rect 4722 34750 4734 34802
rect 4786 34750 4798 34802
rect 2046 34738 2098 34750
rect 11118 34738 11170 34750
rect 11454 34802 11506 34814
rect 16046 34802 16098 34814
rect 15586 34750 15598 34802
rect 15650 34750 15662 34802
rect 11454 34738 11506 34750
rect 16046 34738 16098 34750
rect 22542 34802 22594 34814
rect 37662 34802 37714 34814
rect 27570 34750 27582 34802
rect 27634 34750 27646 34802
rect 22542 34738 22594 34750
rect 37662 34738 37714 34750
rect 39790 34802 39842 34814
rect 39790 34738 39842 34750
rect 40462 34802 40514 34814
rect 45166 34802 45218 34814
rect 43922 34750 43934 34802
rect 43986 34750 43998 34802
rect 40462 34738 40514 34750
rect 45166 34738 45218 34750
rect 2494 34690 2546 34702
rect 2494 34626 2546 34638
rect 3726 34690 3778 34702
rect 3726 34626 3778 34638
rect 4062 34690 4114 34702
rect 5070 34690 5122 34702
rect 21982 34690 22034 34702
rect 37102 34690 37154 34702
rect 4386 34638 4398 34690
rect 4450 34638 4462 34690
rect 8418 34638 8430 34690
rect 8482 34638 8494 34690
rect 23874 34638 23886 34690
rect 23938 34638 23950 34690
rect 4062 34626 4114 34638
rect 5070 34626 5122 34638
rect 21982 34626 22034 34638
rect 37102 34626 37154 34638
rect 37214 34690 37266 34702
rect 37214 34626 37266 34638
rect 37774 34690 37826 34702
rect 37774 34626 37826 34638
rect 44830 34690 44882 34702
rect 44830 34626 44882 34638
rect 1344 34522 46592 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 46592 34522
rect 1344 34436 46592 34470
rect 23326 34354 23378 34366
rect 4722 34302 4734 34354
rect 4786 34302 4798 34354
rect 8306 34302 8318 34354
rect 8370 34302 8382 34354
rect 23326 34290 23378 34302
rect 23886 34354 23938 34366
rect 29934 34354 29986 34366
rect 25554 34302 25566 34354
rect 25618 34302 25630 34354
rect 23886 34290 23938 34302
rect 29934 34290 29986 34302
rect 39454 34354 39506 34366
rect 39454 34290 39506 34302
rect 41134 34354 41186 34366
rect 41134 34290 41186 34302
rect 13694 34242 13746 34254
rect 13694 34178 13746 34190
rect 15598 34242 15650 34254
rect 16158 34242 16210 34254
rect 15810 34190 15822 34242
rect 15874 34190 15886 34242
rect 15598 34178 15650 34190
rect 16158 34178 16210 34190
rect 16830 34242 16882 34254
rect 22430 34242 22482 34254
rect 17826 34190 17838 34242
rect 17890 34190 17902 34242
rect 18162 34190 18174 34242
rect 18226 34190 18238 34242
rect 22082 34190 22094 34242
rect 22146 34190 22158 34242
rect 16830 34178 16882 34190
rect 22430 34178 22482 34190
rect 25230 34242 25282 34254
rect 37662 34242 37714 34254
rect 26450 34190 26462 34242
rect 26514 34190 26526 34242
rect 25230 34178 25282 34190
rect 37662 34178 37714 34190
rect 38334 34242 38386 34254
rect 38334 34178 38386 34190
rect 44942 34242 44994 34254
rect 44942 34178 44994 34190
rect 1822 34130 1874 34142
rect 5630 34130 5682 34142
rect 9102 34130 9154 34142
rect 2146 34078 2158 34130
rect 2210 34078 2222 34130
rect 6066 34078 6078 34130
rect 6130 34078 6142 34130
rect 1822 34066 1874 34078
rect 5630 34066 5682 34078
rect 9102 34066 9154 34078
rect 9662 34130 9714 34142
rect 9662 34066 9714 34078
rect 10782 34130 10834 34142
rect 16494 34130 16546 34142
rect 11330 34078 11342 34130
rect 11394 34078 11406 34130
rect 10782 34066 10834 34078
rect 16494 34066 16546 34078
rect 23214 34130 23266 34142
rect 23214 34066 23266 34078
rect 23438 34130 23490 34142
rect 37998 34130 38050 34142
rect 37426 34078 37438 34130
rect 37490 34078 37502 34130
rect 23438 34066 23490 34078
rect 37998 34066 38050 34078
rect 39790 34130 39842 34142
rect 40910 34130 40962 34142
rect 40226 34078 40238 34130
rect 40290 34078 40302 34130
rect 41458 34078 41470 34130
rect 41522 34078 41534 34130
rect 41794 34078 41806 34130
rect 41858 34078 41870 34130
rect 45378 34078 45390 34130
rect 45442 34078 45454 34130
rect 39790 34066 39842 34078
rect 40910 34066 40962 34078
rect 19294 34018 19346 34030
rect 19294 33954 19346 33966
rect 24446 34018 24498 34030
rect 24446 33954 24498 33966
rect 36990 34018 37042 34030
rect 36990 33954 37042 33966
rect 38894 34018 38946 34030
rect 38894 33954 38946 33966
rect 5294 33906 5346 33918
rect 5294 33842 5346 33854
rect 9550 33906 9602 33918
rect 9550 33842 9602 33854
rect 14478 33906 14530 33918
rect 14478 33842 14530 33854
rect 18398 33906 18450 33918
rect 18398 33842 18450 33854
rect 18734 33906 18786 33918
rect 18734 33842 18786 33854
rect 22878 33906 22930 33918
rect 22878 33842 22930 33854
rect 22990 33906 23042 33918
rect 45938 33854 45950 33906
rect 46002 33854 46014 33906
rect 22990 33842 23042 33854
rect 1344 33738 46592 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 46592 33738
rect 1344 33652 46592 33686
rect 4174 33570 4226 33582
rect 4174 33506 4226 33518
rect 4286 33458 4338 33470
rect 4286 33394 4338 33406
rect 4958 33458 5010 33470
rect 29262 33458 29314 33470
rect 24658 33406 24670 33458
rect 24722 33406 24734 33458
rect 4958 33394 5010 33406
rect 29262 33394 29314 33406
rect 5630 33346 5682 33358
rect 6638 33346 6690 33358
rect 21310 33346 21362 33358
rect 22430 33346 22482 33358
rect 29038 33346 29090 33358
rect 6066 33294 6078 33346
rect 6130 33294 6142 33346
rect 6962 33294 6974 33346
rect 7026 33294 7038 33346
rect 10546 33294 10558 33346
rect 10610 33294 10622 33346
rect 13458 33294 13470 33346
rect 13522 33294 13534 33346
rect 13906 33294 13918 33346
rect 13970 33294 13982 33346
rect 16930 33294 16942 33346
rect 16994 33294 17006 33346
rect 17266 33294 17278 33346
rect 17330 33294 17342 33346
rect 21746 33294 21758 33346
rect 21810 33294 21822 33346
rect 25218 33294 25230 33346
rect 25282 33294 25294 33346
rect 5630 33282 5682 33294
rect 6638 33282 6690 33294
rect 21310 33282 21362 33294
rect 22430 33282 22482 33294
rect 29038 33282 29090 33294
rect 32062 33346 32114 33358
rect 42702 33346 42754 33358
rect 32386 33294 32398 33346
rect 32450 33294 32462 33346
rect 41346 33294 41358 33346
rect 41410 33294 41422 33346
rect 41794 33294 41806 33346
rect 41858 33294 41870 33346
rect 43250 33294 43262 33346
rect 43314 33294 43326 33346
rect 44146 33294 44158 33346
rect 44210 33294 44222 33346
rect 32062 33282 32114 33294
rect 42702 33282 42754 33294
rect 3726 33234 3778 33246
rect 3726 33170 3778 33182
rect 3838 33234 3890 33246
rect 3838 33170 3890 33182
rect 10334 33234 10386 33246
rect 10334 33170 10386 33182
rect 22206 33234 22258 33246
rect 22206 33170 22258 33182
rect 28254 33234 28306 33246
rect 28254 33170 28306 33182
rect 29598 33234 29650 33246
rect 29598 33170 29650 33182
rect 37102 33234 37154 33246
rect 40798 33234 40850 33246
rect 38322 33182 38334 33234
rect 38386 33182 38398 33234
rect 37102 33170 37154 33182
rect 40798 33170 40850 33182
rect 41022 33234 41074 33246
rect 41022 33170 41074 33182
rect 4846 33122 4898 33134
rect 10110 33122 10162 33134
rect 22766 33122 22818 33134
rect 9538 33070 9550 33122
rect 9602 33070 9614 33122
rect 18050 33070 18062 33122
rect 18114 33070 18126 33122
rect 4846 33058 4898 33070
rect 10110 33058 10162 33070
rect 22766 33058 22818 33070
rect 24222 33122 24274 33134
rect 28702 33122 28754 33134
rect 25442 33070 25454 33122
rect 25506 33070 25518 33122
rect 24222 33058 24274 33070
rect 28702 33058 28754 33070
rect 29374 33122 29426 33134
rect 35534 33122 35586 33134
rect 34738 33070 34750 33122
rect 34802 33070 34814 33122
rect 29374 33058 29426 33070
rect 35534 33058 35586 33070
rect 37662 33122 37714 33134
rect 42018 33070 42030 33122
rect 42082 33070 42094 33122
rect 37662 33058 37714 33070
rect 1344 32954 46592 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 46592 32954
rect 1344 32868 46592 32902
rect 5406 32786 5458 32798
rect 4722 32734 4734 32786
rect 4786 32734 4798 32786
rect 5406 32722 5458 32734
rect 8542 32786 8594 32798
rect 8542 32722 8594 32734
rect 12798 32786 12850 32798
rect 41022 32786 41074 32798
rect 38098 32734 38110 32786
rect 38162 32734 38174 32786
rect 39106 32734 39118 32786
rect 39170 32734 39182 32786
rect 12798 32722 12850 32734
rect 41022 32722 41074 32734
rect 8654 32674 8706 32686
rect 8654 32610 8706 32622
rect 12238 32674 12290 32686
rect 12238 32610 12290 32622
rect 22206 32674 22258 32686
rect 22206 32610 22258 32622
rect 22542 32674 22594 32686
rect 24546 32622 24558 32674
rect 24610 32622 24622 32674
rect 25666 32622 25678 32674
rect 25730 32622 25742 32674
rect 28690 32622 28702 32674
rect 28754 32622 28766 32674
rect 22542 32610 22594 32622
rect 1934 32562 1986 32574
rect 12574 32562 12626 32574
rect 21646 32562 21698 32574
rect 29374 32562 29426 32574
rect 32958 32562 33010 32574
rect 38782 32562 38834 32574
rect 2258 32510 2270 32562
rect 2322 32510 2334 32562
rect 12002 32510 12014 32562
rect 12066 32510 12078 32562
rect 13346 32510 13358 32562
rect 13410 32510 13422 32562
rect 13570 32510 13582 32562
rect 13634 32510 13646 32562
rect 17266 32510 17278 32562
rect 17330 32510 17342 32562
rect 17938 32510 17950 32562
rect 18002 32510 18014 32562
rect 21410 32510 21422 32562
rect 21474 32510 21486 32562
rect 24322 32510 24334 32562
rect 24386 32510 24398 32562
rect 25890 32510 25902 32562
rect 25954 32510 25966 32562
rect 28018 32510 28030 32562
rect 28082 32510 28094 32562
rect 28578 32510 28590 32562
rect 28642 32510 28654 32562
rect 29810 32510 29822 32562
rect 29874 32510 29886 32562
rect 30706 32510 30718 32562
rect 30770 32510 30782 32562
rect 33506 32510 33518 32562
rect 33570 32510 33582 32562
rect 36418 32510 36430 32562
rect 36482 32510 36494 32562
rect 36978 32510 36990 32562
rect 37042 32510 37054 32562
rect 37762 32510 37774 32562
rect 37826 32510 37838 32562
rect 38322 32510 38334 32562
rect 38386 32510 38398 32562
rect 1934 32498 1986 32510
rect 12574 32498 12626 32510
rect 21646 32498 21698 32510
rect 29374 32498 29426 32510
rect 32958 32498 33010 32510
rect 38782 32498 38834 32510
rect 39566 32562 39618 32574
rect 42690 32510 42702 32562
rect 42754 32510 42766 32562
rect 43138 32510 43150 32562
rect 43202 32510 43214 32562
rect 44034 32510 44046 32562
rect 44098 32510 44110 32562
rect 39566 32498 39618 32510
rect 11566 32450 11618 32462
rect 25342 32450 25394 32462
rect 20402 32398 20414 32450
rect 20466 32398 20478 32450
rect 11566 32386 11618 32398
rect 25342 32386 25394 32398
rect 26462 32450 26514 32462
rect 26462 32386 26514 32398
rect 27694 32450 27746 32462
rect 27694 32386 27746 32398
rect 32510 32450 32562 32462
rect 41794 32398 41806 32450
rect 41858 32398 41870 32450
rect 32510 32386 32562 32398
rect 16606 32338 16658 32350
rect 45166 32338 45218 32350
rect 21298 32286 21310 32338
rect 21362 32286 21374 32338
rect 24098 32286 24110 32338
rect 24162 32286 24174 32338
rect 16606 32274 16658 32286
rect 45166 32274 45218 32286
rect 1344 32170 46592 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 46592 32170
rect 1344 32084 46592 32118
rect 26898 31950 26910 32002
rect 26962 31950 26974 32002
rect 29810 31950 29822 32002
rect 29874 31950 29886 32002
rect 16158 31890 16210 31902
rect 12338 31838 12350 31890
rect 12402 31838 12414 31890
rect 16158 31826 16210 31838
rect 21310 31890 21362 31902
rect 37550 31890 37602 31902
rect 27794 31838 27806 31890
rect 27858 31838 27870 31890
rect 21310 31826 21362 31838
rect 37550 31826 37602 31838
rect 6974 31778 7026 31790
rect 11342 31778 11394 31790
rect 7410 31726 7422 31778
rect 7474 31726 7486 31778
rect 6974 31714 7026 31726
rect 11342 31714 11394 31726
rect 11566 31778 11618 31790
rect 15038 31778 15090 31790
rect 17614 31778 17666 31790
rect 19854 31778 19906 31790
rect 13570 31726 13582 31778
rect 13634 31726 13646 31778
rect 16594 31726 16606 31778
rect 16658 31726 16670 31778
rect 16930 31726 16942 31778
rect 16994 31726 17006 31778
rect 18162 31726 18174 31778
rect 18226 31726 18238 31778
rect 19282 31726 19294 31778
rect 19346 31726 19358 31778
rect 21746 31726 21758 31778
rect 21810 31726 21822 31778
rect 22082 31738 22094 31790
rect 22146 31738 22158 31790
rect 22766 31778 22818 31790
rect 26126 31778 26178 31790
rect 23314 31726 23326 31778
rect 23378 31726 23390 31778
rect 24322 31726 24334 31778
rect 24386 31726 24398 31778
rect 25218 31726 25230 31778
rect 25282 31726 25294 31778
rect 11566 31714 11618 31726
rect 15038 31714 15090 31726
rect 17614 31714 17666 31726
rect 19854 31714 19906 31726
rect 22766 31714 22818 31726
rect 26126 31714 26178 31726
rect 26350 31778 26402 31790
rect 28354 31726 28366 31778
rect 28418 31726 28430 31778
rect 29250 31726 29262 31778
rect 29314 31726 29326 31778
rect 32050 31726 32062 31778
rect 32114 31726 32126 31778
rect 32386 31726 32398 31778
rect 32450 31726 32462 31778
rect 34626 31726 34638 31778
rect 34690 31726 34702 31778
rect 38882 31726 38894 31778
rect 38946 31726 38958 31778
rect 39666 31726 39678 31778
rect 39730 31726 39742 31778
rect 26350 31714 26402 31726
rect 3950 31666 4002 31678
rect 3950 31602 4002 31614
rect 9662 31666 9714 31678
rect 9662 31602 9714 31614
rect 11902 31666 11954 31678
rect 11902 31602 11954 31614
rect 15374 31666 15426 31678
rect 15374 31602 15426 31614
rect 15710 31666 15762 31678
rect 26574 31666 26626 31678
rect 39454 31666 39506 31678
rect 17154 31614 17166 31666
rect 17218 31614 17230 31666
rect 20402 31614 20414 31666
rect 20466 31614 20478 31666
rect 25442 31614 25454 31666
rect 25506 31614 25518 31666
rect 36194 31614 36206 31666
rect 36258 31614 36270 31666
rect 15710 31602 15762 31614
rect 26574 31602 26626 31614
rect 39454 31602 39506 31614
rect 3838 31554 3890 31566
rect 3838 31490 3890 31502
rect 10446 31554 10498 31566
rect 10446 31490 10498 31502
rect 12798 31554 12850 31566
rect 12798 31490 12850 31502
rect 13806 31554 13858 31566
rect 13806 31490 13858 31502
rect 14478 31554 14530 31566
rect 20750 31554 20802 31566
rect 40238 31554 40290 31566
rect 14690 31502 14702 31554
rect 14754 31502 14766 31554
rect 22306 31502 22318 31554
rect 22370 31502 22382 31554
rect 25554 31502 25566 31554
rect 25618 31502 25630 31554
rect 14478 31490 14530 31502
rect 20750 31490 20802 31502
rect 40238 31490 40290 31502
rect 44942 31554 44994 31566
rect 44942 31490 44994 31502
rect 1344 31386 46592 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 46592 31386
rect 1344 31300 46592 31334
rect 5518 31218 5570 31230
rect 4834 31166 4846 31218
rect 4898 31166 4910 31218
rect 5518 31154 5570 31166
rect 8206 31218 8258 31230
rect 8206 31154 8258 31166
rect 18958 31218 19010 31230
rect 29150 31218 29202 31230
rect 22418 31166 22430 31218
rect 22482 31166 22494 31218
rect 18958 31154 19010 31166
rect 29150 31154 29202 31166
rect 34302 31218 34354 31230
rect 34302 31154 34354 31166
rect 41582 31218 41634 31230
rect 41582 31154 41634 31166
rect 41918 31218 41970 31230
rect 41918 31154 41970 31166
rect 8318 31106 8370 31118
rect 8318 31042 8370 31054
rect 14702 31106 14754 31118
rect 14702 31042 14754 31054
rect 15038 31106 15090 31118
rect 15038 31042 15090 31054
rect 15710 31106 15762 31118
rect 15710 31042 15762 31054
rect 16382 31106 16434 31118
rect 35870 31106 35922 31118
rect 21634 31054 21646 31106
rect 21698 31054 21710 31106
rect 26226 31054 26238 31106
rect 26290 31054 26302 31106
rect 28802 31054 28814 31106
rect 28866 31054 28878 31106
rect 34626 31054 34638 31106
rect 34690 31054 34702 31106
rect 36866 31054 36878 31106
rect 36930 31054 36942 31106
rect 42242 31054 42254 31106
rect 42306 31054 42318 31106
rect 43586 31054 43598 31106
rect 43650 31054 43662 31106
rect 16382 31042 16434 31054
rect 35870 31042 35922 31054
rect 2046 30994 2098 31006
rect 15374 30994 15426 31006
rect 2482 30942 2494 30994
rect 2546 30942 2558 30994
rect 13458 30942 13470 30994
rect 13522 30942 13534 30994
rect 2046 30930 2098 30942
rect 15374 30930 15426 30942
rect 16046 30994 16098 31006
rect 22206 30994 22258 31006
rect 34974 30994 35026 31006
rect 37550 30994 37602 31006
rect 20178 30942 20190 30994
rect 20242 30942 20254 30994
rect 22530 30942 22542 30994
rect 22594 30942 22606 30994
rect 23426 30942 23438 30994
rect 23490 30942 23502 30994
rect 25554 30942 25566 30994
rect 25618 30942 25630 30994
rect 26114 30942 26126 30994
rect 26178 30942 26190 30994
rect 26786 30942 26798 30994
rect 26850 30942 26862 30994
rect 27346 30942 27358 30994
rect 27410 30942 27422 30994
rect 28354 30942 28366 30994
rect 28418 30942 28430 30994
rect 29474 30942 29486 30994
rect 29538 30942 29550 30994
rect 36194 30942 36206 30994
rect 36258 30942 36270 30994
rect 36642 30942 36654 30994
rect 36706 30942 36718 30994
rect 37874 30942 37886 30994
rect 37938 30942 37950 30994
rect 38994 30942 39006 30994
rect 39058 30942 39070 30994
rect 39554 30942 39566 30994
rect 39618 30942 39630 30994
rect 45042 30942 45054 30994
rect 45106 30942 45118 30994
rect 16046 30930 16098 30942
rect 22206 30930 22258 30942
rect 34974 30930 35026 30942
rect 37550 30930 37602 30942
rect 16830 30882 16882 30894
rect 12002 30830 12014 30882
rect 12066 30830 12078 30882
rect 16830 30818 16882 30830
rect 17614 30882 17666 30894
rect 25230 30882 25282 30894
rect 33966 30882 34018 30894
rect 18498 30830 18510 30882
rect 18562 30830 18574 30882
rect 20402 30830 20414 30882
rect 20466 30830 20478 30882
rect 24546 30830 24558 30882
rect 24610 30830 24622 30882
rect 30706 30830 30718 30882
rect 30770 30830 30782 30882
rect 17614 30818 17666 30830
rect 25230 30818 25282 30830
rect 33966 30818 34018 30830
rect 35534 30882 35586 30894
rect 41022 30882 41074 30894
rect 39890 30830 39902 30882
rect 39954 30830 39966 30882
rect 43250 30830 43262 30882
rect 43314 30830 43326 30882
rect 45714 30830 45726 30882
rect 45778 30830 45790 30882
rect 35534 30818 35586 30830
rect 41022 30818 41074 30830
rect 1344 30602 46592 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 46592 30602
rect 1344 30516 46592 30550
rect 37438 30434 37490 30446
rect 37438 30370 37490 30382
rect 14926 30322 14978 30334
rect 20402 30270 20414 30322
rect 20466 30270 20478 30322
rect 14926 30258 14978 30270
rect 3726 30210 3778 30222
rect 13470 30210 13522 30222
rect 12114 30158 12126 30210
rect 12178 30158 12190 30210
rect 12898 30158 12910 30210
rect 12962 30158 12974 30210
rect 3726 30146 3778 30158
rect 13470 30146 13522 30158
rect 14030 30210 14082 30222
rect 22094 30210 22146 30222
rect 26350 30210 26402 30222
rect 29150 30210 29202 30222
rect 35534 30210 35586 30222
rect 45166 30210 45218 30222
rect 14578 30158 14590 30210
rect 14642 30158 14654 30210
rect 19506 30158 19518 30210
rect 19570 30158 19582 30210
rect 20066 30158 20078 30210
rect 20130 30158 20142 30210
rect 22530 30158 22542 30210
rect 22594 30158 22606 30210
rect 23426 30158 23438 30210
rect 23490 30158 23502 30210
rect 24322 30158 24334 30210
rect 24386 30158 24398 30210
rect 25218 30158 25230 30210
rect 25282 30158 25294 30210
rect 25778 30158 25790 30210
rect 25842 30158 25854 30210
rect 27122 30158 27134 30210
rect 27186 30158 27198 30210
rect 28018 30158 28030 30210
rect 28082 30158 28094 30210
rect 29810 30158 29822 30210
rect 29874 30158 29886 30210
rect 37874 30158 37886 30210
rect 37938 30158 37950 30210
rect 39330 30158 39342 30210
rect 39394 30158 39406 30210
rect 40786 30158 40798 30210
rect 40850 30158 40862 30210
rect 41010 30158 41022 30210
rect 41074 30158 41086 30210
rect 41682 30158 41694 30210
rect 41746 30158 41758 30210
rect 44258 30158 44270 30210
rect 44322 30158 44334 30210
rect 14030 30146 14082 30158
rect 22094 30146 22146 30158
rect 26350 30146 26402 30158
rect 29150 30146 29202 30158
rect 35534 30146 35586 30158
rect 45166 30146 45218 30158
rect 45838 30210 45890 30222
rect 45838 30146 45890 30158
rect 3838 30098 3890 30110
rect 24894 30098 24946 30110
rect 33742 30098 33794 30110
rect 17154 30046 17166 30098
rect 17218 30046 17230 30098
rect 21410 30046 21422 30098
rect 21474 30046 21486 30098
rect 23090 30046 23102 30098
rect 23154 30046 23166 30098
rect 30258 30046 30270 30098
rect 30322 30046 30334 30098
rect 3838 30034 3890 30046
rect 24894 30034 24946 30046
rect 33742 30034 33794 30046
rect 34078 30098 34130 30110
rect 34078 30034 34130 30046
rect 34414 30098 34466 30110
rect 34414 30034 34466 30046
rect 34750 30098 34802 30110
rect 38670 30098 38722 30110
rect 44830 30098 44882 30110
rect 35746 30046 35758 30098
rect 35810 30046 35822 30098
rect 36306 30046 36318 30098
rect 36370 30046 36382 30098
rect 38210 30046 38222 30098
rect 38274 30046 38286 30098
rect 42802 30046 42814 30098
rect 42866 30046 42878 30098
rect 34750 30034 34802 30046
rect 38670 30034 38722 30046
rect 44830 30034 44882 30046
rect 45502 30098 45554 30110
rect 45502 30034 45554 30046
rect 17838 29986 17890 29998
rect 17838 29922 17890 29934
rect 19518 29986 19570 29998
rect 19518 29922 19570 29934
rect 21758 29986 21810 29998
rect 30606 29986 30658 29998
rect 25890 29934 25902 29986
rect 25954 29934 25966 29986
rect 21758 29922 21810 29934
rect 30606 29922 30658 29934
rect 33518 29986 33570 29998
rect 33518 29922 33570 29934
rect 35198 29986 35250 29998
rect 35198 29922 35250 29934
rect 37102 29986 37154 29998
rect 37102 29922 37154 29934
rect 39006 29986 39058 29998
rect 42354 29934 42366 29986
rect 42418 29934 42430 29986
rect 39006 29922 39058 29934
rect 1344 29818 46592 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 46592 29818
rect 1344 29732 46592 29766
rect 5406 29650 5458 29662
rect 4834 29598 4846 29650
rect 4898 29598 4910 29650
rect 5406 29586 5458 29598
rect 5630 29650 5682 29662
rect 5630 29586 5682 29598
rect 16494 29650 16546 29662
rect 16494 29586 16546 29598
rect 17390 29650 17442 29662
rect 17390 29586 17442 29598
rect 21198 29650 21250 29662
rect 21198 29586 21250 29598
rect 23662 29650 23714 29662
rect 23662 29586 23714 29598
rect 24110 29650 24162 29662
rect 27694 29650 27746 29662
rect 25218 29598 25230 29650
rect 25282 29598 25294 29650
rect 27346 29598 27358 29650
rect 27410 29598 27422 29650
rect 24110 29586 24162 29598
rect 27694 29586 27746 29598
rect 33182 29650 33234 29662
rect 33182 29586 33234 29598
rect 45502 29650 45554 29662
rect 45502 29586 45554 29598
rect 5966 29538 6018 29550
rect 5966 29474 6018 29486
rect 17726 29538 17778 29550
rect 27806 29538 27858 29550
rect 34750 29538 34802 29550
rect 41918 29538 41970 29550
rect 19506 29486 19518 29538
rect 19570 29486 19582 29538
rect 33506 29486 33518 29538
rect 33570 29486 33582 29538
rect 34178 29486 34190 29538
rect 34242 29486 34254 29538
rect 38210 29486 38222 29538
rect 38274 29486 38286 29538
rect 42914 29486 42926 29538
rect 42978 29486 42990 29538
rect 17726 29474 17778 29486
rect 27806 29474 27858 29486
rect 34750 29474 34802 29486
rect 41918 29474 41970 29486
rect 20526 29426 20578 29438
rect 1810 29374 1822 29426
rect 1874 29374 1886 29426
rect 2258 29374 2270 29426
rect 2322 29374 2334 29426
rect 10770 29374 10782 29426
rect 10834 29374 10846 29426
rect 16706 29374 16718 29426
rect 16770 29374 16782 29426
rect 19170 29374 19182 29426
rect 19234 29374 19246 29426
rect 20526 29362 20578 29374
rect 20862 29426 20914 29438
rect 20862 29362 20914 29374
rect 23326 29426 23378 29438
rect 23326 29362 23378 29374
rect 25790 29426 25842 29438
rect 37214 29426 37266 29438
rect 41470 29426 41522 29438
rect 43598 29426 43650 29438
rect 26786 29374 26798 29426
rect 26850 29374 26862 29426
rect 28578 29374 28590 29426
rect 28642 29374 28654 29426
rect 29250 29374 29262 29426
rect 29314 29374 29326 29426
rect 31490 29374 31502 29426
rect 31554 29374 31566 29426
rect 31826 29374 31838 29426
rect 31890 29374 31902 29426
rect 36754 29374 36766 29426
rect 36818 29374 36830 29426
rect 41010 29374 41022 29426
rect 41074 29374 41086 29426
rect 42242 29374 42254 29426
rect 42306 29374 42318 29426
rect 42690 29374 42702 29426
rect 42754 29374 42766 29426
rect 43922 29374 43934 29426
rect 43986 29374 43998 29426
rect 44930 29374 44942 29426
rect 44994 29374 45006 29426
rect 25790 29362 25842 29374
rect 37214 29362 37266 29374
rect 41470 29362 41522 29374
rect 43598 29362 43650 29374
rect 21982 29314 22034 29326
rect 12786 29262 12798 29314
rect 12850 29262 12862 29314
rect 20066 29262 20078 29314
rect 20130 29262 20142 29314
rect 21982 29250 22034 29262
rect 22990 29314 23042 29326
rect 25566 29314 25618 29326
rect 37774 29314 37826 29326
rect 24546 29262 24558 29314
rect 24610 29262 24622 29314
rect 31154 29262 31166 29314
rect 31218 29262 31230 29314
rect 34626 29262 34638 29314
rect 34690 29262 34702 29314
rect 45938 29262 45950 29314
rect 46002 29262 46014 29314
rect 22990 29250 23042 29262
rect 25566 29250 25618 29262
rect 37774 29250 37826 29262
rect 18398 29202 18450 29214
rect 18398 29138 18450 29150
rect 18734 29202 18786 29214
rect 36094 29202 36146 29214
rect 30146 29150 30158 29202
rect 30210 29150 30222 29202
rect 31266 29150 31278 29202
rect 31330 29150 31342 29202
rect 18734 29138 18786 29150
rect 36094 29138 36146 29150
rect 40126 29202 40178 29214
rect 40126 29138 40178 29150
rect 1344 29034 46592 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 46592 29034
rect 1344 28948 46592 28982
rect 9214 28866 9266 28878
rect 9214 28802 9266 28814
rect 12014 28866 12066 28878
rect 12014 28802 12066 28814
rect 14926 28866 14978 28878
rect 14926 28802 14978 28814
rect 19630 28866 19682 28878
rect 19630 28802 19682 28814
rect 28142 28866 28194 28878
rect 43586 28814 43598 28866
rect 43650 28814 43662 28866
rect 45378 28814 45390 28866
rect 45442 28814 45454 28866
rect 28142 28802 28194 28814
rect 1934 28754 1986 28766
rect 22654 28754 22706 28766
rect 18386 28702 18398 28754
rect 18450 28702 18462 28754
rect 1934 28690 1986 28702
rect 22654 28690 22706 28702
rect 28366 28754 28418 28766
rect 28366 28690 28418 28702
rect 28590 28754 28642 28766
rect 36430 28754 36482 28766
rect 32946 28702 32958 28754
rect 33010 28702 33022 28754
rect 28590 28690 28642 28702
rect 36430 28690 36482 28702
rect 42702 28754 42754 28766
rect 42702 28690 42754 28702
rect 4958 28642 5010 28654
rect 4274 28590 4286 28642
rect 4338 28590 4350 28642
rect 4958 28578 5010 28590
rect 5630 28642 5682 28654
rect 5630 28578 5682 28590
rect 11678 28642 11730 28654
rect 22206 28642 22258 28654
rect 25006 28642 25058 28654
rect 12674 28590 12686 28642
rect 12738 28590 12750 28642
rect 14130 28590 14142 28642
rect 14194 28590 14206 28642
rect 14578 28590 14590 28642
rect 14642 28590 14654 28642
rect 19170 28590 19182 28642
rect 19234 28590 19246 28642
rect 23874 28590 23886 28642
rect 23938 28590 23950 28642
rect 24546 28590 24558 28642
rect 24610 28590 24622 28642
rect 11678 28578 11730 28590
rect 22206 28578 22258 28590
rect 25006 28578 25058 28590
rect 27694 28642 27746 28654
rect 27694 28578 27746 28590
rect 29262 28642 29314 28654
rect 35870 28642 35922 28654
rect 29698 28590 29710 28642
rect 29762 28590 29774 28642
rect 30146 28590 30158 28642
rect 30210 28590 30222 28642
rect 30818 28590 30830 28642
rect 30882 28590 30894 28642
rect 31266 28590 31278 28642
rect 31330 28590 31342 28642
rect 32274 28590 32286 28642
rect 32338 28590 32350 28642
rect 32834 28590 32846 28642
rect 32898 28590 32910 28642
rect 34514 28590 34526 28642
rect 34578 28590 34590 28642
rect 38434 28590 38446 28642
rect 38498 28590 38510 28642
rect 40674 28590 40686 28642
rect 40738 28590 40750 28642
rect 42466 28590 42478 28642
rect 42530 28590 42542 28642
rect 43138 28590 43150 28642
rect 43202 28590 43214 28642
rect 45602 28590 45614 28642
rect 45666 28590 45678 28642
rect 29262 28578 29314 28590
rect 35870 28578 35922 28590
rect 5742 28530 5794 28542
rect 10110 28530 10162 28542
rect 13918 28530 13970 28542
rect 21310 28530 21362 28542
rect 8530 28478 8542 28530
rect 8594 28478 8606 28530
rect 8978 28478 8990 28530
rect 9042 28478 9054 28530
rect 12786 28478 12798 28530
rect 12850 28478 12862 28530
rect 16818 28478 16830 28530
rect 16882 28478 16894 28530
rect 19058 28478 19070 28530
rect 19122 28478 19134 28530
rect 5742 28466 5794 28478
rect 10110 28466 10162 28478
rect 13918 28466 13970 28478
rect 21310 28466 21362 28478
rect 23102 28530 23154 28542
rect 44158 28530 44210 28542
rect 24322 28478 24334 28530
rect 24386 28478 24398 28530
rect 25330 28478 25342 28530
rect 25394 28478 25406 28530
rect 33618 28478 33630 28530
rect 33682 28478 33694 28530
rect 23102 28466 23154 28478
rect 44158 28466 44210 28478
rect 44830 28530 44882 28542
rect 44830 28466 44882 28478
rect 44942 28530 44994 28542
rect 45042 28478 45054 28530
rect 45106 28478 45118 28530
rect 44942 28466 44994 28478
rect 4622 28418 4674 28430
rect 4622 28354 4674 28366
rect 7870 28418 7922 28430
rect 7870 28354 7922 28366
rect 9550 28418 9602 28430
rect 9550 28354 9602 28366
rect 9998 28418 10050 28430
rect 9998 28354 10050 28366
rect 19966 28418 20018 28430
rect 19966 28354 20018 28366
rect 21422 28418 21474 28430
rect 21422 28354 21474 28366
rect 21646 28418 21698 28430
rect 21646 28354 21698 28366
rect 22094 28418 22146 28430
rect 22094 28354 22146 28366
rect 23214 28418 23266 28430
rect 23214 28354 23266 28366
rect 23438 28418 23490 28430
rect 37438 28418 37490 28430
rect 23650 28366 23662 28418
rect 23714 28366 23726 28418
rect 30258 28366 30270 28418
rect 30322 28366 30334 28418
rect 23438 28354 23490 28366
rect 37438 28354 37490 28366
rect 39678 28418 39730 28430
rect 39678 28354 39730 28366
rect 41806 28418 41858 28430
rect 41806 28354 41858 28366
rect 1344 28250 46592 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 46592 28250
rect 1344 28164 46592 28198
rect 5294 28082 5346 28094
rect 13470 28082 13522 28094
rect 23326 28082 23378 28094
rect 25342 28082 25394 28094
rect 4722 28030 4734 28082
rect 4786 28030 4798 28082
rect 10210 28030 10222 28082
rect 10274 28030 10286 28082
rect 21074 28030 21086 28082
rect 21138 28030 21150 28082
rect 23986 28030 23998 28082
rect 24050 28030 24062 28082
rect 5294 28018 5346 28030
rect 13470 28018 13522 28030
rect 23326 28018 23378 28030
rect 25342 28018 25394 28030
rect 28814 28082 28866 28094
rect 28814 28018 28866 28030
rect 33406 28082 33458 28094
rect 34962 28030 34974 28082
rect 35026 28030 35038 28082
rect 33406 28018 33458 28030
rect 6638 27970 6690 27982
rect 9550 27970 9602 27982
rect 7746 27918 7758 27970
rect 7810 27918 7822 27970
rect 6638 27906 6690 27918
rect 9550 27906 9602 27918
rect 15822 27970 15874 27982
rect 19406 27970 19458 27982
rect 25230 27970 25282 27982
rect 17602 27918 17614 27970
rect 17666 27918 17678 27970
rect 19058 27918 19070 27970
rect 19122 27918 19134 27970
rect 20962 27918 20974 27970
rect 21026 27918 21038 27970
rect 21858 27918 21870 27970
rect 21922 27918 21934 27970
rect 24322 27918 24334 27970
rect 24386 27918 24398 27970
rect 15822 27906 15874 27918
rect 19406 27906 19458 27918
rect 25230 27906 25282 27918
rect 26014 27970 26066 27982
rect 26014 27906 26066 27918
rect 26126 27970 26178 27982
rect 26126 27906 26178 27918
rect 27134 27970 27186 27982
rect 27134 27906 27186 27918
rect 27246 27970 27298 27982
rect 27246 27906 27298 27918
rect 32174 27970 32226 27982
rect 32174 27906 32226 27918
rect 33070 27970 33122 27982
rect 33070 27906 33122 27918
rect 35310 27970 35362 27982
rect 36306 27918 36318 27970
rect 36370 27918 36382 27970
rect 35310 27906 35362 27918
rect 6750 27858 6802 27870
rect 14030 27858 14082 27870
rect 23662 27858 23714 27870
rect 1698 27806 1710 27858
rect 1762 27806 1774 27858
rect 2258 27806 2270 27858
rect 2322 27806 2334 27858
rect 7186 27806 7198 27858
rect 7250 27806 7262 27858
rect 9762 27806 9774 27858
rect 9826 27806 9838 27858
rect 10434 27806 10446 27858
rect 10498 27806 10510 27858
rect 13234 27806 13246 27858
rect 13298 27806 13310 27858
rect 13794 27806 13806 27858
rect 13858 27806 13870 27858
rect 17490 27806 17502 27858
rect 17554 27806 17566 27858
rect 20178 27806 20190 27858
rect 20242 27806 20254 27858
rect 20850 27806 20862 27858
rect 20914 27806 20926 27858
rect 21746 27806 21758 27858
rect 21810 27806 21822 27858
rect 6750 27794 6802 27806
rect 14030 27794 14082 27806
rect 23662 27794 23714 27806
rect 24670 27858 24722 27870
rect 24670 27794 24722 27806
rect 25566 27858 25618 27870
rect 25566 27794 25618 27806
rect 26910 27858 26962 27870
rect 34302 27858 34354 27870
rect 36766 27858 36818 27870
rect 28578 27806 28590 27858
rect 28642 27806 28654 27858
rect 29810 27806 29822 27858
rect 29874 27806 29886 27858
rect 32386 27806 32398 27858
rect 32450 27806 32462 27858
rect 34738 27806 34750 27858
rect 34802 27806 34814 27858
rect 35746 27806 35758 27858
rect 35810 27806 35822 27858
rect 36082 27806 36094 27858
rect 36146 27806 36158 27858
rect 37426 27806 37438 27858
rect 37490 27806 37502 27858
rect 38322 27806 38334 27858
rect 38386 27806 38398 27858
rect 40114 27806 40126 27858
rect 40178 27806 40190 27858
rect 41010 27806 41022 27858
rect 41074 27806 41086 27858
rect 41906 27806 41918 27858
rect 41970 27806 41982 27858
rect 42914 27806 42926 27858
rect 42978 27806 42990 27858
rect 44034 27806 44046 27858
rect 44098 27806 44110 27858
rect 26910 27794 26962 27806
rect 34302 27794 34354 27806
rect 36766 27794 36818 27806
rect 33854 27746 33906 27758
rect 22866 27694 22878 27746
rect 22930 27694 22942 27746
rect 31490 27694 31502 27746
rect 31554 27694 31566 27746
rect 39554 27694 39566 27746
rect 39618 27694 39630 27746
rect 40002 27694 40014 27746
rect 40066 27694 40078 27746
rect 42802 27694 42814 27746
rect 42866 27694 42878 27746
rect 44482 27694 44494 27746
rect 44546 27694 44558 27746
rect 33854 27682 33906 27694
rect 8878 27634 8930 27646
rect 18286 27634 18338 27646
rect 16594 27582 16606 27634
rect 16658 27582 16670 27634
rect 8878 27570 8930 27582
rect 18286 27570 18338 27582
rect 18622 27634 18674 27646
rect 18622 27570 18674 27582
rect 26126 27634 26178 27646
rect 26126 27570 26178 27582
rect 39118 27634 39170 27646
rect 39118 27570 39170 27582
rect 1344 27466 46592 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 46592 27466
rect 1344 27380 46592 27414
rect 11566 27298 11618 27310
rect 11566 27234 11618 27246
rect 35422 27298 35474 27310
rect 35422 27234 35474 27246
rect 37438 27298 37490 27310
rect 38322 27246 38334 27298
rect 38386 27246 38398 27298
rect 37438 27234 37490 27246
rect 1934 27186 1986 27198
rect 1934 27122 1986 27134
rect 13806 27186 13858 27198
rect 13806 27122 13858 27134
rect 14926 27186 14978 27198
rect 14926 27122 14978 27134
rect 16494 27186 16546 27198
rect 24670 27186 24722 27198
rect 17602 27134 17614 27186
rect 17666 27134 17678 27186
rect 24322 27134 24334 27186
rect 24386 27134 24398 27186
rect 16494 27122 16546 27134
rect 24670 27122 24722 27134
rect 30382 27186 30434 27198
rect 30382 27122 30434 27134
rect 30718 27186 30770 27198
rect 30718 27122 30770 27134
rect 37214 27186 37266 27198
rect 37214 27122 37266 27134
rect 39566 27186 39618 27198
rect 39566 27122 39618 27134
rect 8094 27074 8146 27086
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 7858 27022 7870 27074
rect 7922 27022 7934 27074
rect 8094 27010 8146 27022
rect 11342 27074 11394 27086
rect 11342 27010 11394 27022
rect 11678 27074 11730 27086
rect 15486 27074 15538 27086
rect 23998 27074 24050 27086
rect 14466 27022 14478 27074
rect 14530 27022 14542 27074
rect 17378 27022 17390 27074
rect 17442 27022 17454 27074
rect 18722 27022 18734 27074
rect 18786 27022 18798 27074
rect 19394 27022 19406 27074
rect 19458 27022 19470 27074
rect 20514 27022 20526 27074
rect 20578 27022 20590 27074
rect 21522 27022 21534 27074
rect 21586 27022 21598 27074
rect 22194 27022 22206 27074
rect 22258 27022 22270 27074
rect 23090 27022 23102 27074
rect 23154 27022 23166 27074
rect 11678 27010 11730 27022
rect 15486 27010 15538 27022
rect 23998 27010 24050 27022
rect 24894 27074 24946 27086
rect 24894 27010 24946 27022
rect 25342 27074 25394 27086
rect 25342 27010 25394 27022
rect 25454 27074 25506 27086
rect 25454 27010 25506 27022
rect 25790 27074 25842 27086
rect 25790 27010 25842 27022
rect 26126 27074 26178 27086
rect 26126 27010 26178 27022
rect 26350 27074 26402 27086
rect 26350 27010 26402 27022
rect 28590 27074 28642 27086
rect 32174 27074 32226 27086
rect 37886 27074 37938 27086
rect 29362 27022 29374 27074
rect 29426 27022 29438 27074
rect 29922 27022 29934 27074
rect 29986 27022 29998 27074
rect 31154 27022 31166 27074
rect 31218 27022 31230 27074
rect 31490 27022 31502 27074
rect 31554 27022 31566 27074
rect 32946 27022 32958 27074
rect 33010 27022 33022 27074
rect 33842 27022 33854 27074
rect 33906 27022 33918 27074
rect 34514 27022 34526 27074
rect 34578 27022 34590 27074
rect 36082 27022 36094 27074
rect 36146 27022 36158 27074
rect 28590 27010 28642 27022
rect 32174 27010 32226 27022
rect 37886 27010 37938 27022
rect 38222 27074 38274 27086
rect 38894 27074 38946 27086
rect 38546 27022 38558 27074
rect 38610 27022 38622 27074
rect 40002 27022 40014 27074
rect 40066 27022 40078 27074
rect 40338 27022 40350 27074
rect 40402 27022 40414 27074
rect 41346 27022 41358 27074
rect 41410 27022 41422 27074
rect 41794 27022 41806 27074
rect 41858 27022 41870 27074
rect 42802 27022 42814 27074
rect 42866 27022 42878 27074
rect 38222 27010 38274 27022
rect 38894 27010 38946 27022
rect 4622 26962 4674 26974
rect 4622 26898 4674 26910
rect 4734 26962 4786 26974
rect 11006 26962 11058 26974
rect 9986 26910 9998 26962
rect 10050 26910 10062 26962
rect 4734 26898 4786 26910
rect 11006 26898 11058 26910
rect 11118 26962 11170 26974
rect 11118 26898 11170 26910
rect 14254 26962 14306 26974
rect 14254 26898 14306 26910
rect 17054 26962 17106 26974
rect 26014 26962 26066 26974
rect 28254 26962 28306 26974
rect 18834 26910 18846 26962
rect 18898 26910 18910 26962
rect 19282 26910 19294 26962
rect 19346 26910 19358 26962
rect 21410 26910 21422 26962
rect 21474 26910 21486 26962
rect 22082 26910 22094 26962
rect 22146 26910 22158 26962
rect 27570 26910 27582 26962
rect 27634 26910 27646 26962
rect 17054 26898 17106 26910
rect 26014 26898 26066 26910
rect 28254 26898 28306 26910
rect 29150 26962 29202 26974
rect 38110 26962 38162 26974
rect 31714 26910 31726 26962
rect 31778 26910 31790 26962
rect 34290 26910 34302 26962
rect 34354 26910 34366 26962
rect 36194 26910 36206 26962
rect 36258 26910 36270 26962
rect 39218 26910 39230 26962
rect 39282 26910 39294 26962
rect 29150 26898 29202 26910
rect 38110 26898 38162 26910
rect 10670 26850 10722 26862
rect 10670 26786 10722 26798
rect 16270 26850 16322 26862
rect 25230 26850 25282 26862
rect 19170 26798 19182 26850
rect 19234 26798 19246 26850
rect 22194 26798 22206 26850
rect 22258 26798 22270 26850
rect 16270 26786 16322 26798
rect 25230 26786 25282 26798
rect 27918 26850 27970 26862
rect 27918 26786 27970 26798
rect 35086 26850 35138 26862
rect 35086 26786 35138 26798
rect 40686 26850 40738 26862
rect 40686 26786 40738 26798
rect 1344 26682 46592 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 46592 26682
rect 1344 26596 46592 26630
rect 9662 26514 9714 26526
rect 9662 26450 9714 26462
rect 19742 26514 19794 26526
rect 19742 26450 19794 26462
rect 24110 26514 24162 26526
rect 24110 26450 24162 26462
rect 24782 26514 24834 26526
rect 24782 26450 24834 26462
rect 27470 26514 27522 26526
rect 33070 26514 33122 26526
rect 28018 26462 28030 26514
rect 28082 26462 28094 26514
rect 30258 26462 30270 26514
rect 30322 26462 30334 26514
rect 27470 26450 27522 26462
rect 33070 26450 33122 26462
rect 35758 26514 35810 26526
rect 35758 26450 35810 26462
rect 36430 26514 36482 26526
rect 36430 26450 36482 26462
rect 39678 26514 39730 26526
rect 39678 26450 39730 26462
rect 43822 26514 43874 26526
rect 44146 26462 44158 26514
rect 44210 26462 44222 26514
rect 43822 26450 43874 26462
rect 5406 26402 5458 26414
rect 22430 26402 22482 26414
rect 10210 26350 10222 26402
rect 10274 26350 10286 26402
rect 10658 26350 10670 26402
rect 10722 26350 10734 26402
rect 21298 26350 21310 26402
rect 21362 26350 21374 26402
rect 21970 26350 21982 26402
rect 22034 26350 22046 26402
rect 5406 26338 5458 26350
rect 22430 26338 22482 26350
rect 24446 26402 24498 26414
rect 24446 26338 24498 26350
rect 24558 26402 24610 26414
rect 33742 26402 33794 26414
rect 26338 26350 26350 26402
rect 26402 26350 26414 26402
rect 24558 26338 24610 26350
rect 33742 26338 33794 26350
rect 2718 26290 2770 26302
rect 6414 26290 6466 26302
rect 3154 26238 3166 26290
rect 3218 26238 3230 26290
rect 2718 26226 2770 26238
rect 6414 26226 6466 26238
rect 6974 26290 7026 26302
rect 9998 26290 10050 26302
rect 17950 26290 18002 26302
rect 23550 26290 23602 26302
rect 28366 26290 28418 26302
rect 30942 26290 30994 26302
rect 37774 26290 37826 26302
rect 8194 26238 8206 26290
rect 8258 26238 8270 26290
rect 11666 26238 11678 26290
rect 11730 26238 11742 26290
rect 17490 26238 17502 26290
rect 17554 26238 17566 26290
rect 18610 26238 18622 26290
rect 18674 26238 18686 26290
rect 18834 26238 18846 26290
rect 18898 26238 18910 26290
rect 20178 26238 20190 26290
rect 20242 26238 20254 26290
rect 20850 26238 20862 26290
rect 20914 26238 20926 26290
rect 21746 26238 21758 26290
rect 21810 26238 21822 26290
rect 22530 26238 22542 26290
rect 22594 26238 22606 26290
rect 22978 26238 22990 26290
rect 23042 26238 23054 26290
rect 25218 26238 25230 26290
rect 25282 26238 25294 26290
rect 25666 26238 25678 26290
rect 25730 26238 25742 26290
rect 26786 26238 26798 26290
rect 26850 26238 26862 26290
rect 27794 26238 27806 26290
rect 27858 26238 27870 26290
rect 29698 26238 29710 26290
rect 29762 26238 29774 26290
rect 30146 26238 30158 26290
rect 30210 26238 30222 26290
rect 31266 26238 31278 26290
rect 31330 26238 31342 26290
rect 32386 26238 32398 26290
rect 32450 26238 32462 26290
rect 33282 26238 33294 26290
rect 33346 26238 33358 26290
rect 33954 26238 33966 26290
rect 34018 26238 34030 26290
rect 34850 26238 34862 26290
rect 34914 26238 34926 26290
rect 37090 26238 37102 26290
rect 37154 26238 37166 26290
rect 38770 26238 38782 26290
rect 38834 26238 38846 26290
rect 6974 26226 7026 26238
rect 9998 26226 10050 26238
rect 17950 26226 18002 26238
rect 23550 26226 23602 26238
rect 28366 26226 28418 26238
rect 30942 26226 30994 26238
rect 37774 26226 37826 26238
rect 26126 26178 26178 26190
rect 8642 26126 8654 26178
rect 8706 26126 8718 26178
rect 11330 26126 11342 26178
rect 11394 26126 11406 26178
rect 19394 26126 19406 26178
rect 19458 26126 19470 26178
rect 26126 26114 26178 26126
rect 28926 26178 28978 26190
rect 28926 26114 28978 26126
rect 29262 26178 29314 26190
rect 35186 26126 35198 26178
rect 35250 26126 35262 26178
rect 36754 26126 36766 26178
rect 36818 26126 36830 26178
rect 38210 26126 38222 26178
rect 38274 26126 38286 26178
rect 39106 26126 39118 26178
rect 39170 26126 39182 26178
rect 29262 26114 29314 26126
rect 6190 26066 6242 26078
rect 8082 26014 8094 26066
rect 8146 26014 8158 26066
rect 18498 26014 18510 26066
rect 18562 26014 18574 26066
rect 6190 26002 6242 26014
rect 1344 25898 46592 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 46592 25898
rect 1344 25812 46592 25846
rect 1934 25730 1986 25742
rect 1934 25666 1986 25678
rect 4622 25730 4674 25742
rect 4622 25666 4674 25678
rect 26574 25730 26626 25742
rect 26574 25666 26626 25678
rect 5854 25618 5906 25630
rect 13694 25618 13746 25630
rect 25006 25618 25058 25630
rect 34862 25618 34914 25630
rect 40126 25618 40178 25630
rect 12114 25566 12126 25618
rect 12178 25566 12190 25618
rect 16930 25566 16942 25618
rect 16994 25566 17006 25618
rect 31266 25566 31278 25618
rect 31330 25566 31342 25618
rect 37314 25566 37326 25618
rect 37378 25566 37390 25618
rect 45266 25566 45278 25618
rect 45330 25566 45342 25618
rect 5854 25554 5906 25566
rect 13694 25554 13746 25566
rect 25006 25554 25058 25566
rect 34862 25554 34914 25566
rect 40126 25554 40178 25566
rect 17614 25506 17666 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 7746 25454 7758 25506
rect 7810 25454 7822 25506
rect 9202 25454 9214 25506
rect 9266 25454 9278 25506
rect 14018 25454 14030 25506
rect 14082 25454 14094 25506
rect 17614 25442 17666 25454
rect 18062 25506 18114 25518
rect 19854 25506 19906 25518
rect 23774 25506 23826 25518
rect 18498 25454 18510 25506
rect 18562 25454 18574 25506
rect 19058 25454 19070 25506
rect 19122 25454 19134 25506
rect 19394 25454 19406 25506
rect 19458 25454 19470 25506
rect 20514 25454 20526 25506
rect 20578 25454 20590 25506
rect 21298 25454 21310 25506
rect 21362 25454 21374 25506
rect 22306 25454 22318 25506
rect 22370 25454 22382 25506
rect 23090 25454 23102 25506
rect 23154 25454 23166 25506
rect 18062 25442 18114 25454
rect 19854 25442 19906 25454
rect 23774 25442 23826 25454
rect 24110 25506 24162 25518
rect 25342 25506 25394 25518
rect 24546 25454 24558 25506
rect 24610 25454 24622 25506
rect 24110 25442 24162 25454
rect 25342 25442 25394 25454
rect 25566 25506 25618 25518
rect 28254 25506 28306 25518
rect 36430 25506 36482 25518
rect 44830 25506 44882 25518
rect 26226 25454 26238 25506
rect 26290 25454 26302 25506
rect 30034 25454 30046 25506
rect 30098 25454 30110 25506
rect 40898 25454 40910 25506
rect 40962 25454 40974 25506
rect 41346 25454 41358 25506
rect 41410 25454 41422 25506
rect 42466 25454 42478 25506
rect 42530 25454 42542 25506
rect 43474 25454 43486 25506
rect 43538 25454 43550 25506
rect 25566 25442 25618 25454
rect 28254 25442 28306 25454
rect 36430 25442 36482 25454
rect 44830 25442 44882 25454
rect 4734 25394 4786 25406
rect 4734 25330 4786 25342
rect 8542 25394 8594 25406
rect 8542 25330 8594 25342
rect 8878 25394 8930 25406
rect 17726 25394 17778 25406
rect 25902 25394 25954 25406
rect 40462 25394 40514 25406
rect 9986 25342 9998 25394
rect 10050 25342 10062 25394
rect 12450 25342 12462 25394
rect 12514 25342 12526 25394
rect 14802 25342 14814 25394
rect 14866 25342 14878 25394
rect 20402 25342 20414 25394
rect 20466 25342 20478 25394
rect 22418 25342 22430 25394
rect 22482 25342 22494 25394
rect 23426 25342 23438 25394
rect 23490 25342 23502 25394
rect 27906 25342 27918 25394
rect 27970 25342 27982 25394
rect 8878 25330 8930 25342
rect 17726 25330 17778 25342
rect 25902 25330 25954 25342
rect 40462 25330 40514 25342
rect 41918 25394 41970 25406
rect 41918 25330 41970 25342
rect 12798 25282 12850 25294
rect 12798 25218 12850 25230
rect 21198 25282 21250 25294
rect 21198 25218 21250 25230
rect 23998 25282 24050 25294
rect 23998 25218 24050 25230
rect 25454 25282 25506 25294
rect 25454 25218 25506 25230
rect 26462 25282 26514 25294
rect 27246 25282 27298 25294
rect 26898 25230 26910 25282
rect 26962 25230 26974 25282
rect 26462 25218 26514 25230
rect 27246 25218 27298 25230
rect 27582 25282 27634 25294
rect 27582 25218 27634 25230
rect 28590 25282 28642 25294
rect 28590 25218 28642 25230
rect 37774 25282 37826 25294
rect 38446 25282 38498 25294
rect 39118 25282 39170 25294
rect 38098 25230 38110 25282
rect 38162 25230 38174 25282
rect 38770 25230 38782 25282
rect 38834 25230 38846 25282
rect 37774 25218 37826 25230
rect 38446 25218 38498 25230
rect 39118 25218 39170 25230
rect 39678 25282 39730 25294
rect 41458 25230 41470 25282
rect 41522 25230 41534 25282
rect 39678 25218 39730 25230
rect 1344 25114 46592 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 46592 25114
rect 1344 25028 46592 25062
rect 6638 24946 6690 24958
rect 6638 24882 6690 24894
rect 10110 24946 10162 24958
rect 10110 24882 10162 24894
rect 10782 24946 10834 24958
rect 10782 24882 10834 24894
rect 12462 24946 12514 24958
rect 12462 24882 12514 24894
rect 19182 24946 19234 24958
rect 19182 24882 19234 24894
rect 32286 24946 32338 24958
rect 32286 24882 32338 24894
rect 33630 24946 33682 24958
rect 35186 24894 35198 24946
rect 35250 24894 35262 24946
rect 33630 24882 33682 24894
rect 5070 24834 5122 24846
rect 5070 24770 5122 24782
rect 6974 24834 7026 24846
rect 9550 24834 9602 24846
rect 12350 24834 12402 24846
rect 8418 24782 8430 24834
rect 8482 24782 8494 24834
rect 8866 24782 8878 24834
rect 8930 24782 8942 24834
rect 11330 24782 11342 24834
rect 11394 24782 11406 24834
rect 11778 24782 11790 24834
rect 11842 24782 11854 24834
rect 6974 24770 7026 24782
rect 9550 24770 9602 24782
rect 12350 24770 12402 24782
rect 13358 24834 13410 24846
rect 27470 24834 27522 24846
rect 35646 24834 35698 24846
rect 44494 24834 44546 24846
rect 19730 24782 19742 24834
rect 19794 24782 19806 24834
rect 20178 24782 20190 24834
rect 20242 24782 20254 24834
rect 22866 24782 22878 24834
rect 22930 24782 22942 24834
rect 26338 24782 26350 24834
rect 26402 24782 26414 24834
rect 29250 24782 29262 24834
rect 29314 24782 29326 24834
rect 39666 24782 39678 24834
rect 39730 24782 39742 24834
rect 40226 24782 40238 24834
rect 40290 24782 40302 24834
rect 41906 24782 41918 24834
rect 41970 24782 41982 24834
rect 13358 24770 13410 24782
rect 27470 24770 27522 24782
rect 35646 24770 35698 24782
rect 44494 24770 44546 24782
rect 7310 24722 7362 24734
rect 2258 24670 2270 24722
rect 2322 24670 2334 24722
rect 2706 24670 2718 24722
rect 2770 24670 2782 24722
rect 6402 24670 6414 24722
rect 6466 24670 6478 24722
rect 7310 24658 7362 24670
rect 7758 24722 7810 24734
rect 7758 24658 7810 24670
rect 8094 24722 8146 24734
rect 8094 24658 8146 24670
rect 11118 24722 11170 24734
rect 11118 24658 11170 24670
rect 12574 24722 12626 24734
rect 12574 24658 12626 24670
rect 13022 24722 13074 24734
rect 13022 24658 13074 24670
rect 13246 24722 13298 24734
rect 13246 24658 13298 24670
rect 16718 24722 16770 24734
rect 18622 24722 18674 24734
rect 26126 24722 26178 24734
rect 31726 24722 31778 24734
rect 38334 24722 38386 24734
rect 17826 24670 17838 24722
rect 17890 24670 17902 24722
rect 19506 24670 19518 24722
rect 19570 24670 19582 24722
rect 20514 24670 20526 24722
rect 20578 24670 20590 24722
rect 20962 24670 20974 24722
rect 21026 24670 21038 24722
rect 21858 24670 21870 24722
rect 21922 24670 21934 24722
rect 22530 24670 22542 24722
rect 22594 24670 22606 24722
rect 23874 24670 23886 24722
rect 23938 24670 23950 24722
rect 24210 24670 24222 24722
rect 24274 24670 24286 24722
rect 25666 24670 25678 24722
rect 25730 24670 25742 24722
rect 26786 24670 26798 24722
rect 26850 24670 26862 24722
rect 27122 24670 27134 24722
rect 27186 24670 27198 24722
rect 30034 24670 30046 24722
rect 30098 24670 30110 24722
rect 34514 24670 34526 24722
rect 34578 24670 34590 24722
rect 34962 24670 34974 24722
rect 35026 24670 35038 24722
rect 36306 24670 36318 24722
rect 36370 24670 36382 24722
rect 37202 24670 37214 24722
rect 37266 24670 37278 24722
rect 16718 24658 16770 24670
rect 18622 24658 18674 24670
rect 26126 24658 26178 24670
rect 31726 24658 31778 24670
rect 38334 24658 38386 24670
rect 39454 24722 39506 24734
rect 42590 24722 42642 24734
rect 45502 24722 45554 24734
rect 41234 24670 41246 24722
rect 41298 24670 41310 24722
rect 41794 24670 41806 24722
rect 41858 24670 41870 24722
rect 42914 24670 42926 24722
rect 42978 24670 42990 24722
rect 44034 24670 44046 24722
rect 44098 24670 44110 24722
rect 44706 24670 44718 24722
rect 44770 24670 44782 24722
rect 45714 24670 45726 24722
rect 45778 24670 45790 24722
rect 39454 24658 39506 24670
rect 42590 24658 42642 24670
rect 45502 24658 45554 24670
rect 1822 24610 1874 24622
rect 1822 24546 1874 24558
rect 5854 24610 5906 24622
rect 22206 24610 22258 24622
rect 18162 24558 18174 24610
rect 18226 24558 18238 24610
rect 5854 24546 5906 24558
rect 22206 24546 22258 24558
rect 22318 24610 22370 24622
rect 26014 24610 26066 24622
rect 23986 24558 23998 24610
rect 24050 24558 24062 24610
rect 22318 24546 22370 24558
rect 26014 24546 26066 24558
rect 33070 24610 33122 24622
rect 33070 24546 33122 24558
rect 34190 24610 34242 24622
rect 39118 24610 39170 24622
rect 37874 24558 37886 24610
rect 37938 24558 37950 24610
rect 34190 24546 34242 24558
rect 39118 24546 39170 24558
rect 40910 24610 40962 24622
rect 40910 24546 40962 24558
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 16830 24498 16882 24510
rect 27134 24498 27186 24510
rect 23538 24446 23550 24498
rect 23602 24446 23614 24498
rect 44818 24446 44830 24498
rect 44882 24446 44894 24498
rect 16830 24434 16882 24446
rect 27134 24434 27186 24446
rect 1344 24330 46592 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 46592 24330
rect 1344 24244 46592 24278
rect 30606 24162 30658 24174
rect 2818 24110 2830 24162
rect 2882 24110 2894 24162
rect 38434 24110 38446 24162
rect 38498 24110 38510 24162
rect 30606 24098 30658 24110
rect 14590 24050 14642 24062
rect 14590 23986 14642 23998
rect 15374 24050 15426 24062
rect 27806 24050 27858 24062
rect 18610 23998 18622 24050
rect 18674 23998 18686 24050
rect 19282 23998 19294 24050
rect 19346 23998 19358 24050
rect 15374 23986 15426 23998
rect 27806 23986 27858 23998
rect 28366 24050 28418 24062
rect 28366 23986 28418 23998
rect 29598 24050 29650 24062
rect 41918 24050 41970 24062
rect 31826 23998 31838 24050
rect 31890 23998 31902 24050
rect 37202 23998 37214 24050
rect 37266 23998 37278 24050
rect 45266 23998 45278 24050
rect 45330 23998 45342 24050
rect 29598 23986 29650 23998
rect 41918 23986 41970 23998
rect 14478 23938 14530 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 4946 23886 4958 23938
rect 5010 23886 5022 23938
rect 5618 23886 5630 23938
rect 5682 23886 5694 23938
rect 10098 23886 10110 23938
rect 10162 23886 10174 23938
rect 10546 23886 10558 23938
rect 10610 23886 10622 23938
rect 11890 23886 11902 23938
rect 11954 23886 11966 23938
rect 12786 23886 12798 23938
rect 12850 23886 12862 23938
rect 14478 23874 14530 23886
rect 14702 23938 14754 23950
rect 26798 23938 26850 23950
rect 29822 23938 29874 23950
rect 15698 23886 15710 23938
rect 15762 23886 15774 23938
rect 19618 23886 19630 23938
rect 19682 23886 19694 23938
rect 20178 23886 20190 23938
rect 20242 23886 20254 23938
rect 20738 23886 20750 23938
rect 20802 23886 20814 23938
rect 21970 23886 21982 23938
rect 22034 23886 22046 23938
rect 22642 23886 22654 23938
rect 22706 23886 22718 23938
rect 23314 23886 23326 23938
rect 23378 23886 23390 23938
rect 24322 23886 24334 23938
rect 24386 23886 24398 23938
rect 24994 23886 25006 23938
rect 25058 23886 25070 23938
rect 25330 23886 25342 23938
rect 25394 23886 25406 23938
rect 26450 23886 26462 23938
rect 26514 23886 26526 23938
rect 27458 23886 27470 23938
rect 27522 23886 27534 23938
rect 14702 23874 14754 23886
rect 26798 23874 26850 23886
rect 29822 23874 29874 23886
rect 29934 23938 29986 23950
rect 29934 23874 29986 23886
rect 30382 23938 30434 23950
rect 30382 23874 30434 23886
rect 31054 23938 31106 23950
rect 31054 23874 31106 23886
rect 32286 23938 32338 23950
rect 34862 23938 34914 23950
rect 40462 23938 40514 23950
rect 44830 23938 44882 23950
rect 33618 23886 33630 23938
rect 33682 23886 33694 23938
rect 33954 23886 33966 23938
rect 34018 23886 34030 23938
rect 35410 23886 35422 23938
rect 35474 23886 35486 23938
rect 36194 23886 36206 23938
rect 36258 23886 36270 23938
rect 37426 23886 37438 23938
rect 37490 23886 37502 23938
rect 37762 23886 37774 23938
rect 37826 23886 37838 23938
rect 38770 23886 38782 23938
rect 38834 23886 38846 23938
rect 41122 23886 41134 23938
rect 41186 23886 41198 23938
rect 42578 23886 42590 23938
rect 42642 23886 42654 23938
rect 43026 23886 43038 23938
rect 43090 23886 43102 23938
rect 44146 23886 44158 23938
rect 44210 23886 44222 23938
rect 45938 23886 45950 23938
rect 46002 23886 46014 23938
rect 32286 23874 32338 23886
rect 34862 23874 34914 23886
rect 40462 23874 40514 23886
rect 44830 23874 44882 23886
rect 8654 23826 8706 23838
rect 8654 23762 8706 23774
rect 9662 23826 9714 23838
rect 9662 23762 9714 23774
rect 11118 23826 11170 23838
rect 11118 23762 11170 23774
rect 14142 23826 14194 23838
rect 24558 23826 24610 23838
rect 33182 23826 33234 23838
rect 36990 23826 37042 23838
rect 40798 23826 40850 23838
rect 16482 23774 16494 23826
rect 16546 23774 16558 23826
rect 19282 23774 19294 23826
rect 19346 23774 19358 23826
rect 22866 23774 22878 23826
rect 22930 23774 22942 23826
rect 23650 23774 23662 23826
rect 23714 23774 23726 23826
rect 25778 23774 25790 23826
rect 25842 23774 25854 23826
rect 26338 23774 26350 23826
rect 26402 23774 26414 23826
rect 32610 23774 32622 23826
rect 32674 23774 32686 23826
rect 34178 23774 34190 23826
rect 34242 23774 34254 23826
rect 38994 23774 39006 23826
rect 39058 23774 39070 23826
rect 14142 23762 14194 23774
rect 24558 23762 24610 23774
rect 33182 23762 33234 23774
rect 36990 23762 37042 23774
rect 40798 23762 40850 23774
rect 4734 23714 4786 23726
rect 4734 23650 4786 23662
rect 6638 23714 6690 23726
rect 6638 23650 6690 23662
rect 8542 23714 8594 23726
rect 21422 23714 21474 23726
rect 27694 23714 27746 23726
rect 10658 23662 10670 23714
rect 10722 23662 10734 23714
rect 27122 23662 27134 23714
rect 27186 23662 27198 23714
rect 8542 23650 8594 23662
rect 21422 23650 21474 23662
rect 27694 23650 27746 23662
rect 29374 23714 29426 23726
rect 29374 23650 29426 23662
rect 31390 23714 31442 23726
rect 31390 23650 31442 23662
rect 37214 23714 37266 23726
rect 37214 23650 37266 23662
rect 41582 23714 41634 23726
rect 45714 23662 45726 23714
rect 45778 23662 45790 23714
rect 41582 23650 41634 23662
rect 1344 23546 46592 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 46592 23546
rect 1344 23460 46592 23494
rect 5854 23378 5906 23390
rect 4834 23326 4846 23378
rect 4898 23326 4910 23378
rect 5854 23314 5906 23326
rect 7646 23378 7698 23390
rect 7646 23314 7698 23326
rect 14926 23378 14978 23390
rect 14926 23314 14978 23326
rect 15934 23378 15986 23390
rect 15934 23314 15986 23326
rect 20750 23378 20802 23390
rect 26462 23378 26514 23390
rect 27918 23378 27970 23390
rect 23986 23326 23998 23378
rect 24050 23326 24062 23378
rect 27458 23326 27470 23378
rect 27522 23326 27534 23378
rect 20750 23314 20802 23326
rect 26462 23314 26514 23326
rect 27918 23314 27970 23326
rect 31838 23378 31890 23390
rect 31838 23314 31890 23326
rect 32286 23378 32338 23390
rect 32286 23314 32338 23326
rect 42030 23378 42082 23390
rect 42030 23314 42082 23326
rect 9662 23266 9714 23278
rect 16606 23266 16658 23278
rect 25678 23266 25730 23278
rect 6962 23214 6974 23266
rect 7026 23214 7038 23266
rect 8754 23214 8766 23266
rect 8818 23214 8830 23266
rect 10658 23214 10670 23266
rect 10722 23214 10734 23266
rect 23538 23214 23550 23266
rect 23602 23214 23614 23266
rect 24546 23214 24558 23266
rect 24610 23214 24622 23266
rect 9662 23202 9714 23214
rect 16606 23202 16658 23214
rect 25678 23202 25730 23214
rect 29038 23266 29090 23278
rect 31502 23266 31554 23278
rect 30594 23214 30606 23266
rect 30658 23214 30670 23266
rect 31042 23214 31054 23266
rect 31106 23214 31118 23266
rect 44482 23214 44494 23266
rect 44546 23214 44558 23266
rect 29038 23202 29090 23214
rect 31502 23202 31554 23214
rect 5518 23154 5570 23166
rect 1922 23102 1934 23154
rect 1986 23102 1998 23154
rect 2370 23102 2382 23154
rect 2434 23102 2446 23154
rect 5518 23090 5570 23102
rect 6190 23154 6242 23166
rect 7982 23154 8034 23166
rect 11118 23154 11170 23166
rect 14142 23154 14194 23166
rect 6850 23102 6862 23154
rect 6914 23102 6926 23154
rect 8418 23102 8430 23154
rect 8482 23102 8494 23154
rect 10098 23102 10110 23154
rect 10162 23102 10174 23154
rect 10434 23102 10446 23154
rect 10498 23102 10510 23154
rect 11890 23102 11902 23154
rect 11954 23102 11966 23154
rect 12786 23102 12798 23154
rect 12850 23102 12862 23154
rect 6190 23090 6242 23102
rect 7982 23090 8034 23102
rect 11118 23090 11170 23102
rect 14142 23090 14194 23102
rect 14814 23154 14866 23166
rect 14814 23090 14866 23102
rect 15598 23154 15650 23166
rect 25230 23154 25282 23166
rect 16370 23102 16382 23154
rect 16434 23102 16446 23154
rect 17378 23102 17390 23154
rect 17442 23102 17454 23154
rect 21186 23102 21198 23154
rect 21250 23102 21262 23154
rect 21410 23102 21422 23154
rect 21474 23102 21486 23154
rect 22530 23102 22542 23154
rect 22594 23102 22606 23154
rect 23426 23102 23438 23154
rect 23490 23102 23502 23154
rect 24210 23102 24222 23154
rect 24274 23102 24286 23154
rect 15598 23090 15650 23102
rect 25230 23090 25282 23102
rect 25902 23154 25954 23166
rect 25902 23090 25954 23102
rect 26238 23154 26290 23166
rect 28702 23154 28754 23166
rect 33854 23154 33906 23166
rect 35758 23154 35810 23166
rect 26786 23102 26798 23154
rect 26850 23102 26862 23154
rect 27234 23102 27246 23154
rect 27298 23102 27310 23154
rect 33506 23102 33518 23154
rect 33570 23102 33582 23154
rect 34962 23102 34974 23154
rect 35026 23102 35038 23154
rect 36194 23102 36206 23154
rect 36258 23102 36270 23154
rect 38994 23102 39006 23154
rect 39058 23102 39070 23154
rect 42578 23102 42590 23154
rect 42642 23102 42654 23154
rect 44930 23102 44942 23154
rect 44994 23102 45006 23154
rect 45490 23102 45502 23154
rect 45554 23102 45566 23154
rect 26238 23090 26290 23102
rect 28702 23090 28754 23102
rect 33854 23090 33906 23102
rect 35758 23090 35810 23102
rect 14478 23042 14530 23054
rect 25790 23042 25842 23054
rect 18162 22990 18174 23042
rect 18226 22990 18238 23042
rect 20290 22990 20302 23042
rect 20354 22990 20366 23042
rect 21522 22990 21534 23042
rect 21586 22990 21598 23042
rect 14478 22978 14530 22990
rect 25790 22978 25842 22990
rect 26350 23042 26402 23054
rect 26350 22978 26402 22990
rect 28366 23042 28418 23054
rect 33170 22990 33182 23042
rect 33234 22990 33246 23042
rect 38546 22990 38558 23042
rect 38610 22990 38622 23042
rect 28366 22978 28418 22990
rect 14926 22930 14978 22942
rect 14926 22866 14978 22878
rect 29486 22930 29538 22942
rect 29486 22866 29538 22878
rect 30270 22930 30322 22942
rect 36418 22878 36430 22930
rect 36482 22878 36494 22930
rect 30270 22866 30322 22878
rect 1344 22762 46592 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 46592 22762
rect 1344 22676 46592 22710
rect 9550 22594 9602 22606
rect 9550 22530 9602 22542
rect 9886 22594 9938 22606
rect 9886 22530 9938 22542
rect 13806 22594 13858 22606
rect 37102 22594 37154 22606
rect 32386 22542 32398 22594
rect 32450 22542 32462 22594
rect 13806 22530 13858 22542
rect 37102 22530 37154 22542
rect 37438 22594 37490 22606
rect 37438 22530 37490 22542
rect 11678 22482 11730 22494
rect 2034 22430 2046 22482
rect 2098 22430 2110 22482
rect 11678 22418 11730 22430
rect 13694 22482 13746 22494
rect 15710 22482 15762 22494
rect 20526 22482 20578 22494
rect 39790 22482 39842 22494
rect 14578 22430 14590 22482
rect 14642 22430 14654 22482
rect 19282 22430 19294 22482
rect 19346 22430 19358 22482
rect 25890 22430 25902 22482
rect 25954 22430 25966 22482
rect 30594 22430 30606 22482
rect 30658 22430 30670 22482
rect 13694 22418 13746 22430
rect 15710 22418 15762 22430
rect 20526 22418 20578 22430
rect 39790 22418 39842 22430
rect 41358 22482 41410 22494
rect 41358 22418 41410 22430
rect 4734 22370 4786 22382
rect 4274 22318 4286 22370
rect 4338 22318 4350 22370
rect 4734 22306 4786 22318
rect 5966 22370 6018 22382
rect 5966 22306 6018 22318
rect 6302 22370 6354 22382
rect 7870 22370 7922 22382
rect 12238 22370 12290 22382
rect 6850 22318 6862 22370
rect 6914 22318 6926 22370
rect 8418 22318 8430 22370
rect 8482 22318 8494 22370
rect 10434 22318 10446 22370
rect 10498 22318 10510 22370
rect 6302 22306 6354 22318
rect 7870 22306 7922 22318
rect 12238 22306 12290 22318
rect 15038 22370 15090 22382
rect 15822 22370 15874 22382
rect 19966 22370 20018 22382
rect 15362 22318 15374 22370
rect 15426 22318 15438 22370
rect 16370 22318 16382 22370
rect 16434 22318 16446 22370
rect 15038 22306 15090 22318
rect 15822 22306 15874 22318
rect 19966 22306 20018 22318
rect 21422 22370 21474 22382
rect 27022 22370 27074 22382
rect 21858 22318 21870 22370
rect 21922 22318 21934 22370
rect 22642 22318 22654 22370
rect 22706 22318 22718 22370
rect 23202 22318 23214 22370
rect 23266 22318 23278 22370
rect 24210 22318 24222 22370
rect 24274 22318 24286 22370
rect 26674 22318 26686 22370
rect 26738 22318 26750 22370
rect 21422 22306 21474 22318
rect 27022 22306 27074 22318
rect 27582 22370 27634 22382
rect 27582 22306 27634 22318
rect 29262 22370 29314 22382
rect 33518 22370 33570 22382
rect 42142 22370 42194 22382
rect 32274 22318 32286 22370
rect 32338 22318 32350 22370
rect 32610 22318 32622 22370
rect 32674 22318 32686 22370
rect 33394 22318 33406 22370
rect 33458 22318 33470 22370
rect 34290 22318 34302 22370
rect 34354 22318 34366 22370
rect 40226 22318 40238 22370
rect 40290 22318 40302 22370
rect 42466 22318 42478 22370
rect 42530 22318 42542 22370
rect 43474 22318 43486 22370
rect 43538 22318 43550 22370
rect 29262 22306 29314 22318
rect 33518 22306 33570 22318
rect 42142 22306 42194 22318
rect 5070 22258 5122 22270
rect 16046 22258 16098 22270
rect 26126 22258 26178 22270
rect 7074 22206 7086 22258
rect 7138 22206 7150 22258
rect 10546 22206 10558 22258
rect 10610 22206 10622 22258
rect 17154 22206 17166 22258
rect 17218 22206 17230 22258
rect 23426 22206 23438 22258
rect 23490 22206 23502 22258
rect 24322 22206 24334 22258
rect 24386 22206 24398 22258
rect 25330 22206 25342 22258
rect 25394 22206 25406 22258
rect 5070 22194 5122 22206
rect 16046 22194 16098 22206
rect 26126 22194 26178 22206
rect 27918 22258 27970 22270
rect 34526 22258 34578 22270
rect 31154 22206 31166 22258
rect 31218 22206 31230 22258
rect 35186 22206 35198 22258
rect 35250 22206 35262 22258
rect 37650 22206 37662 22258
rect 37714 22206 37726 22258
rect 38210 22206 38222 22258
rect 38274 22206 38286 22258
rect 27918 22194 27970 22206
rect 34526 22194 34578 22206
rect 7534 22146 7586 22158
rect 7534 22082 7586 22094
rect 8206 22146 8258 22158
rect 8206 22082 8258 22094
rect 11902 22146 11954 22158
rect 11902 22082 11954 22094
rect 13022 22146 13074 22158
rect 13022 22082 13074 22094
rect 13582 22146 13634 22158
rect 13582 22082 13634 22094
rect 15598 22146 15650 22158
rect 15598 22082 15650 22094
rect 21310 22146 21362 22158
rect 21310 22082 21362 22094
rect 21534 22146 21586 22158
rect 25006 22146 25058 22158
rect 23314 22094 23326 22146
rect 23378 22094 23390 22146
rect 21534 22082 21586 22094
rect 25006 22082 25058 22094
rect 25902 22146 25954 22158
rect 25902 22082 25954 22094
rect 27134 22146 27186 22158
rect 27134 22082 27186 22094
rect 27246 22146 27298 22158
rect 27246 22082 27298 22094
rect 28254 22146 28306 22158
rect 31278 22146 31330 22158
rect 28578 22094 28590 22146
rect 28642 22094 28654 22146
rect 28254 22082 28306 22094
rect 31278 22082 31330 22094
rect 34862 22146 34914 22158
rect 34862 22082 34914 22094
rect 35646 22146 35698 22158
rect 35646 22082 35698 22094
rect 40574 22146 40626 22158
rect 40574 22082 40626 22094
rect 1344 21978 46592 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 46592 21978
rect 1344 21892 46592 21926
rect 5630 21810 5682 21822
rect 4834 21758 4846 21810
rect 4898 21758 4910 21810
rect 5630 21746 5682 21758
rect 6302 21810 6354 21822
rect 6302 21746 6354 21758
rect 8094 21810 8146 21822
rect 8094 21746 8146 21758
rect 11566 21810 11618 21822
rect 11566 21746 11618 21758
rect 12238 21810 12290 21822
rect 12238 21746 12290 21758
rect 13806 21810 13858 21822
rect 13806 21746 13858 21758
rect 15038 21810 15090 21822
rect 15038 21746 15090 21758
rect 15150 21810 15202 21822
rect 15150 21746 15202 21758
rect 16046 21810 16098 21822
rect 16046 21746 16098 21758
rect 19966 21810 20018 21822
rect 19966 21746 20018 21758
rect 20414 21810 20466 21822
rect 20414 21746 20466 21758
rect 21982 21810 22034 21822
rect 21982 21746 22034 21758
rect 22094 21810 22146 21822
rect 22094 21746 22146 21758
rect 22318 21810 22370 21822
rect 22318 21746 22370 21758
rect 22654 21810 22706 21822
rect 22654 21746 22706 21758
rect 24334 21810 24386 21822
rect 24334 21746 24386 21758
rect 26126 21810 26178 21822
rect 26126 21746 26178 21758
rect 26238 21810 26290 21822
rect 26238 21746 26290 21758
rect 26798 21810 26850 21822
rect 26798 21746 26850 21758
rect 27806 21810 27858 21822
rect 27806 21746 27858 21758
rect 28478 21810 28530 21822
rect 36766 21810 36818 21822
rect 34738 21758 34750 21810
rect 34802 21758 34814 21810
rect 37986 21758 37998 21810
rect 38050 21758 38062 21810
rect 28478 21746 28530 21758
rect 36766 21746 36818 21758
rect 11902 21698 11954 21710
rect 6850 21646 6862 21698
rect 6914 21646 6926 21698
rect 7410 21646 7422 21698
rect 7474 21646 7486 21698
rect 11218 21646 11230 21698
rect 11282 21646 11294 21698
rect 11902 21634 11954 21646
rect 13134 21698 13186 21710
rect 13134 21634 13186 21646
rect 13470 21698 13522 21710
rect 13470 21634 13522 21646
rect 16830 21698 16882 21710
rect 16830 21634 16882 21646
rect 17614 21698 17666 21710
rect 17614 21634 17666 21646
rect 20526 21698 20578 21710
rect 28030 21698 28082 21710
rect 24658 21646 24670 21698
rect 24722 21646 24734 21698
rect 20526 21634 20578 21646
rect 28030 21634 28082 21646
rect 29262 21698 29314 21710
rect 35982 21698 36034 21710
rect 30258 21646 30270 21698
rect 30322 21646 30334 21698
rect 29262 21634 29314 21646
rect 35982 21634 36034 21646
rect 41134 21698 41186 21710
rect 41458 21646 41470 21698
rect 41522 21646 41534 21698
rect 45154 21646 45166 21698
rect 45218 21646 45230 21698
rect 41134 21634 41186 21646
rect 2158 21586 2210 21598
rect 10670 21586 10722 21598
rect 12574 21586 12626 21598
rect 2482 21534 2494 21586
rect 2546 21534 2558 21586
rect 10994 21534 11006 21586
rect 11058 21534 11070 21586
rect 2158 21522 2210 21534
rect 10670 21522 10722 21534
rect 12574 21522 12626 21534
rect 14814 21586 14866 21598
rect 14814 21522 14866 21534
rect 14926 21586 14978 21598
rect 15934 21586 15986 21598
rect 15362 21534 15374 21586
rect 15426 21534 15438 21586
rect 15698 21534 15710 21586
rect 15762 21534 15774 21586
rect 14926 21522 14978 21534
rect 15934 21522 15986 21534
rect 16158 21586 16210 21598
rect 17502 21586 17554 21598
rect 16370 21534 16382 21586
rect 16434 21534 16446 21586
rect 16158 21522 16210 21534
rect 17502 21522 17554 21534
rect 19406 21586 19458 21598
rect 19406 21522 19458 21534
rect 20302 21586 20354 21598
rect 20302 21522 20354 21534
rect 20974 21586 21026 21598
rect 20974 21522 21026 21534
rect 21870 21586 21922 21598
rect 27022 21586 27074 21598
rect 23090 21534 23102 21586
rect 23154 21534 23166 21586
rect 23426 21534 23438 21586
rect 23490 21534 23502 21586
rect 21870 21522 21922 21534
rect 27022 21522 27074 21534
rect 27246 21586 27298 21598
rect 30942 21586 30994 21598
rect 32958 21586 33010 21598
rect 35086 21586 35138 21598
rect 37662 21586 37714 21598
rect 29698 21534 29710 21586
rect 29762 21534 29774 21586
rect 30034 21534 30046 21586
rect 30098 21534 30110 21586
rect 31490 21534 31502 21586
rect 31554 21534 31566 21586
rect 32386 21534 32398 21586
rect 32450 21534 32462 21586
rect 33282 21534 33294 21586
rect 33346 21534 33358 21586
rect 33730 21534 33742 21586
rect 33794 21534 33806 21586
rect 36194 21534 36206 21586
rect 36258 21534 36270 21586
rect 42466 21534 42478 21586
rect 42530 21534 42542 21586
rect 43586 21534 43598 21586
rect 43650 21534 43662 21586
rect 44706 21534 44718 21586
rect 44770 21534 44782 21586
rect 27246 21522 27298 21534
rect 30942 21522 30994 21534
rect 32958 21522 33010 21534
rect 35086 21522 35138 21534
rect 37662 21522 37714 21534
rect 14366 21474 14418 21486
rect 14366 21410 14418 21422
rect 18062 21474 18114 21486
rect 27134 21474 27186 21486
rect 41918 21474 41970 21486
rect 23202 21422 23214 21474
rect 23266 21422 23278 21474
rect 27682 21422 27694 21474
rect 27746 21422 27758 21474
rect 28354 21422 28366 21474
rect 28418 21422 28430 21474
rect 35522 21422 35534 21474
rect 35586 21422 35598 21474
rect 18062 21410 18114 21422
rect 27134 21410 27186 21422
rect 41918 21410 41970 21422
rect 6638 21362 6690 21374
rect 6638 21298 6690 21310
rect 26350 21362 26402 21374
rect 26350 21298 26402 21310
rect 28702 21362 28754 21374
rect 43362 21310 43374 21362
rect 43426 21310 43438 21362
rect 28702 21298 28754 21310
rect 1344 21194 46592 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 46592 21194
rect 1344 21108 46592 21142
rect 13582 21026 13634 21038
rect 13582 20962 13634 20974
rect 22654 21026 22706 21038
rect 22654 20962 22706 20974
rect 27806 21026 27858 21038
rect 27806 20962 27858 20974
rect 33742 21026 33794 21038
rect 33742 20962 33794 20974
rect 11342 20914 11394 20926
rect 20302 20914 20354 20926
rect 2706 20862 2718 20914
rect 2770 20862 2782 20914
rect 10546 20862 10558 20914
rect 10610 20862 10622 20914
rect 13906 20862 13918 20914
rect 13970 20862 13982 20914
rect 11342 20850 11394 20862
rect 20302 20850 20354 20862
rect 27358 20914 27410 20926
rect 27358 20850 27410 20862
rect 28590 20914 28642 20926
rect 41134 20914 41186 20926
rect 29698 20862 29710 20914
rect 29762 20862 29774 20914
rect 35186 20862 35198 20914
rect 35250 20862 35262 20914
rect 28590 20850 28642 20862
rect 41134 20850 41186 20862
rect 6302 20802 6354 20814
rect 17166 20802 17218 20814
rect 4274 20750 4286 20802
rect 4338 20750 4350 20802
rect 6850 20750 6862 20802
rect 6914 20750 6926 20802
rect 7634 20750 7646 20802
rect 7698 20750 7710 20802
rect 12114 20750 12126 20802
rect 12178 20750 12190 20802
rect 16818 20750 16830 20802
rect 16882 20750 16894 20802
rect 6302 20738 6354 20750
rect 17166 20738 17218 20750
rect 17838 20802 17890 20814
rect 17838 20738 17890 20750
rect 20414 20802 20466 20814
rect 20414 20738 20466 20750
rect 20862 20802 20914 20814
rect 20862 20738 20914 20750
rect 22990 20802 23042 20814
rect 29262 20802 29314 20814
rect 33854 20802 33906 20814
rect 34526 20802 34578 20814
rect 27122 20750 27134 20802
rect 27186 20750 27198 20802
rect 27794 20750 27806 20802
rect 27858 20750 27870 20802
rect 30482 20750 30494 20802
rect 30546 20750 30558 20802
rect 30930 20750 30942 20802
rect 30994 20750 31006 20802
rect 32386 20750 32398 20802
rect 32450 20750 32462 20802
rect 33282 20750 33294 20802
rect 33346 20750 33358 20802
rect 34402 20750 34414 20802
rect 34466 20750 34478 20802
rect 22990 20738 23042 20750
rect 29262 20738 29314 20750
rect 33854 20738 33906 20750
rect 34526 20738 34578 20750
rect 34638 20802 34690 20814
rect 34638 20738 34690 20750
rect 35646 20802 35698 20814
rect 37986 20750 37998 20802
rect 38050 20750 38062 20802
rect 39106 20750 39118 20802
rect 39170 20750 39182 20802
rect 42690 20750 42702 20802
rect 42754 20750 42766 20802
rect 35646 20738 35698 20750
rect 13470 20690 13522 20702
rect 17278 20690 17330 20702
rect 27470 20690 27522 20702
rect 8418 20638 8430 20690
rect 8482 20638 8494 20690
rect 12002 20638 12014 20690
rect 12066 20638 12078 20690
rect 12898 20638 12910 20690
rect 12962 20638 12974 20690
rect 16034 20638 16046 20690
rect 16098 20638 16110 20690
rect 23202 20638 23214 20690
rect 23266 20638 23278 20690
rect 23762 20638 23774 20690
rect 23826 20638 23838 20690
rect 13470 20626 13522 20638
rect 17278 20626 17330 20638
rect 27470 20626 27522 20638
rect 28142 20690 28194 20702
rect 28142 20626 28194 20638
rect 30158 20690 30210 20702
rect 31614 20690 31666 20702
rect 31154 20638 31166 20690
rect 31218 20638 31230 20690
rect 30158 20626 30210 20638
rect 31614 20626 31666 20638
rect 34078 20690 34130 20702
rect 34078 20626 34130 20638
rect 35982 20690 36034 20702
rect 35982 20626 36034 20638
rect 36318 20690 36370 20702
rect 42142 20690 42194 20702
rect 36978 20638 36990 20690
rect 37042 20638 37054 20690
rect 39218 20638 39230 20690
rect 39282 20638 39294 20690
rect 36318 20626 36370 20638
rect 42142 20626 42194 20638
rect 5070 20578 5122 20590
rect 4722 20526 4734 20578
rect 4786 20526 4798 20578
rect 5070 20514 5122 20526
rect 5966 20578 6018 20590
rect 5966 20514 6018 20526
rect 6638 20578 6690 20590
rect 6638 20514 6690 20526
rect 11006 20578 11058 20590
rect 11006 20514 11058 20526
rect 12574 20578 12626 20590
rect 12574 20514 12626 20526
rect 17390 20578 17442 20590
rect 17390 20514 17442 20526
rect 20190 20578 20242 20590
rect 20190 20514 20242 20526
rect 24334 20578 24386 20590
rect 38098 20526 38110 20578
rect 38162 20526 38174 20578
rect 42466 20526 42478 20578
rect 42530 20526 42542 20578
rect 24334 20514 24386 20526
rect 1344 20410 46592 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 46592 20410
rect 1344 20324 46592 20358
rect 6078 20242 6130 20254
rect 6078 20178 6130 20190
rect 9550 20242 9602 20254
rect 24446 20242 24498 20254
rect 23090 20190 23102 20242
rect 23154 20190 23166 20242
rect 9550 20178 9602 20190
rect 24446 20178 24498 20190
rect 30830 20242 30882 20254
rect 30830 20178 30882 20190
rect 1710 20130 1762 20142
rect 5294 20130 5346 20142
rect 2034 20078 2046 20130
rect 2098 20078 2110 20130
rect 1710 20066 1762 20078
rect 5294 20066 5346 20078
rect 8542 20130 8594 20142
rect 8542 20066 8594 20078
rect 9886 20130 9938 20142
rect 22542 20130 22594 20142
rect 10658 20078 10670 20130
rect 10722 20078 10734 20130
rect 11666 20078 11678 20130
rect 11730 20078 11742 20130
rect 12002 20078 12014 20130
rect 12066 20078 12078 20130
rect 14018 20078 14030 20130
rect 14082 20078 14094 20130
rect 15250 20078 15262 20130
rect 15314 20078 15326 20130
rect 17378 20078 17390 20130
rect 17442 20078 17454 20130
rect 9886 20066 9938 20078
rect 22542 20066 22594 20078
rect 23774 20130 23826 20142
rect 33518 20130 33570 20142
rect 41806 20130 41858 20142
rect 43262 20130 43314 20142
rect 24098 20078 24110 20130
rect 24162 20078 24174 20130
rect 28690 20078 28702 20130
rect 28754 20078 28766 20130
rect 29586 20078 29598 20130
rect 29650 20078 29662 20130
rect 36082 20078 36094 20130
rect 36146 20078 36158 20130
rect 39890 20078 39902 20130
rect 39954 20078 39966 20130
rect 42802 20078 42814 20130
rect 42866 20078 42878 20130
rect 23774 20066 23826 20078
rect 33518 20066 33570 20078
rect 41806 20066 41858 20078
rect 43262 20066 43314 20078
rect 2382 20018 2434 20030
rect 6414 20018 6466 20030
rect 2930 19966 2942 20018
rect 2994 19966 3006 20018
rect 2382 19954 2434 19966
rect 6414 19954 6466 19966
rect 8878 20018 8930 20030
rect 11454 20018 11506 20030
rect 10434 19966 10446 20018
rect 10498 19966 10510 20018
rect 8878 19954 8930 19966
rect 11454 19954 11506 19966
rect 12798 20018 12850 20030
rect 18174 20018 18226 20030
rect 13458 19966 13470 20018
rect 13522 19966 13534 20018
rect 16706 19966 16718 20018
rect 16770 19966 16782 20018
rect 17602 19966 17614 20018
rect 17666 19966 17678 20018
rect 12798 19954 12850 19966
rect 18174 19954 18226 19966
rect 18622 20018 18674 20030
rect 18622 19954 18674 19966
rect 19854 20018 19906 20030
rect 19854 19954 19906 19966
rect 28366 20018 28418 20030
rect 31726 20018 31778 20030
rect 29250 19966 29262 20018
rect 29314 19966 29326 20018
rect 28366 19954 28418 19966
rect 31726 19954 31778 19966
rect 32510 20018 32562 20030
rect 32510 19954 32562 19966
rect 33182 20018 33234 20030
rect 33182 19954 33234 19966
rect 34526 20018 34578 20030
rect 34526 19954 34578 19966
rect 35086 20018 35138 20030
rect 36766 20018 36818 20030
rect 39230 20018 39282 20030
rect 35522 19966 35534 20018
rect 35586 19966 35598 20018
rect 35970 19966 35982 20018
rect 36034 19966 36046 20018
rect 37090 19966 37102 20018
rect 37154 19966 37166 20018
rect 38098 19966 38110 20018
rect 38162 19966 38174 20018
rect 35086 19954 35138 19966
rect 36766 19954 36818 19966
rect 39230 19954 39282 19966
rect 39566 20018 39618 20030
rect 41010 19966 41022 20018
rect 41074 19966 41086 20018
rect 42130 19966 42142 20018
rect 42194 19966 42206 20018
rect 42690 19966 42702 20018
rect 42754 19966 42766 20018
rect 44034 19966 44046 20018
rect 44098 19966 44110 20018
rect 44930 19966 44942 20018
rect 44994 19966 45006 20018
rect 39566 19954 39618 19966
rect 19630 19906 19682 19918
rect 13570 19854 13582 19906
rect 13634 19854 13646 19906
rect 19630 19842 19682 19854
rect 24558 19906 24610 19918
rect 40350 19906 40402 19918
rect 32050 19854 32062 19906
rect 32114 19854 32126 19906
rect 38770 19854 38782 19906
rect 38834 19854 38846 19906
rect 41346 19854 41358 19906
rect 41410 19854 41422 19906
rect 24558 19842 24610 19854
rect 40350 19842 40402 19854
rect 11118 19794 11170 19806
rect 11118 19730 11170 19742
rect 18062 19794 18114 19806
rect 18062 19730 18114 19742
rect 18510 19794 18562 19806
rect 33966 19794 34018 19806
rect 20290 19742 20302 19794
rect 20354 19742 20366 19794
rect 18510 19730 18562 19742
rect 33966 19730 34018 19742
rect 34190 19794 34242 19806
rect 34190 19730 34242 19742
rect 34638 19794 34690 19806
rect 34638 19730 34690 19742
rect 34750 19794 34802 19806
rect 34750 19730 34802 19742
rect 1344 19626 46592 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 46592 19626
rect 1344 19540 46592 19574
rect 4510 19458 4562 19470
rect 4510 19394 4562 19406
rect 10558 19458 10610 19470
rect 10558 19394 10610 19406
rect 10894 19458 10946 19470
rect 15698 19406 15710 19458
rect 15762 19406 15774 19458
rect 44034 19406 44046 19458
rect 44098 19406 44110 19458
rect 10894 19394 10946 19406
rect 3166 19346 3218 19358
rect 3166 19282 3218 19294
rect 4622 19346 4674 19358
rect 14478 19346 14530 19358
rect 21758 19346 21810 19358
rect 36990 19346 37042 19358
rect 7970 19294 7982 19346
rect 8034 19294 8046 19346
rect 10098 19294 10110 19346
rect 10162 19294 10174 19346
rect 15586 19294 15598 19346
rect 15650 19294 15662 19346
rect 20066 19294 20078 19346
rect 20130 19294 20142 19346
rect 33506 19294 33518 19346
rect 33570 19294 33582 19346
rect 4622 19282 4674 19294
rect 14478 19282 14530 19294
rect 21758 19282 21810 19294
rect 36990 19282 37042 19294
rect 2270 19234 2322 19246
rect 1810 19182 1822 19234
rect 1874 19182 1886 19234
rect 2270 19170 2322 19182
rect 3502 19234 3554 19246
rect 3502 19170 3554 19182
rect 5630 19234 5682 19246
rect 12350 19234 12402 19246
rect 7186 19182 7198 19234
rect 7250 19182 7262 19234
rect 11330 19182 11342 19234
rect 11394 19182 11406 19234
rect 5630 19170 5682 19182
rect 12350 19170 12402 19182
rect 13470 19234 13522 19246
rect 13470 19170 13522 19182
rect 14030 19234 14082 19246
rect 14030 19170 14082 19182
rect 15934 19234 15986 19246
rect 15934 19170 15986 19182
rect 16606 19234 16658 19246
rect 29374 19234 29426 19246
rect 17154 19182 17166 19234
rect 17218 19182 17230 19234
rect 23202 19182 23214 19234
rect 23266 19182 23278 19234
rect 16606 19170 16658 19182
rect 29374 19170 29426 19182
rect 32734 19234 32786 19246
rect 37886 19234 37938 19246
rect 35074 19182 35086 19234
rect 35138 19182 35150 19234
rect 35634 19182 35646 19234
rect 35698 19182 35710 19234
rect 36082 19182 36094 19234
rect 36146 19182 36158 19234
rect 37426 19182 37438 19234
rect 37490 19182 37502 19234
rect 32734 19170 32786 19182
rect 37886 19170 37938 19182
rect 38894 19234 38946 19246
rect 39330 19182 39342 19234
rect 39394 19182 39406 19234
rect 39778 19182 39790 19234
rect 39842 19182 39854 19234
rect 38894 19170 38946 19182
rect 2606 19122 2658 19134
rect 2606 19058 2658 19070
rect 5070 19122 5122 19134
rect 5070 19058 5122 19070
rect 6638 19122 6690 19134
rect 16270 19122 16322 19134
rect 11666 19070 11678 19122
rect 11730 19070 11742 19122
rect 6638 19058 6690 19070
rect 16270 19058 16322 19070
rect 16718 19122 16770 19134
rect 16718 19058 16770 19070
rect 16830 19122 16882 19134
rect 17938 19070 17950 19122
rect 18002 19070 18014 19122
rect 24546 19070 24558 19122
rect 24610 19070 24622 19122
rect 29698 19070 29710 19122
rect 29762 19070 29774 19122
rect 34514 19070 34526 19122
rect 34578 19070 34590 19122
rect 36418 19070 36430 19122
rect 36482 19070 36494 19122
rect 42578 19070 42590 19122
rect 42642 19070 42654 19122
rect 16830 19058 16882 19070
rect 4958 19010 5010 19022
rect 3826 18958 3838 19010
rect 3890 18958 3902 19010
rect 4958 18946 5010 18958
rect 6190 19010 6242 19022
rect 6190 18946 6242 18958
rect 12910 19010 12962 19022
rect 21646 19010 21698 19022
rect 13794 18958 13806 19010
rect 13858 18958 13870 19010
rect 12910 18946 12962 18958
rect 21646 18946 21698 18958
rect 32174 19010 32226 19022
rect 32174 18946 32226 18958
rect 33070 19010 33122 19022
rect 33070 18946 33122 18958
rect 34078 19010 34130 19022
rect 34078 18946 34130 18958
rect 36542 19010 36594 19022
rect 38670 19010 38722 19022
rect 38210 18958 38222 19010
rect 38274 18958 38286 19010
rect 36542 18946 36594 18958
rect 38670 18946 38722 18958
rect 1344 18842 46592 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 46592 18842
rect 1344 18756 46592 18790
rect 12798 18674 12850 18686
rect 12798 18610 12850 18622
rect 13022 18674 13074 18686
rect 13022 18610 13074 18622
rect 14030 18674 14082 18686
rect 14030 18610 14082 18622
rect 14254 18674 14306 18686
rect 14254 18610 14306 18622
rect 41582 18674 41634 18686
rect 41582 18610 41634 18622
rect 5630 18562 5682 18574
rect 5630 18498 5682 18510
rect 8318 18562 8370 18574
rect 8318 18498 8370 18510
rect 8990 18562 9042 18574
rect 8990 18498 9042 18510
rect 18398 18562 18450 18574
rect 18398 18498 18450 18510
rect 18510 18562 18562 18574
rect 29710 18562 29762 18574
rect 24546 18510 24558 18562
rect 24610 18510 24622 18562
rect 18510 18498 18562 18510
rect 29710 18498 29762 18510
rect 30382 18562 30434 18574
rect 30382 18498 30434 18510
rect 31950 18562 32002 18574
rect 31950 18498 32002 18510
rect 38894 18562 38946 18574
rect 38894 18498 38946 18510
rect 41358 18562 41410 18574
rect 41358 18498 41410 18510
rect 45054 18562 45106 18574
rect 45054 18498 45106 18510
rect 1710 18450 1762 18462
rect 1710 18386 1762 18398
rect 2942 18450 2994 18462
rect 14702 18450 14754 18462
rect 3378 18398 3390 18450
rect 3442 18398 3454 18450
rect 8082 18398 8094 18450
rect 8146 18398 8158 18450
rect 8754 18398 8766 18450
rect 8818 18398 8830 18450
rect 9538 18398 9550 18450
rect 9602 18398 9614 18450
rect 10322 18398 10334 18450
rect 10386 18398 10398 18450
rect 13346 18398 13358 18450
rect 13410 18398 13422 18450
rect 2942 18386 2994 18398
rect 14702 18386 14754 18398
rect 15486 18450 15538 18462
rect 16382 18450 16434 18462
rect 15922 18398 15934 18450
rect 15986 18398 15998 18450
rect 15486 18386 15538 18398
rect 16382 18386 16434 18398
rect 17390 18450 17442 18462
rect 17390 18386 17442 18398
rect 18174 18450 18226 18462
rect 18174 18386 18226 18398
rect 19182 18450 19234 18462
rect 19182 18386 19234 18398
rect 19742 18450 19794 18462
rect 22654 18450 22706 18462
rect 20514 18398 20526 18450
rect 20578 18398 20590 18450
rect 19742 18386 19794 18398
rect 22654 18386 22706 18398
rect 23438 18450 23490 18462
rect 39454 18450 39506 18462
rect 45950 18450 46002 18462
rect 24210 18398 24222 18450
rect 24274 18398 24286 18450
rect 29474 18398 29486 18450
rect 29538 18398 29550 18450
rect 30146 18398 30158 18450
rect 30210 18398 30222 18450
rect 34626 18398 34638 18450
rect 34690 18398 34702 18450
rect 35410 18398 35422 18450
rect 35474 18398 35486 18450
rect 36642 18398 36654 18450
rect 36706 18398 36718 18450
rect 38322 18398 38334 18450
rect 38386 18398 38398 18450
rect 42018 18398 42030 18450
rect 42082 18398 42094 18450
rect 42466 18398 42478 18450
rect 42530 18398 42542 18450
rect 23438 18386 23490 18398
rect 39454 18386 39506 18398
rect 45950 18386 46002 18398
rect 2270 18338 2322 18350
rect 12910 18338 12962 18350
rect 12450 18286 12462 18338
rect 12514 18286 12526 18338
rect 2270 18274 2322 18286
rect 12910 18274 12962 18286
rect 14142 18338 14194 18350
rect 16830 18338 16882 18350
rect 15026 18286 15038 18338
rect 15090 18286 15102 18338
rect 14142 18274 14194 18286
rect 16830 18274 16882 18286
rect 17950 18338 18002 18350
rect 25342 18338 25394 18350
rect 21746 18286 21758 18338
rect 21810 18286 21822 18338
rect 17950 18274 18002 18286
rect 25342 18274 25394 18286
rect 31726 18338 31778 18350
rect 31726 18274 31778 18286
rect 32510 18338 32562 18350
rect 34738 18286 34750 18338
rect 34802 18286 34814 18338
rect 35970 18286 35982 18338
rect 36034 18286 36046 18338
rect 37426 18286 37438 18338
rect 37490 18286 37502 18338
rect 32510 18274 32562 18286
rect 6414 18226 6466 18238
rect 6414 18162 6466 18174
rect 23774 18226 23826 18238
rect 23774 18162 23826 18174
rect 1344 18058 46592 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 46592 18058
rect 1344 17972 46592 18006
rect 4062 17890 4114 17902
rect 4062 17826 4114 17838
rect 4958 17890 5010 17902
rect 4958 17826 5010 17838
rect 10670 17890 10722 17902
rect 10670 17826 10722 17838
rect 11006 17890 11058 17902
rect 23762 17838 23774 17890
rect 23826 17838 23838 17890
rect 34402 17838 34414 17890
rect 34466 17838 34478 17890
rect 36306 17838 36318 17890
rect 36370 17887 36382 17890
rect 36530 17887 36542 17890
rect 36370 17841 36542 17887
rect 36370 17838 36382 17841
rect 36530 17838 36542 17841
rect 36594 17838 36606 17890
rect 42578 17838 42590 17890
rect 42642 17838 42654 17890
rect 11006 17826 11058 17838
rect 3278 17778 3330 17790
rect 3278 17714 3330 17726
rect 4174 17778 4226 17790
rect 4174 17714 4226 17726
rect 4622 17778 4674 17790
rect 4622 17714 4674 17726
rect 5070 17778 5122 17790
rect 5070 17714 5122 17726
rect 9662 17778 9714 17790
rect 17950 17778 18002 17790
rect 14802 17726 14814 17778
rect 14866 17726 14878 17778
rect 16930 17726 16942 17778
rect 16994 17726 17006 17778
rect 9662 17714 9714 17726
rect 17950 17714 18002 17726
rect 18622 17778 18674 17790
rect 18622 17714 18674 17726
rect 19854 17778 19906 17790
rect 29374 17778 29426 17790
rect 35870 17778 35922 17790
rect 37886 17778 37938 17790
rect 21970 17726 21982 17778
rect 22034 17726 22046 17778
rect 34962 17726 34974 17778
rect 35026 17726 35038 17778
rect 37426 17726 37438 17778
rect 37490 17726 37502 17778
rect 19854 17714 19906 17726
rect 29374 17714 29426 17726
rect 35870 17714 35922 17726
rect 37886 17714 37938 17726
rect 1710 17666 1762 17678
rect 1710 17602 1762 17614
rect 3502 17666 3554 17678
rect 3502 17602 3554 17614
rect 5518 17666 5570 17678
rect 12910 17666 12962 17678
rect 6066 17614 6078 17666
rect 6130 17614 6142 17666
rect 12450 17614 12462 17666
rect 12514 17614 12526 17666
rect 5518 17602 5570 17614
rect 12910 17602 12962 17614
rect 13358 17666 13410 17678
rect 13358 17602 13410 17614
rect 13694 17666 13746 17678
rect 18958 17666 19010 17678
rect 14018 17614 14030 17666
rect 14082 17614 14094 17666
rect 13694 17602 13746 17614
rect 18958 17602 19010 17614
rect 19518 17666 19570 17678
rect 19518 17602 19570 17614
rect 20414 17666 20466 17678
rect 20414 17602 20466 17614
rect 20638 17666 20690 17678
rect 20638 17602 20690 17614
rect 21422 17666 21474 17678
rect 21422 17602 21474 17614
rect 21646 17666 21698 17678
rect 35422 17666 35474 17678
rect 23202 17614 23214 17666
rect 23266 17614 23278 17666
rect 29810 17614 29822 17666
rect 29874 17614 29886 17666
rect 31266 17614 31278 17666
rect 31330 17614 31342 17666
rect 31714 17614 31726 17666
rect 31778 17614 31790 17666
rect 34066 17614 34078 17666
rect 34130 17614 34142 17666
rect 21646 17602 21698 17614
rect 35422 17602 35474 17614
rect 38446 17666 38498 17678
rect 38446 17602 38498 17614
rect 2382 17554 2434 17566
rect 2382 17490 2434 17502
rect 3614 17554 3666 17566
rect 3614 17490 3666 17502
rect 9214 17554 9266 17566
rect 9214 17490 9266 17502
rect 9886 17554 9938 17566
rect 9886 17490 9938 17502
rect 10222 17554 10274 17566
rect 13582 17554 13634 17566
rect 11330 17502 11342 17554
rect 11394 17502 11406 17554
rect 11554 17502 11566 17554
rect 11618 17502 11630 17554
rect 10222 17490 10274 17502
rect 13582 17490 13634 17502
rect 20078 17554 20130 17566
rect 20078 17490 20130 17502
rect 21982 17554 22034 17566
rect 21982 17490 22034 17502
rect 22206 17554 22258 17566
rect 28254 17554 28306 17566
rect 22866 17502 22878 17554
rect 22930 17502 22942 17554
rect 22206 17490 22258 17502
rect 28254 17490 28306 17502
rect 28590 17554 28642 17566
rect 28590 17490 28642 17502
rect 36430 17554 36482 17566
rect 36430 17490 36482 17502
rect 36990 17554 37042 17566
rect 39106 17502 39118 17554
rect 39170 17502 39182 17554
rect 36990 17490 37042 17502
rect 2046 17442 2098 17454
rect 2046 17378 2098 17390
rect 2718 17442 2770 17454
rect 17390 17442 17442 17454
rect 8418 17390 8430 17442
rect 8482 17390 8494 17442
rect 2718 17378 2770 17390
rect 17390 17378 17442 17390
rect 20750 17442 20802 17454
rect 20750 17378 20802 17390
rect 22542 17442 22594 17454
rect 22542 17378 22594 17390
rect 29598 17442 29650 17454
rect 29598 17378 29650 17390
rect 30942 17442 30994 17454
rect 30942 17378 30994 17390
rect 1344 17274 46592 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 46592 17274
rect 1344 17188 46592 17222
rect 5294 17106 5346 17118
rect 13022 17106 13074 17118
rect 4722 17054 4734 17106
rect 4786 17054 4798 17106
rect 8418 17054 8430 17106
rect 8482 17054 8494 17106
rect 12674 17054 12686 17106
rect 12738 17054 12750 17106
rect 5294 17042 5346 17054
rect 13022 17042 13074 17054
rect 18062 17106 18114 17118
rect 18062 17042 18114 17054
rect 23102 17106 23154 17118
rect 23102 17042 23154 17054
rect 23886 17106 23938 17118
rect 23886 17042 23938 17054
rect 24670 17106 24722 17118
rect 37550 17106 37602 17118
rect 35970 17054 35982 17106
rect 36034 17054 36046 17106
rect 24670 17042 24722 17054
rect 37550 17042 37602 17054
rect 38558 17106 38610 17118
rect 38558 17042 38610 17054
rect 40014 17106 40066 17118
rect 40014 17042 40066 17054
rect 9662 16994 9714 17006
rect 9662 16930 9714 16942
rect 9998 16994 10050 17006
rect 9998 16930 10050 16942
rect 10670 16994 10722 17006
rect 23326 16994 23378 17006
rect 39678 16994 39730 17006
rect 12114 16942 12126 16994
rect 12178 16942 12190 16994
rect 15698 16942 15710 16994
rect 15762 16942 15774 16994
rect 19618 16942 19630 16994
rect 19682 16942 19694 16994
rect 28466 16942 28478 16994
rect 28530 16942 28542 16994
rect 33282 16942 33294 16994
rect 33346 16942 33358 16994
rect 36306 16942 36318 16994
rect 36370 16942 36382 16994
rect 38882 16942 38894 16994
rect 38946 16942 38958 16994
rect 10670 16930 10722 16942
rect 23326 16930 23378 16942
rect 39678 16930 39730 16942
rect 5406 16882 5458 16894
rect 9102 16882 9154 16894
rect 17502 16882 17554 16894
rect 22766 16882 22818 16894
rect 1698 16830 1710 16882
rect 1762 16830 1774 16882
rect 2146 16830 2158 16882
rect 2210 16830 2222 16882
rect 5954 16830 5966 16882
rect 6018 16830 6030 16882
rect 10434 16830 10446 16882
rect 10498 16830 10510 16882
rect 12226 16830 12238 16882
rect 12290 16830 12302 16882
rect 16370 16830 16382 16882
rect 16434 16830 16446 16882
rect 21858 16830 21870 16882
rect 21922 16830 21934 16882
rect 5406 16818 5458 16830
rect 9102 16818 9154 16830
rect 17502 16818 17554 16830
rect 22766 16818 22818 16830
rect 26126 16882 26178 16894
rect 26126 16818 26178 16830
rect 26350 16882 26402 16894
rect 34750 16882 34802 16894
rect 39454 16882 39506 16894
rect 28354 16830 28366 16882
rect 28418 16830 28430 16882
rect 30258 16830 30270 16882
rect 30322 16830 30334 16882
rect 33170 16830 33182 16882
rect 33234 16830 33246 16882
rect 35746 16830 35758 16882
rect 35810 16830 35822 16882
rect 36530 16830 36542 16882
rect 36594 16830 36606 16882
rect 43474 16830 43486 16882
rect 43538 16830 43550 16882
rect 44370 16830 44382 16882
rect 44434 16830 44446 16882
rect 26350 16818 26402 16830
rect 34750 16818 34802 16830
rect 39454 16818 39506 16830
rect 11454 16770 11506 16782
rect 22990 16770 23042 16782
rect 13570 16718 13582 16770
rect 13634 16718 13646 16770
rect 18722 16718 18734 16770
rect 18786 16718 18798 16770
rect 11454 16706 11506 16718
rect 22990 16706 23042 16718
rect 23774 16770 23826 16782
rect 23774 16706 23826 16718
rect 26798 16770 26850 16782
rect 26798 16706 26850 16718
rect 27246 16770 27298 16782
rect 27246 16706 27298 16718
rect 32286 16770 32338 16782
rect 35186 16718 35198 16770
rect 35250 16718 35262 16770
rect 45490 16718 45502 16770
rect 45554 16718 45566 16770
rect 32286 16706 32338 16718
rect 11118 16658 11170 16670
rect 23662 16658 23714 16670
rect 21522 16606 21534 16658
rect 21586 16606 21598 16658
rect 11118 16594 11170 16606
rect 23662 16594 23714 16606
rect 25678 16658 25730 16670
rect 25678 16594 25730 16606
rect 25902 16658 25954 16670
rect 25902 16594 25954 16606
rect 26238 16658 26290 16670
rect 26238 16594 26290 16606
rect 26574 16658 26626 16670
rect 33966 16658 34018 16670
rect 31490 16606 31502 16658
rect 31554 16606 31566 16658
rect 26574 16594 26626 16606
rect 33966 16594 34018 16606
rect 34302 16658 34354 16670
rect 34302 16594 34354 16606
rect 1344 16490 46592 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 46592 16490
rect 1344 16404 46592 16438
rect 3502 16322 3554 16334
rect 3502 16258 3554 16270
rect 14366 16322 14418 16334
rect 20190 16322 20242 16334
rect 16594 16270 16606 16322
rect 16658 16270 16670 16322
rect 14366 16258 14418 16270
rect 20190 16258 20242 16270
rect 1822 16210 1874 16222
rect 1822 16146 1874 16158
rect 2270 16210 2322 16222
rect 2270 16146 2322 16158
rect 2718 16210 2770 16222
rect 2718 16146 2770 16158
rect 6078 16210 6130 16222
rect 11902 16210 11954 16222
rect 8978 16158 8990 16210
rect 9042 16158 9054 16210
rect 11106 16158 11118 16210
rect 11170 16158 11182 16210
rect 6078 16146 6130 16158
rect 11902 16146 11954 16158
rect 15262 16210 15314 16222
rect 30046 16210 30098 16222
rect 23650 16158 23662 16210
rect 23714 16158 23726 16210
rect 25442 16158 25454 16210
rect 25506 16158 25518 16210
rect 29250 16158 29262 16210
rect 29314 16158 29326 16210
rect 15262 16146 15314 16158
rect 30046 16146 30098 16158
rect 31726 16210 31778 16222
rect 35746 16158 35758 16210
rect 35810 16158 35822 16210
rect 38994 16158 39006 16210
rect 39058 16158 39070 16210
rect 31726 16146 31778 16158
rect 19966 16098 20018 16110
rect 25902 16098 25954 16110
rect 27358 16098 27410 16110
rect 8306 16046 8318 16098
rect 8370 16046 8382 16098
rect 12338 16046 12350 16098
rect 12402 16046 12414 16098
rect 13794 16046 13806 16098
rect 13858 16046 13870 16098
rect 16258 16046 16270 16098
rect 16322 16046 16334 16098
rect 19730 16046 19742 16098
rect 19794 16046 19806 16098
rect 20290 16046 20302 16098
rect 20354 16046 20366 16098
rect 21634 16046 21646 16098
rect 21698 16046 21710 16098
rect 24994 16046 25006 16098
rect 25058 16046 25070 16098
rect 26002 16046 26014 16098
rect 26066 16046 26078 16098
rect 26898 16046 26910 16098
rect 26962 16046 26974 16098
rect 19966 16034 20018 16046
rect 25902 16034 25954 16046
rect 27358 16034 27410 16046
rect 28030 16098 28082 16110
rect 28030 16034 28082 16046
rect 28590 16098 28642 16110
rect 28590 16034 28642 16046
rect 29710 16098 29762 16110
rect 29710 16034 29762 16046
rect 30606 16098 30658 16110
rect 30606 16034 30658 16046
rect 31278 16098 31330 16110
rect 38222 16098 38274 16110
rect 32162 16046 32174 16098
rect 32226 16046 32238 16098
rect 32498 16046 32510 16098
rect 32562 16046 32574 16098
rect 33730 16046 33742 16098
rect 33794 16046 33806 16098
rect 34850 16046 34862 16098
rect 34914 16046 34926 16098
rect 35410 16046 35422 16098
rect 35474 16046 35486 16098
rect 31278 16034 31330 16046
rect 38222 16034 38274 16046
rect 39454 16098 39506 16110
rect 41246 16098 41298 16110
rect 40114 16046 40126 16098
rect 40178 16046 40190 16098
rect 40674 16046 40686 16098
rect 40738 16046 40750 16098
rect 41906 16046 41918 16098
rect 41970 16046 41982 16098
rect 42914 16046 42926 16098
rect 42978 16046 42990 16098
rect 43586 16046 43598 16098
rect 43650 16046 43662 16098
rect 39454 16034 39506 16046
rect 41246 16034 41298 16046
rect 3614 15986 3666 15998
rect 15934 15986 15986 15998
rect 12674 15934 12686 15986
rect 12738 15934 12750 15986
rect 13570 15934 13582 15986
rect 13634 15934 13646 15986
rect 3614 15922 3666 15934
rect 15934 15922 15986 15934
rect 18622 15986 18674 15998
rect 33182 15986 33234 15998
rect 25330 15934 25342 15986
rect 25394 15934 25406 15986
rect 30930 15934 30942 15986
rect 30994 15934 31006 15986
rect 32722 15934 32734 15986
rect 32786 15934 32798 15986
rect 18622 15922 18674 15934
rect 33182 15922 33234 15934
rect 38558 15986 38610 15998
rect 38558 15922 38610 15934
rect 39790 15986 39842 15998
rect 43362 15934 43374 15986
rect 43426 15934 43438 15986
rect 39790 15922 39842 15934
rect 5966 15874 6018 15886
rect 5966 15810 6018 15822
rect 11566 15874 11618 15886
rect 11566 15810 11618 15822
rect 14702 15874 14754 15886
rect 14702 15810 14754 15822
rect 20526 15874 20578 15886
rect 20526 15810 20578 15822
rect 24334 15874 24386 15886
rect 40786 15822 40798 15874
rect 40850 15822 40862 15874
rect 24334 15810 24386 15822
rect 1344 15706 46592 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 46592 15706
rect 1344 15620 46592 15654
rect 9102 15538 9154 15550
rect 7970 15486 7982 15538
rect 8034 15486 8046 15538
rect 9102 15474 9154 15486
rect 11566 15538 11618 15550
rect 11566 15474 11618 15486
rect 12238 15538 12290 15550
rect 12238 15474 12290 15486
rect 13134 15538 13186 15550
rect 13134 15474 13186 15486
rect 16830 15538 16882 15550
rect 16830 15474 16882 15486
rect 20302 15538 20354 15550
rect 20302 15474 20354 15486
rect 21870 15538 21922 15550
rect 21870 15474 21922 15486
rect 22430 15538 22482 15550
rect 24110 15538 24162 15550
rect 23314 15486 23326 15538
rect 23378 15486 23390 15538
rect 22430 15474 22482 15486
rect 24110 15474 24162 15486
rect 25566 15538 25618 15550
rect 32398 15538 32450 15550
rect 37662 15538 37714 15550
rect 31042 15486 31054 15538
rect 31106 15486 31118 15538
rect 37314 15486 37326 15538
rect 37378 15486 37390 15538
rect 40002 15486 40014 15538
rect 40066 15486 40078 15538
rect 25566 15474 25618 15486
rect 32398 15474 32450 15486
rect 37662 15474 37714 15486
rect 4286 15426 4338 15438
rect 4286 15362 4338 15374
rect 4622 15426 4674 15438
rect 10558 15426 10610 15438
rect 9874 15374 9886 15426
rect 9938 15374 9950 15426
rect 4622 15362 4674 15374
rect 10558 15362 10610 15374
rect 10894 15426 10946 15438
rect 10894 15362 10946 15374
rect 11230 15426 11282 15438
rect 11230 15362 11282 15374
rect 14254 15426 14306 15438
rect 21646 15426 21698 15438
rect 33070 15426 33122 15438
rect 19506 15374 19518 15426
rect 19570 15374 19582 15426
rect 26002 15374 26014 15426
rect 26066 15374 26078 15426
rect 27682 15374 27694 15426
rect 27746 15374 27758 15426
rect 29922 15374 29934 15426
rect 29986 15374 29998 15426
rect 14254 15362 14306 15374
rect 21646 15362 21698 15374
rect 33070 15362 33122 15374
rect 33406 15426 33458 15438
rect 39678 15426 39730 15438
rect 35858 15374 35870 15426
rect 35922 15374 35934 15426
rect 38098 15374 38110 15426
rect 38162 15374 38174 15426
rect 33406 15362 33458 15374
rect 39678 15362 39730 15374
rect 5070 15314 5122 15326
rect 9550 15314 9602 15326
rect 12574 15314 12626 15326
rect 21310 15314 21362 15326
rect 23662 15314 23714 15326
rect 5506 15262 5518 15314
rect 5570 15262 5582 15314
rect 10322 15262 10334 15314
rect 10386 15262 10398 15314
rect 11778 15262 11790 15314
rect 11842 15262 11854 15314
rect 12898 15262 12910 15314
rect 12962 15262 12974 15314
rect 14018 15262 14030 15314
rect 14082 15262 14094 15314
rect 17490 15262 17502 15314
rect 17554 15262 17566 15314
rect 17714 15262 17726 15314
rect 17778 15262 17790 15314
rect 22642 15262 22654 15314
rect 22706 15262 22718 15314
rect 5070 15250 5122 15262
rect 9550 15250 9602 15262
rect 12574 15250 12626 15262
rect 21310 15250 21362 15262
rect 23662 15250 23714 15262
rect 25230 15314 25282 15326
rect 34414 15314 34466 15326
rect 25890 15262 25902 15314
rect 25954 15262 25966 15314
rect 27570 15262 27582 15314
rect 27634 15262 27646 15314
rect 30034 15262 30046 15314
rect 30098 15262 30110 15314
rect 30482 15262 30494 15314
rect 30546 15262 30558 15314
rect 34178 15262 34190 15314
rect 34242 15262 34254 15314
rect 35074 15262 35086 15314
rect 35138 15262 35150 15314
rect 35522 15262 35534 15314
rect 35586 15262 35598 15314
rect 40226 15262 40238 15314
rect 40290 15262 40302 15314
rect 41346 15262 41358 15314
rect 41410 15262 41422 15314
rect 42242 15262 42254 15314
rect 42306 15262 42318 15314
rect 25230 15250 25282 15262
rect 34414 15250 34466 15262
rect 3502 15202 3554 15214
rect 3502 15138 3554 15150
rect 3614 15202 3666 15214
rect 3614 15138 3666 15150
rect 8542 15202 8594 15214
rect 8542 15138 8594 15150
rect 13246 15202 13298 15214
rect 13246 15138 13298 15150
rect 20750 15202 20802 15214
rect 22318 15202 22370 15214
rect 21970 15150 21982 15202
rect 22034 15150 22046 15202
rect 20750 15138 20802 15150
rect 22318 15138 22370 15150
rect 24670 15202 24722 15214
rect 34850 15150 34862 15202
rect 34914 15150 34926 15202
rect 24670 15138 24722 15150
rect 45390 15090 45442 15102
rect 45390 15026 45442 15038
rect 1344 14922 46592 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 46592 14922
rect 1344 14836 46592 14870
rect 21310 14754 21362 14766
rect 21310 14690 21362 14702
rect 33854 14754 33906 14766
rect 33854 14690 33906 14702
rect 43038 14754 43090 14766
rect 43038 14690 43090 14702
rect 7310 14642 7362 14654
rect 23662 14642 23714 14654
rect 9762 14590 9774 14642
rect 9826 14590 9838 14642
rect 11890 14590 11902 14642
rect 11954 14590 11966 14642
rect 14690 14590 14702 14642
rect 14754 14590 14766 14642
rect 16818 14590 16830 14642
rect 16882 14590 16894 14642
rect 18610 14590 18622 14642
rect 18674 14590 18686 14642
rect 7310 14578 7362 14590
rect 23662 14578 23714 14590
rect 24110 14642 24162 14654
rect 24110 14578 24162 14590
rect 24670 14642 24722 14654
rect 24670 14578 24722 14590
rect 25006 14642 25058 14654
rect 25006 14578 25058 14590
rect 25342 14642 25394 14654
rect 25342 14578 25394 14590
rect 31726 14642 31778 14654
rect 31726 14578 31778 14590
rect 32622 14642 32674 14654
rect 32622 14578 32674 14590
rect 7982 14530 8034 14542
rect 19294 14530 19346 14542
rect 21422 14530 21474 14542
rect 29374 14530 29426 14542
rect 4834 14478 4846 14530
rect 4898 14478 4910 14530
rect 12562 14478 12574 14530
rect 12626 14478 12638 14530
rect 13906 14478 13918 14530
rect 13970 14478 13982 14530
rect 19730 14478 19742 14530
rect 19794 14478 19806 14530
rect 20514 14478 20526 14530
rect 20578 14478 20590 14530
rect 21634 14478 21646 14530
rect 21698 14478 21710 14530
rect 25778 14478 25790 14530
rect 25842 14478 25854 14530
rect 26114 14478 26126 14530
rect 26178 14478 26190 14530
rect 27570 14478 27582 14530
rect 27634 14478 27646 14530
rect 28466 14478 28478 14530
rect 28530 14478 28542 14530
rect 29138 14478 29150 14530
rect 29202 14478 29214 14530
rect 7982 14466 8034 14478
rect 19294 14466 19346 14478
rect 21422 14466 21474 14478
rect 29374 14466 29426 14478
rect 29486 14530 29538 14542
rect 29486 14466 29538 14478
rect 29598 14530 29650 14542
rect 30158 14530 30210 14542
rect 29810 14478 29822 14530
rect 29874 14478 29886 14530
rect 29598 14466 29650 14478
rect 30158 14466 30210 14478
rect 30830 14530 30882 14542
rect 30830 14466 30882 14478
rect 32062 14530 32114 14542
rect 34190 14530 34242 14542
rect 35534 14530 35586 14542
rect 33170 14478 33182 14530
rect 33234 14478 33246 14530
rect 34850 14478 34862 14530
rect 34914 14478 34926 14530
rect 32062 14466 32114 14478
rect 34190 14466 34242 14478
rect 35534 14466 35586 14478
rect 38670 14530 38722 14542
rect 38994 14478 39006 14530
rect 39058 14478 39070 14530
rect 39330 14478 39342 14530
rect 39394 14478 39406 14530
rect 38670 14466 38722 14478
rect 8318 14418 8370 14430
rect 26798 14418 26850 14430
rect 26338 14366 26350 14418
rect 26402 14366 26414 14418
rect 8318 14354 8370 14366
rect 26798 14354 26850 14366
rect 32958 14418 33010 14430
rect 36990 14418 37042 14430
rect 34962 14366 34974 14418
rect 35026 14366 35038 14418
rect 32958 14354 33010 14366
rect 36990 14354 37042 14366
rect 37774 14418 37826 14430
rect 37774 14354 37826 14366
rect 7198 14306 7250 14318
rect 4610 14254 4622 14306
rect 4674 14254 4686 14306
rect 7198 14242 7250 14254
rect 18174 14306 18226 14318
rect 18174 14242 18226 14254
rect 19966 14306 20018 14318
rect 19966 14242 20018 14254
rect 20302 14306 20354 14318
rect 20302 14242 20354 14254
rect 30494 14306 30546 14318
rect 30494 14242 30546 14254
rect 31166 14306 31218 14318
rect 31166 14242 31218 14254
rect 37326 14306 37378 14318
rect 37326 14242 37378 14254
rect 38110 14306 38162 14318
rect 38110 14242 38162 14254
rect 38446 14306 38498 14318
rect 42354 14254 42366 14306
rect 42418 14254 42430 14306
rect 38446 14242 38498 14254
rect 1344 14138 46592 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 46592 14138
rect 1344 14052 46592 14086
rect 5294 13970 5346 13982
rect 18734 13970 18786 13982
rect 4498 13918 4510 13970
rect 4562 13918 4574 13970
rect 8306 13918 8318 13970
rect 8370 13918 8382 13970
rect 5294 13906 5346 13918
rect 18734 13906 18786 13918
rect 24110 13970 24162 13982
rect 24110 13906 24162 13918
rect 25454 13970 25506 13982
rect 25454 13906 25506 13918
rect 27806 13970 27858 13982
rect 27806 13906 27858 13918
rect 29038 13970 29090 13982
rect 29038 13906 29090 13918
rect 29598 13970 29650 13982
rect 29598 13906 29650 13918
rect 34974 13970 35026 13982
rect 34974 13906 35026 13918
rect 38782 13970 38834 13982
rect 38782 13906 38834 13918
rect 40910 13970 40962 13982
rect 40910 13906 40962 13918
rect 14142 13858 14194 13870
rect 11106 13806 11118 13858
rect 11170 13806 11182 13858
rect 14142 13794 14194 13806
rect 15150 13858 15202 13870
rect 15150 13794 15202 13806
rect 15822 13858 15874 13870
rect 25678 13858 25730 13870
rect 17938 13806 17950 13858
rect 18002 13806 18014 13858
rect 22306 13806 22318 13858
rect 22370 13806 22382 13858
rect 15822 13794 15874 13806
rect 25678 13794 25730 13806
rect 26014 13858 26066 13870
rect 27470 13858 27522 13870
rect 33966 13858 34018 13870
rect 26338 13806 26350 13858
rect 26402 13806 26414 13858
rect 28466 13806 28478 13858
rect 28530 13806 28542 13858
rect 32050 13806 32062 13858
rect 32114 13806 32126 13858
rect 35410 13806 35422 13858
rect 35474 13806 35486 13858
rect 37986 13806 37998 13858
rect 38050 13806 38062 13858
rect 39330 13806 39342 13858
rect 39394 13806 39406 13858
rect 39890 13806 39902 13858
rect 39954 13806 39966 13858
rect 45266 13806 45278 13858
rect 45330 13806 45342 13858
rect 26014 13794 26066 13806
rect 27470 13794 27522 13806
rect 33966 13794 34018 13806
rect 1822 13746 1874 13758
rect 5630 13746 5682 13758
rect 14478 13746 14530 13758
rect 2146 13694 2158 13746
rect 2210 13694 2222 13746
rect 6066 13694 6078 13746
rect 6130 13694 6142 13746
rect 10322 13694 10334 13746
rect 10386 13694 10398 13746
rect 1822 13682 1874 13694
rect 5630 13682 5682 13694
rect 14478 13682 14530 13694
rect 14814 13746 14866 13758
rect 14814 13682 14866 13694
rect 15486 13746 15538 13758
rect 15486 13682 15538 13694
rect 18286 13746 18338 13758
rect 26686 13746 26738 13758
rect 19618 13694 19630 13746
rect 19682 13694 19694 13746
rect 18286 13682 18338 13694
rect 26686 13682 26738 13694
rect 28142 13746 28194 13758
rect 28142 13682 28194 13694
rect 29262 13746 29314 13758
rect 29262 13682 29314 13694
rect 30494 13746 30546 13758
rect 33630 13746 33682 13758
rect 31602 13694 31614 13746
rect 31666 13694 31678 13746
rect 32274 13694 32286 13746
rect 32338 13694 32350 13746
rect 34402 13694 34414 13746
rect 34466 13694 34478 13746
rect 35298 13694 35310 13746
rect 35362 13694 35374 13746
rect 37650 13694 37662 13746
rect 37714 13694 37726 13746
rect 38210 13694 38222 13746
rect 38274 13694 38286 13746
rect 41122 13694 41134 13746
rect 41186 13694 41198 13746
rect 42690 13694 42702 13746
rect 42754 13694 42766 13746
rect 43698 13694 43710 13746
rect 43762 13694 43774 13746
rect 30494 13682 30546 13694
rect 33630 13682 33682 13694
rect 17614 13634 17666 13646
rect 13234 13582 13246 13634
rect 13298 13582 13310 13634
rect 17614 13570 17666 13582
rect 29934 13634 29986 13646
rect 33070 13634 33122 13646
rect 31266 13582 31278 13634
rect 31330 13582 31342 13634
rect 36306 13582 36318 13634
rect 36370 13582 36382 13634
rect 29934 13570 29986 13582
rect 33070 13570 33122 13582
rect 9102 13522 9154 13534
rect 9102 13458 9154 13470
rect 39118 13522 39170 13534
rect 39118 13458 39170 13470
rect 1344 13354 46592 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 46592 13354
rect 1344 13268 46592 13302
rect 16942 13186 16994 13198
rect 32286 13186 32338 13198
rect 30034 13134 30046 13186
rect 30098 13134 30110 13186
rect 16942 13122 16994 13134
rect 32286 13122 32338 13134
rect 8654 13074 8706 13086
rect 8654 13010 8706 13022
rect 18174 13074 18226 13086
rect 18174 13010 18226 13022
rect 37326 13074 37378 13086
rect 37986 13022 37998 13074
rect 38050 13022 38062 13074
rect 37326 13010 37378 13022
rect 13694 12962 13746 12974
rect 13694 12898 13746 12910
rect 14254 12962 14306 12974
rect 14254 12898 14306 12910
rect 14590 12962 14642 12974
rect 14590 12898 14642 12910
rect 15262 12962 15314 12974
rect 15262 12898 15314 12910
rect 15822 12962 15874 12974
rect 19070 12962 19122 12974
rect 20414 12962 20466 12974
rect 17714 12910 17726 12962
rect 17778 12910 17790 12962
rect 19842 12910 19854 12962
rect 19906 12910 19918 12962
rect 15822 12898 15874 12910
rect 19070 12898 19122 12910
rect 20414 12898 20466 12910
rect 23886 12962 23938 12974
rect 23886 12898 23938 12910
rect 24446 12962 24498 12974
rect 30382 12962 30434 12974
rect 31390 12962 31442 12974
rect 26450 12910 26462 12962
rect 26514 12910 26526 12962
rect 26898 12910 26910 12962
rect 26962 12910 26974 12962
rect 27570 12910 27582 12962
rect 27634 12910 27646 12962
rect 29810 12910 29822 12962
rect 29874 12910 29886 12962
rect 30258 12910 30270 12962
rect 30322 12910 30334 12962
rect 31042 12910 31054 12962
rect 31106 12910 31118 12962
rect 24446 12898 24498 12910
rect 30382 12898 30434 12910
rect 31390 12898 31442 12910
rect 32510 12962 32562 12974
rect 32510 12898 32562 12910
rect 32734 12962 32786 12974
rect 34862 12962 34914 12974
rect 37550 12962 37602 12974
rect 33618 12910 33630 12962
rect 33682 12910 33694 12962
rect 33954 12910 33966 12962
rect 34018 12910 34030 12962
rect 35410 12910 35422 12962
rect 35474 12910 35486 12962
rect 36306 12910 36318 12962
rect 36370 12910 36382 12962
rect 40226 12910 40238 12962
rect 40290 12910 40302 12962
rect 40674 12910 40686 12962
rect 40738 12910 40750 12962
rect 42130 12910 42142 12962
rect 42194 12910 42206 12962
rect 43026 12910 43038 12962
rect 43090 12910 43102 12962
rect 32734 12898 32786 12910
rect 34862 12898 34914 12910
rect 37550 12898 37602 12910
rect 3614 12850 3666 12862
rect 13918 12850 13970 12862
rect 12898 12798 12910 12850
rect 12962 12798 12974 12850
rect 3614 12786 3666 12798
rect 13918 12786 13970 12798
rect 14926 12850 14978 12862
rect 14926 12786 14978 12798
rect 16718 12850 16770 12862
rect 16718 12786 16770 12798
rect 18510 12850 18562 12862
rect 18510 12786 18562 12798
rect 19406 12850 19458 12862
rect 19406 12786 19458 12798
rect 23326 12850 23378 12862
rect 31838 12850 31890 12862
rect 33182 12850 33234 12862
rect 38670 12850 38722 12862
rect 25554 12798 25566 12850
rect 25618 12798 25630 12850
rect 27794 12798 27806 12850
rect 27858 12798 27870 12850
rect 32050 12798 32062 12850
rect 32114 12798 32126 12850
rect 34178 12798 34190 12850
rect 34242 12798 34254 12850
rect 23326 12786 23378 12798
rect 31838 12786 31890 12798
rect 33182 12786 33234 12798
rect 38670 12786 38722 12798
rect 39678 12850 39730 12862
rect 39678 12786 39730 12798
rect 39902 12850 39954 12862
rect 41358 12850 41410 12862
rect 40898 12798 40910 12850
rect 40962 12798 40974 12850
rect 39902 12786 39954 12798
rect 41358 12786 41410 12798
rect 3502 12738 3554 12750
rect 3502 12674 3554 12686
rect 8542 12738 8594 12750
rect 8542 12674 8594 12686
rect 12574 12738 12626 12750
rect 24558 12738 24610 12750
rect 17266 12686 17278 12738
rect 17330 12686 17342 12738
rect 12574 12674 12626 12686
rect 24558 12674 24610 12686
rect 24782 12738 24834 12750
rect 24782 12674 24834 12686
rect 25230 12738 25282 12750
rect 27458 12686 27470 12738
rect 27522 12686 27534 12738
rect 32162 12686 32174 12738
rect 32226 12686 32238 12738
rect 25230 12674 25282 12686
rect 1344 12570 46592 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 46592 12570
rect 1344 12484 46592 12518
rect 5294 12402 5346 12414
rect 4722 12350 4734 12402
rect 4786 12350 4798 12402
rect 5294 12338 5346 12350
rect 11790 12402 11842 12414
rect 11790 12338 11842 12350
rect 12014 12402 12066 12414
rect 12014 12338 12066 12350
rect 12686 12402 12738 12414
rect 12686 12338 12738 12350
rect 18174 12402 18226 12414
rect 18174 12338 18226 12350
rect 20302 12402 20354 12414
rect 20302 12338 20354 12350
rect 21534 12402 21586 12414
rect 21534 12338 21586 12350
rect 22206 12402 22258 12414
rect 41134 12402 41186 12414
rect 26226 12350 26238 12402
rect 26290 12350 26302 12402
rect 30258 12350 30270 12402
rect 30322 12350 30334 12402
rect 35746 12350 35758 12402
rect 35810 12350 35822 12402
rect 40226 12350 40238 12402
rect 40290 12350 40302 12402
rect 22206 12338 22258 12350
rect 41134 12338 41186 12350
rect 41806 12402 41858 12414
rect 41806 12338 41858 12350
rect 45838 12402 45890 12414
rect 45838 12338 45890 12350
rect 6190 12290 6242 12302
rect 13022 12290 13074 12302
rect 21086 12290 21138 12302
rect 12338 12238 12350 12290
rect 12402 12238 12414 12290
rect 19282 12238 19294 12290
rect 19346 12238 19358 12290
rect 19730 12238 19742 12290
rect 19794 12238 19806 12290
rect 6190 12226 6242 12238
rect 13022 12226 13074 12238
rect 21086 12226 21138 12238
rect 22542 12290 22594 12302
rect 22542 12226 22594 12238
rect 22878 12290 22930 12302
rect 23202 12238 23214 12290
rect 23266 12238 23278 12290
rect 33730 12238 33742 12290
rect 33794 12238 33806 12290
rect 35634 12238 35646 12290
rect 35698 12238 35710 12290
rect 36530 12238 36542 12290
rect 36594 12238 36606 12290
rect 37650 12238 37662 12290
rect 37714 12238 37726 12290
rect 22878 12226 22930 12238
rect 1822 12178 1874 12190
rect 8878 12178 8930 12190
rect 17838 12178 17890 12190
rect 2146 12126 2158 12178
rect 2210 12126 2222 12178
rect 8418 12126 8430 12178
rect 8482 12126 8494 12178
rect 13458 12126 13470 12178
rect 13522 12126 13534 12178
rect 16482 12126 16494 12178
rect 16546 12126 16558 12178
rect 1822 12114 1874 12126
rect 8878 12114 8930 12126
rect 17838 12114 17890 12126
rect 17950 12178 18002 12190
rect 17950 12114 18002 12126
rect 18398 12178 18450 12190
rect 18398 12114 18450 12126
rect 20750 12178 20802 12190
rect 30942 12178 30994 12190
rect 42030 12178 42082 12190
rect 23426 12126 23438 12178
rect 23490 12126 23502 12178
rect 24322 12126 24334 12178
rect 24386 12126 24398 12178
rect 25554 12126 25566 12178
rect 25618 12126 25630 12178
rect 26114 12126 26126 12178
rect 26178 12126 26190 12178
rect 26786 12126 26798 12178
rect 26850 12126 26862 12178
rect 27458 12126 27470 12178
rect 27522 12126 27534 12178
rect 28242 12126 28254 12178
rect 28306 12126 28318 12178
rect 29586 12126 29598 12178
rect 29650 12126 29662 12178
rect 30034 12126 30046 12178
rect 30098 12126 30110 12178
rect 31490 12126 31502 12178
rect 31554 12126 31566 12178
rect 32386 12126 32398 12178
rect 32450 12126 32462 12178
rect 33058 12126 33070 12178
rect 33122 12126 33134 12178
rect 33618 12126 33630 12178
rect 33682 12126 33694 12178
rect 34962 12126 34974 12178
rect 35026 12126 35038 12178
rect 35522 12126 35534 12178
rect 35586 12126 35598 12178
rect 36642 12126 36654 12178
rect 36706 12126 36718 12178
rect 42354 12126 42366 12178
rect 42418 12126 42430 12178
rect 42802 12126 42814 12178
rect 42866 12126 42878 12178
rect 20750 12114 20802 12126
rect 30942 12114 30994 12126
rect 42030 12114 42082 12126
rect 9662 12066 9714 12078
rect 9662 12002 9714 12014
rect 10110 12066 10162 12078
rect 10110 12002 10162 12014
rect 13918 12066 13970 12078
rect 23886 12066 23938 12078
rect 15362 12014 15374 12066
rect 15426 12014 15438 12066
rect 13918 12002 13970 12014
rect 23886 12002 23938 12014
rect 25230 12066 25282 12078
rect 25230 12002 25282 12014
rect 29262 12066 29314 12078
rect 34066 12014 34078 12066
rect 34130 12014 34142 12066
rect 29262 12002 29314 12014
rect 5406 11954 5458 11966
rect 5406 11890 5458 11902
rect 9550 11954 9602 11966
rect 9550 11890 9602 11902
rect 9998 11954 10050 11966
rect 9998 11890 10050 11902
rect 18286 11954 18338 11966
rect 18286 11890 18338 11902
rect 19966 11954 20018 11966
rect 19966 11890 20018 11902
rect 1344 11786 46592 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 46592 11786
rect 1344 11700 46592 11734
rect 4062 11618 4114 11630
rect 4062 11554 4114 11566
rect 11006 11618 11058 11630
rect 11006 11554 11058 11566
rect 42478 11618 42530 11630
rect 42478 11554 42530 11566
rect 3726 11506 3778 11518
rect 3726 11442 3778 11454
rect 6190 11506 6242 11518
rect 6190 11442 6242 11454
rect 19854 11506 19906 11518
rect 19854 11442 19906 11454
rect 26126 11506 26178 11518
rect 30606 11506 30658 11518
rect 29586 11454 29598 11506
rect 29650 11454 29662 11506
rect 32162 11454 32174 11506
rect 32226 11454 32238 11506
rect 33954 11454 33966 11506
rect 34018 11454 34030 11506
rect 34626 11454 34638 11506
rect 34690 11454 34702 11506
rect 26126 11442 26178 11454
rect 30606 11442 30658 11454
rect 3614 11394 3666 11406
rect 3614 11330 3666 11342
rect 5630 11394 5682 11406
rect 5630 11330 5682 11342
rect 7310 11394 7362 11406
rect 19630 11394 19682 11406
rect 23102 11394 23154 11406
rect 7970 11342 7982 11394
rect 8034 11342 8046 11394
rect 11330 11342 11342 11394
rect 11394 11342 11406 11394
rect 12002 11342 12014 11394
rect 12066 11342 12078 11394
rect 12674 11342 12686 11394
rect 12738 11342 12750 11394
rect 14690 11342 14702 11394
rect 14754 11342 14766 11394
rect 15026 11342 15038 11394
rect 15090 11342 15102 11394
rect 16370 11342 16382 11394
rect 16434 11342 16446 11394
rect 16818 11342 16830 11394
rect 16882 11342 16894 11394
rect 18050 11342 18062 11394
rect 18114 11342 18126 11394
rect 19170 11342 19182 11394
rect 19234 11342 19246 11394
rect 20066 11342 20078 11394
rect 20130 11342 20142 11394
rect 21298 11342 21310 11394
rect 21362 11342 21374 11394
rect 22642 11342 22654 11394
rect 22706 11342 22718 11394
rect 7310 11330 7362 11342
rect 19630 11330 19682 11342
rect 23102 11330 23154 11342
rect 23886 11394 23938 11406
rect 23886 11330 23938 11342
rect 24222 11394 24274 11406
rect 24222 11330 24274 11342
rect 26014 11394 26066 11406
rect 37774 11394 37826 11406
rect 26338 11342 26350 11394
rect 26402 11342 26414 11394
rect 27794 11342 27806 11394
rect 27858 11342 27870 11394
rect 30146 11342 30158 11394
rect 30210 11342 30222 11394
rect 31714 11342 31726 11394
rect 31778 11342 31790 11394
rect 33506 11342 33518 11394
rect 33570 11342 33582 11394
rect 34514 11342 34526 11394
rect 34578 11342 34590 11394
rect 37202 11342 37214 11394
rect 37266 11342 37278 11394
rect 26014 11330 26066 11342
rect 37774 11330 37826 11342
rect 37998 11394 38050 11406
rect 38322 11342 38334 11394
rect 38386 11342 38398 11394
rect 38658 11342 38670 11394
rect 38722 11342 38734 11394
rect 37998 11330 38050 11342
rect 4174 11282 4226 11294
rect 12910 11282 12962 11294
rect 16046 11282 16098 11294
rect 17502 11282 17554 11294
rect 11554 11230 11566 11282
rect 11618 11230 11630 11282
rect 15698 11230 15710 11282
rect 15762 11230 15774 11282
rect 17042 11230 17054 11282
rect 17106 11230 17118 11282
rect 4174 11218 4226 11230
rect 12910 11218 12962 11230
rect 16046 11218 16098 11230
rect 17502 11218 17554 11230
rect 27358 11282 27410 11294
rect 36978 11230 36990 11282
rect 37042 11230 37054 11282
rect 41570 11230 41582 11282
rect 41634 11230 41646 11282
rect 27358 11218 27410 11230
rect 12238 11170 12290 11182
rect 10322 11118 10334 11170
rect 10386 11118 10398 11170
rect 12238 11106 12290 11118
rect 21422 11170 21474 11182
rect 21422 11106 21474 11118
rect 29150 11170 29202 11182
rect 29150 11106 29202 11118
rect 1344 11002 46592 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 46592 11002
rect 1344 10916 46592 10950
rect 5294 10834 5346 10846
rect 23662 10834 23714 10846
rect 4722 10782 4734 10834
rect 4786 10782 4798 10834
rect 6066 10782 6078 10834
rect 6130 10782 6142 10834
rect 12450 10782 12462 10834
rect 12514 10782 12526 10834
rect 19506 10782 19518 10834
rect 19570 10782 19582 10834
rect 5294 10770 5346 10782
rect 23662 10770 23714 10782
rect 24446 10834 24498 10846
rect 24446 10770 24498 10782
rect 24558 10834 24610 10846
rect 24558 10770 24610 10782
rect 24670 10834 24722 10846
rect 24670 10770 24722 10782
rect 33182 10834 33234 10846
rect 33182 10770 33234 10782
rect 33294 10834 33346 10846
rect 33294 10770 33346 10782
rect 33406 10834 33458 10846
rect 33406 10770 33458 10782
rect 14814 10722 14866 10734
rect 26238 10722 26290 10734
rect 22530 10670 22542 10722
rect 22594 10670 22606 10722
rect 23090 10670 23102 10722
rect 23154 10670 23166 10722
rect 28242 10670 28254 10722
rect 28306 10670 28318 10722
rect 14814 10658 14866 10670
rect 26238 10658 26290 10670
rect 1822 10610 1874 10622
rect 9102 10610 9154 10622
rect 2146 10558 2158 10610
rect 2210 10558 2222 10610
rect 8418 10558 8430 10610
rect 8482 10558 8494 10610
rect 1822 10546 1874 10558
rect 9102 10546 9154 10558
rect 9662 10610 9714 10622
rect 13918 10610 13970 10622
rect 9986 10558 9998 10610
rect 10050 10558 10062 10610
rect 13458 10558 13470 10610
rect 13522 10558 13534 10610
rect 9662 10546 9714 10558
rect 13918 10546 13970 10558
rect 14366 10610 14418 10622
rect 14366 10546 14418 10558
rect 16046 10610 16098 10622
rect 17614 10610 17666 10622
rect 17378 10558 17390 10610
rect 17442 10558 17454 10610
rect 16046 10546 16098 10558
rect 17614 10546 17666 10558
rect 17726 10610 17778 10622
rect 19966 10610 20018 10622
rect 23998 10610 24050 10622
rect 18946 10558 18958 10610
rect 19010 10558 19022 10610
rect 19282 10558 19294 10610
rect 19346 10558 19358 10610
rect 20738 10558 20750 10610
rect 20802 10558 20814 10610
rect 21634 10558 21646 10610
rect 21698 10558 21710 10610
rect 27010 10558 27022 10610
rect 27074 10558 27086 10610
rect 29922 10558 29934 10610
rect 29986 10558 29998 10610
rect 30370 10558 30382 10610
rect 30434 10558 30446 10610
rect 31490 10558 31502 10610
rect 31554 10558 31566 10610
rect 17726 10546 17778 10558
rect 19966 10546 20018 10558
rect 23998 10546 24050 10558
rect 16606 10498 16658 10510
rect 18510 10498 18562 10510
rect 33630 10498 33682 10510
rect 18162 10446 18174 10498
rect 18226 10446 18238 10498
rect 25666 10446 25678 10498
rect 25730 10446 25742 10498
rect 29586 10446 29598 10498
rect 29650 10446 29662 10498
rect 16606 10434 16658 10446
rect 18510 10434 18562 10446
rect 33630 10434 33682 10446
rect 33854 10498 33906 10510
rect 33854 10434 33906 10446
rect 5406 10386 5458 10398
rect 5406 10322 5458 10334
rect 13134 10386 13186 10398
rect 13134 10322 13186 10334
rect 23326 10386 23378 10398
rect 23326 10322 23378 10334
rect 1344 10218 46592 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 46592 10218
rect 1344 10132 46592 10166
rect 6078 10050 6130 10062
rect 6078 9986 6130 9998
rect 11454 10050 11506 10062
rect 11454 9986 11506 9998
rect 13918 10050 13970 10062
rect 13918 9986 13970 9998
rect 14030 10050 14082 10062
rect 14030 9986 14082 9998
rect 14254 10050 14306 10062
rect 14254 9986 14306 9998
rect 21870 10050 21922 10062
rect 21870 9986 21922 9998
rect 23214 10050 23266 10062
rect 23214 9986 23266 9998
rect 5966 9938 6018 9950
rect 32622 9938 32674 9950
rect 19282 9886 19294 9938
rect 19346 9886 19358 9938
rect 30258 9886 30270 9938
rect 30322 9886 30334 9938
rect 5966 9874 6018 9886
rect 32622 9874 32674 9886
rect 7982 9826 8034 9838
rect 12910 9826 12962 9838
rect 16830 9826 16882 9838
rect 22990 9826 23042 9838
rect 32062 9826 32114 9838
rect 34638 9826 34690 9838
rect 39902 9826 39954 9838
rect 8418 9774 8430 9826
rect 8482 9774 8494 9826
rect 15474 9774 15486 9826
rect 15538 9774 15550 9826
rect 15922 9774 15934 9826
rect 15986 9774 15998 9826
rect 17266 9774 17278 9826
rect 17330 9774 17342 9826
rect 18274 9774 18286 9826
rect 18338 9774 18350 9826
rect 20178 9774 20190 9826
rect 20242 9774 20254 9826
rect 21298 9774 21310 9826
rect 21362 9774 21374 9826
rect 24434 9774 24446 9826
rect 24498 9774 24510 9826
rect 24770 9774 24782 9826
rect 24834 9774 24846 9826
rect 26114 9774 26126 9826
rect 26178 9774 26190 9826
rect 27122 9774 27134 9826
rect 27186 9774 27198 9826
rect 29586 9774 29598 9826
rect 29650 9774 29662 9826
rect 31154 9774 31166 9826
rect 31218 9774 31230 9826
rect 33282 9774 33294 9826
rect 33346 9774 33358 9826
rect 33730 9774 33742 9826
rect 33794 9774 33806 9826
rect 35074 9774 35086 9826
rect 35138 9774 35150 9826
rect 35970 9774 35982 9826
rect 36034 9774 36046 9826
rect 38770 9774 38782 9826
rect 38834 9774 38846 9826
rect 39330 9774 39342 9826
rect 39394 9774 39406 9826
rect 40674 9774 40686 9826
rect 40738 9774 40750 9826
rect 41570 9774 41582 9826
rect 41634 9774 41646 9826
rect 7982 9762 8034 9774
rect 12910 9762 12962 9774
rect 16830 9762 16882 9774
rect 22990 9762 23042 9774
rect 32062 9762 32114 9774
rect 34638 9762 34690 9774
rect 39902 9762 39954 9774
rect 4286 9714 4338 9726
rect 4286 9650 4338 9662
rect 4958 9714 5010 9726
rect 4958 9650 5010 9662
rect 10670 9714 10722 9726
rect 10670 9650 10722 9662
rect 12574 9714 12626 9726
rect 15150 9714 15202 9726
rect 23998 9714 24050 9726
rect 25454 9714 25506 9726
rect 31390 9714 31442 9726
rect 32958 9714 33010 9726
rect 38446 9714 38498 9726
rect 14802 9662 14814 9714
rect 14866 9662 14878 9714
rect 19954 9662 19966 9714
rect 20018 9662 20030 9714
rect 23538 9662 23550 9714
rect 23602 9662 23614 9714
rect 24994 9662 25006 9714
rect 25058 9662 25070 9714
rect 29810 9662 29822 9714
rect 29874 9662 29886 9714
rect 31714 9662 31726 9714
rect 31778 9662 31790 9714
rect 33954 9662 33966 9714
rect 34018 9662 34030 9714
rect 39442 9662 39454 9714
rect 39506 9662 39518 9714
rect 12574 9650 12626 9662
rect 15150 9650 15202 9662
rect 23998 9650 24050 9662
rect 25454 9650 25506 9662
rect 31390 9650 31442 9662
rect 32958 9650 33010 9662
rect 38446 9650 38498 9662
rect 4174 9602 4226 9614
rect 4174 9538 4226 9550
rect 4846 9602 4898 9614
rect 20638 9602 20690 9614
rect 16146 9550 16158 9602
rect 16210 9550 16222 9602
rect 4846 9538 4898 9550
rect 20638 9538 20690 9550
rect 30718 9602 30770 9614
rect 30718 9538 30770 9550
rect 1344 9434 46592 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 46592 9434
rect 1344 9348 46592 9382
rect 2942 9266 2994 9278
rect 9886 9266 9938 9278
rect 3714 9214 3726 9266
rect 3778 9214 3790 9266
rect 2942 9202 2994 9214
rect 9886 9202 9938 9214
rect 18174 9266 18226 9278
rect 18174 9202 18226 9214
rect 30942 9266 30994 9278
rect 30942 9202 30994 9214
rect 31726 9266 31778 9278
rect 32398 9266 32450 9278
rect 38558 9266 38610 9278
rect 32050 9214 32062 9266
rect 32114 9214 32126 9266
rect 33394 9214 33406 9266
rect 33458 9214 33470 9266
rect 31726 9202 31778 9214
rect 32398 9202 32450 9214
rect 38558 9202 38610 9214
rect 43374 9266 43426 9278
rect 43374 9202 43426 9214
rect 23326 9154 23378 9166
rect 13570 9102 13582 9154
rect 13634 9102 13646 9154
rect 15586 9102 15598 9154
rect 15650 9102 15662 9154
rect 18610 9102 18622 9154
rect 18674 9102 18686 9154
rect 19058 9102 19070 9154
rect 19122 9102 19134 9154
rect 23326 9090 23378 9102
rect 26126 9154 26178 9166
rect 26126 9090 26178 9102
rect 29598 9154 29650 9166
rect 41806 9154 41858 9166
rect 37538 9102 37550 9154
rect 37602 9102 37614 9154
rect 41234 9102 41246 9154
rect 41298 9102 41310 9154
rect 29598 9090 29650 9102
rect 41806 9090 41858 9102
rect 6638 9042 6690 9054
rect 5954 8990 5966 9042
rect 6018 8990 6030 9042
rect 6638 8978 6690 8990
rect 9998 9042 10050 9054
rect 14366 9042 14418 9054
rect 13458 8990 13470 9042
rect 13522 8990 13534 9042
rect 9998 8978 10050 8990
rect 14366 8978 14418 8990
rect 20638 9042 20690 9054
rect 20638 8978 20690 8990
rect 22990 9042 23042 9054
rect 22990 8978 23042 8990
rect 23662 9042 23714 9054
rect 25230 9042 25282 9054
rect 24098 8990 24110 9042
rect 24162 8990 24174 9042
rect 26226 8990 26238 9042
rect 26290 8990 26302 9042
rect 29810 8990 29822 9042
rect 29874 8990 29886 9042
rect 33170 8990 33182 9042
rect 33234 8990 33246 9042
rect 34850 8990 34862 9042
rect 34914 8990 34926 9042
rect 35410 8990 35422 9042
rect 35474 8990 35486 9042
rect 23662 8978 23714 8990
rect 25230 8978 25282 8990
rect 14478 8930 14530 8942
rect 20178 8878 20190 8930
rect 20242 8878 20254 8930
rect 25666 8878 25678 8930
rect 25730 8878 25742 8930
rect 31266 8878 31278 8930
rect 31330 8878 31342 8930
rect 41570 8878 41582 8930
rect 41634 8878 41646 8930
rect 14478 8866 14530 8878
rect 19294 8818 19346 8830
rect 19294 8754 19346 8766
rect 19630 8818 19682 8830
rect 19630 8754 19682 8766
rect 1344 8650 46592 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 46592 8650
rect 1344 8564 46592 8598
rect 23326 8370 23378 8382
rect 13570 8318 13582 8370
rect 13634 8318 13646 8370
rect 15810 8318 15822 8370
rect 15874 8318 15886 8370
rect 35074 8318 35086 8370
rect 35138 8318 35150 8370
rect 23326 8306 23378 8318
rect 18734 8258 18786 8270
rect 20302 8258 20354 8270
rect 13682 8206 13694 8258
rect 13746 8206 13758 8258
rect 15026 8206 15038 8258
rect 15090 8206 15102 8258
rect 19170 8206 19182 8258
rect 19234 8206 19246 8258
rect 19730 8206 19742 8258
rect 19794 8206 19806 8258
rect 18734 8194 18786 8206
rect 20302 8194 20354 8206
rect 21646 8258 21698 8270
rect 21646 8194 21698 8206
rect 22990 8258 23042 8270
rect 26910 8258 26962 8270
rect 31278 8258 31330 8270
rect 35758 8258 35810 8270
rect 24882 8206 24894 8258
rect 24946 8206 24958 8258
rect 30818 8206 30830 8258
rect 30882 8206 30894 8258
rect 31826 8206 31838 8258
rect 31890 8206 31902 8258
rect 37874 8206 37886 8258
rect 37938 8206 37950 8258
rect 38434 8206 38446 8258
rect 38498 8206 38510 8258
rect 40898 8206 40910 8258
rect 40962 8206 40974 8258
rect 22990 8194 23042 8206
rect 26910 8194 26962 8206
rect 31278 8194 31330 8206
rect 35758 8194 35810 8206
rect 19966 8146 20018 8158
rect 24670 8146 24722 8158
rect 26686 8146 26738 8158
rect 30606 8146 30658 8158
rect 22306 8094 22318 8146
rect 22370 8094 22382 8146
rect 22754 8094 22766 8146
rect 22818 8094 22830 8146
rect 25106 8094 25118 8146
rect 25170 8094 25182 8146
rect 27010 8094 27022 8146
rect 27074 8094 27086 8146
rect 27570 8094 27582 8146
rect 27634 8094 27646 8146
rect 34066 8094 34078 8146
rect 34130 8094 34142 8146
rect 19966 8082 20018 8094
rect 24670 8082 24722 8094
rect 26686 8082 26738 8094
rect 30606 8082 30658 8094
rect 20638 8034 20690 8046
rect 23886 8034 23938 8046
rect 36094 8034 36146 8046
rect 18946 7982 18958 8034
rect 19010 7982 19022 8034
rect 21298 7982 21310 8034
rect 21362 7982 21374 8034
rect 24210 7982 24222 8034
rect 24274 7982 24286 8034
rect 25890 7982 25902 8034
rect 25954 7982 25966 8034
rect 20638 7970 20690 7982
rect 23886 7970 23938 7982
rect 36094 7970 36146 7982
rect 1344 7866 46592 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 46592 7866
rect 1344 7780 46592 7814
rect 5518 7698 5570 7710
rect 4946 7646 4958 7698
rect 5010 7646 5022 7698
rect 5518 7634 5570 7646
rect 21982 7698 22034 7710
rect 35534 7698 35586 7710
rect 26786 7646 26798 7698
rect 26850 7646 26862 7698
rect 32386 7646 32398 7698
rect 32450 7646 32462 7698
rect 38546 7646 38558 7698
rect 38610 7646 38622 7698
rect 21982 7634 22034 7646
rect 35534 7634 35586 7646
rect 19070 7586 19122 7598
rect 25790 7586 25842 7598
rect 19842 7534 19854 7586
rect 19906 7534 19918 7586
rect 21298 7534 21310 7586
rect 21362 7534 21374 7586
rect 19070 7522 19122 7534
rect 25790 7522 25842 7534
rect 27246 7586 27298 7598
rect 30146 7534 30158 7586
rect 30210 7534 30222 7586
rect 27246 7522 27298 7534
rect 2046 7474 2098 7486
rect 22878 7474 22930 7486
rect 2482 7422 2494 7474
rect 2546 7422 2558 7474
rect 18834 7422 18846 7474
rect 18898 7422 18910 7474
rect 2046 7410 2098 7422
rect 22878 7410 22930 7422
rect 24110 7474 24162 7486
rect 24110 7410 24162 7422
rect 24670 7474 24722 7486
rect 33966 7474 34018 7486
rect 35646 7474 35698 7486
rect 26114 7422 26126 7474
rect 26178 7422 26190 7474
rect 26674 7422 26686 7474
rect 26738 7422 26750 7474
rect 28018 7422 28030 7474
rect 28082 7422 28094 7474
rect 28802 7422 28814 7474
rect 28866 7422 28878 7474
rect 29474 7422 29486 7474
rect 29538 7422 29550 7474
rect 33618 7422 33630 7474
rect 33682 7422 33694 7474
rect 34290 7422 34302 7474
rect 34354 7422 34366 7474
rect 36194 7422 36206 7474
rect 36258 7422 36270 7474
rect 24670 7410 24722 7422
rect 33966 7410 34018 7422
rect 35646 7410 35698 7422
rect 21646 7362 21698 7374
rect 23438 7362 23490 7374
rect 19506 7310 19518 7362
rect 19570 7310 19582 7362
rect 22418 7310 22430 7362
rect 22482 7310 22494 7362
rect 21646 7298 21698 7310
rect 23438 7298 23490 7310
rect 39342 7250 39394 7262
rect 39342 7186 39394 7198
rect 1344 7082 46592 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 46592 7082
rect 1344 6996 46592 7030
rect 28018 6862 28030 6914
rect 28082 6862 28094 6914
rect 33730 6862 33742 6914
rect 33794 6862 33806 6914
rect 19282 6750 19294 6802
rect 19346 6750 19358 6802
rect 24894 6690 24946 6702
rect 15474 6638 15486 6690
rect 15538 6638 15550 6690
rect 21634 6638 21646 6690
rect 21698 6638 21710 6690
rect 22082 6638 22094 6690
rect 22146 6638 22158 6690
rect 22866 6638 22878 6690
rect 22930 6638 22942 6690
rect 23314 6638 23326 6690
rect 23378 6638 23390 6690
rect 24434 6638 24446 6690
rect 24498 6638 24510 6690
rect 24894 6626 24946 6638
rect 25454 6690 25506 6702
rect 29486 6690 29538 6702
rect 28354 6638 28366 6690
rect 28418 6638 28430 6690
rect 30146 6638 30158 6690
rect 30210 6638 30222 6690
rect 30594 6638 30606 6690
rect 30658 6638 30670 6690
rect 32834 6638 32846 6690
rect 32898 6638 32910 6690
rect 25454 6626 25506 6638
rect 29486 6626 29538 6638
rect 20638 6578 20690 6590
rect 19842 6526 19854 6578
rect 19906 6526 19918 6578
rect 20638 6514 20690 6526
rect 21310 6578 21362 6590
rect 22306 6526 22318 6578
rect 22370 6526 22382 6578
rect 29138 6526 29150 6578
rect 29202 6526 29214 6578
rect 21310 6514 21362 6526
rect 18274 6414 18286 6466
rect 18338 6414 18350 6466
rect 1344 6298 46592 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 46592 6298
rect 1344 6212 46592 6246
rect 5854 6130 5906 6142
rect 25342 6130 25394 6142
rect 5058 6078 5070 6130
rect 5122 6078 5134 6130
rect 22418 6078 22430 6130
rect 22482 6078 22494 6130
rect 5854 6066 5906 6078
rect 25342 6066 25394 6078
rect 15934 6018 15986 6030
rect 15934 5954 15986 5966
rect 16158 6018 16210 6030
rect 16158 5954 16210 5966
rect 17502 6018 17554 6030
rect 18498 5966 18510 6018
rect 18562 5966 18574 6018
rect 19842 5966 19854 6018
rect 19906 5966 19918 6018
rect 17502 5954 17554 5966
rect 2158 5906 2210 5918
rect 15598 5906 15650 5918
rect 21198 5906 21250 5918
rect 22878 5906 22930 5918
rect 25678 5906 25730 5918
rect 2706 5854 2718 5906
rect 2770 5854 2782 5906
rect 16370 5854 16382 5906
rect 16434 5854 16446 5906
rect 18610 5854 18622 5906
rect 18674 5854 18686 5906
rect 21746 5854 21758 5906
rect 21810 5854 21822 5906
rect 22194 5854 22206 5906
rect 22258 5854 22270 5906
rect 23650 5854 23662 5906
rect 23714 5854 23726 5906
rect 24546 5854 24558 5906
rect 24610 5854 24622 5906
rect 25218 5854 25230 5906
rect 25282 5854 25294 5906
rect 27570 5854 27582 5906
rect 27634 5854 27646 5906
rect 2158 5842 2210 5854
rect 15598 5842 15650 5854
rect 21198 5842 21250 5854
rect 22878 5842 22930 5854
rect 25678 5842 25730 5854
rect 21422 5794 21474 5806
rect 28802 5742 28814 5794
rect 28866 5742 28878 5794
rect 21422 5730 21474 5742
rect 25454 5682 25506 5694
rect 16706 5630 16718 5682
rect 16770 5630 16782 5682
rect 25454 5618 25506 5630
rect 1344 5514 46592 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 46592 5514
rect 1344 5428 46592 5462
rect 27582 5346 27634 5358
rect 27582 5282 27634 5294
rect 21410 5182 21422 5234
rect 21474 5182 21486 5234
rect 22978 5182 22990 5234
rect 23042 5182 23054 5234
rect 24546 5182 24558 5234
rect 24610 5182 24622 5234
rect 15262 5122 15314 5134
rect 15262 5058 15314 5070
rect 20414 5122 20466 5134
rect 21522 5070 21534 5122
rect 21586 5070 21598 5122
rect 23538 5070 23550 5122
rect 23602 5070 23614 5122
rect 24994 5070 25006 5122
rect 25058 5070 25070 5122
rect 28578 5070 28590 5122
rect 28642 5070 28654 5122
rect 20414 5058 20466 5070
rect 20750 5010 20802 5022
rect 23874 4958 23886 5010
rect 23938 4958 23950 5010
rect 24882 4958 24894 5010
rect 24946 4958 24958 5010
rect 20750 4946 20802 4958
rect 1710 4898 1762 4910
rect 18498 4846 18510 4898
rect 18562 4846 18574 4898
rect 1710 4834 1762 4846
rect 1344 4730 46592 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 46592 4730
rect 1344 4644 46592 4678
rect 22094 4562 22146 4574
rect 19618 4510 19630 4562
rect 19682 4510 19694 4562
rect 23650 4510 23662 4562
rect 23714 4510 23726 4562
rect 22094 4498 22146 4510
rect 19182 4450 19234 4462
rect 19182 4386 19234 4398
rect 20638 4450 20690 4462
rect 20638 4386 20690 4398
rect 20974 4450 21026 4462
rect 23090 4398 23102 4450
rect 23154 4398 23166 4450
rect 24658 4398 24670 4450
rect 24722 4398 24734 4450
rect 20974 4386 21026 4398
rect 21422 4338 21474 4350
rect 17490 4286 17502 4338
rect 17554 4286 17566 4338
rect 18498 4286 18510 4338
rect 18562 4286 18574 4338
rect 19730 4286 19742 4338
rect 19794 4286 19806 4338
rect 20290 4286 20302 4338
rect 20354 4286 20366 4338
rect 21422 4274 21474 4286
rect 21646 4338 21698 4350
rect 24110 4338 24162 4350
rect 23538 4286 23550 4338
rect 23602 4286 23614 4338
rect 21646 4274 21698 4286
rect 24110 4274 24162 4286
rect 21198 4114 21250 4126
rect 21198 4050 21250 4062
rect 1344 3946 46592 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 46592 3946
rect 1344 3860 46592 3894
rect 19854 3554 19906 3566
rect 19854 3490 19906 3502
rect 19506 3390 19518 3442
rect 19570 3390 19582 3442
rect 1344 3162 46592 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 46592 3162
rect 1344 3076 46592 3110
<< via1 >>
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 1710 43710 1762 43762
rect 28366 43710 28418 43762
rect 13246 43598 13298 43650
rect 28254 43598 28306 43650
rect 30494 43598 30546 43650
rect 13022 43486 13074 43538
rect 19182 43486 19234 43538
rect 25342 43486 25394 43538
rect 26126 43486 26178 43538
rect 29486 43486 29538 43538
rect 30830 43486 30882 43538
rect 19854 43374 19906 43426
rect 22318 43374 22370 43426
rect 25790 43374 25842 43426
rect 28702 43374 28754 43426
rect 27246 43262 27298 43314
rect 30270 43262 30322 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 13582 42702 13634 42754
rect 14926 42702 14978 42754
rect 20078 42702 20130 42754
rect 21982 42702 22034 42754
rect 22430 42702 22482 42754
rect 22878 42702 22930 42754
rect 23326 42702 23378 42754
rect 29262 42702 29314 42754
rect 30494 42702 30546 42754
rect 17950 42590 18002 42642
rect 19742 42590 19794 42642
rect 20750 42590 20802 42642
rect 25566 42590 25618 42642
rect 26686 42590 26738 42642
rect 27918 42590 27970 42642
rect 28478 42590 28530 42642
rect 33518 42590 33570 42642
rect 1710 42478 1762 42530
rect 20414 42478 20466 42530
rect 28142 42478 28194 42530
rect 46174 42478 46226 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 33518 42030 33570 42082
rect 12798 41918 12850 41970
rect 14142 41918 14194 41970
rect 19518 41918 19570 41970
rect 20190 41918 20242 41970
rect 22990 41918 23042 41970
rect 23438 41918 23490 41970
rect 25678 41918 25730 41970
rect 26462 41918 26514 41970
rect 30046 41918 30098 41970
rect 30606 41918 30658 41970
rect 30830 41918 30882 41970
rect 31726 41918 31778 41970
rect 32510 41918 32562 41970
rect 16046 41806 16098 41858
rect 18510 41806 18562 41858
rect 28926 41806 28978 41858
rect 24222 41694 24274 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 13694 41134 13746 41186
rect 14142 41134 14194 41186
rect 14590 41134 14642 41186
rect 23438 41134 23490 41186
rect 24110 41134 24162 41186
rect 26350 41134 26402 41186
rect 26910 41134 26962 41186
rect 29486 41134 29538 41186
rect 29934 41134 29986 41186
rect 31390 41134 31442 41186
rect 32286 41134 32338 41186
rect 19294 41022 19346 41074
rect 19630 41022 19682 41074
rect 22878 41022 22930 41074
rect 23214 41022 23266 41074
rect 27582 41022 27634 41074
rect 29150 41022 29202 41074
rect 30606 41022 30658 41074
rect 12574 40910 12626 40962
rect 12910 40910 12962 40962
rect 13470 40910 13522 40962
rect 17390 40910 17442 40962
rect 18062 40910 18114 40962
rect 19070 40910 19122 40962
rect 27918 40910 27970 40962
rect 28254 40910 28306 40962
rect 30158 40910 30210 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 24110 40574 24162 40626
rect 11454 40462 11506 40514
rect 12126 40462 12178 40514
rect 12574 40462 12626 40514
rect 15934 40462 15986 40514
rect 26798 40462 26850 40514
rect 27806 40462 27858 40514
rect 30382 40462 30434 40514
rect 37886 40462 37938 40514
rect 11230 40350 11282 40402
rect 11902 40350 11954 40402
rect 14254 40350 14306 40402
rect 15150 40350 15202 40402
rect 16270 40350 16322 40402
rect 17390 40350 17442 40402
rect 19406 40350 19458 40402
rect 19854 40350 19906 40402
rect 22094 40350 22146 40402
rect 23886 40350 23938 40402
rect 27134 40350 27186 40402
rect 27582 40350 27634 40402
rect 28478 40350 28530 40402
rect 28926 40350 28978 40402
rect 29934 40350 29986 40402
rect 30830 40350 30882 40402
rect 31278 40350 31330 40402
rect 31838 40350 31890 40402
rect 35086 40350 35138 40402
rect 35534 40350 35586 40402
rect 13918 40238 13970 40290
rect 18286 40238 18338 40290
rect 15486 40126 15538 40178
rect 23102 40126 23154 40178
rect 38670 40126 38722 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 34190 39790 34242 39842
rect 13694 39678 13746 39730
rect 22094 39678 22146 39730
rect 22430 39678 22482 39730
rect 37662 39678 37714 39730
rect 14366 39566 14418 39618
rect 15038 39566 15090 39618
rect 15598 39566 15650 39618
rect 16158 39566 16210 39618
rect 19406 39566 19458 39618
rect 21310 39566 21362 39618
rect 22766 39566 22818 39618
rect 23214 39566 23266 39618
rect 24110 39566 24162 39618
rect 24446 39566 24498 39618
rect 25566 39566 25618 39618
rect 28030 39566 28082 39618
rect 29822 39566 29874 39618
rect 30046 39566 30098 39618
rect 33630 39566 33682 39618
rect 9214 39454 9266 39506
rect 19070 39454 19122 39506
rect 21646 39454 21698 39506
rect 27694 39454 27746 39506
rect 28254 39454 28306 39506
rect 29374 39454 29426 39506
rect 33182 39454 33234 39506
rect 37326 39454 37378 39506
rect 37886 39454 37938 39506
rect 38670 39454 38722 39506
rect 39454 39454 39506 39506
rect 12798 39342 12850 39394
rect 14814 39342 14866 39394
rect 15262 39342 15314 39394
rect 20526 39342 20578 39394
rect 23438 39342 23490 39394
rect 29150 39342 29202 39394
rect 34750 39342 34802 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 4846 39006 4898 39058
rect 21758 39006 21810 39058
rect 29374 39006 29426 39058
rect 39454 39006 39506 39058
rect 11678 38894 11730 38946
rect 16718 38894 16770 38946
rect 18398 38894 18450 38946
rect 20974 38894 21026 38946
rect 21310 38894 21362 38946
rect 22430 38894 22482 38946
rect 23998 38894 24050 38946
rect 27582 38894 27634 38946
rect 32510 38894 32562 38946
rect 1934 38782 1986 38834
rect 2382 38782 2434 38834
rect 14366 38782 14418 38834
rect 15262 38782 15314 38834
rect 16270 38782 16322 38834
rect 17726 38782 17778 38834
rect 18286 38782 18338 38834
rect 19070 38782 19122 38834
rect 19630 38782 19682 38834
rect 20526 38782 20578 38834
rect 22206 38782 22258 38834
rect 23214 38782 23266 38834
rect 23774 38782 23826 38834
rect 32286 38782 32338 38834
rect 33070 38782 33122 38834
rect 33518 38782 33570 38834
rect 35870 38782 35922 38834
rect 36318 38782 36370 38834
rect 37774 38782 37826 38834
rect 38558 38782 38610 38834
rect 39118 38782 39170 38834
rect 39678 38782 39730 38834
rect 41582 38782 41634 38834
rect 41806 38782 41858 38834
rect 13806 38670 13858 38722
rect 17390 38670 17442 38722
rect 24558 38670 24610 38722
rect 38222 38670 38274 38722
rect 41134 38670 41186 38722
rect 41358 38670 41410 38722
rect 41694 38670 41746 38722
rect 5406 38558 5458 38610
rect 22878 38558 22930 38610
rect 37214 38558 37266 38610
rect 40910 38558 40962 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 14814 38110 14866 38162
rect 20190 38110 20242 38162
rect 22094 38110 22146 38162
rect 43150 38110 43202 38162
rect 13694 37998 13746 38050
rect 15150 37998 15202 38050
rect 15598 37998 15650 38050
rect 16494 37998 16546 38050
rect 16830 37998 16882 38050
rect 17950 37998 18002 38050
rect 19182 37998 19234 38050
rect 20638 37998 20690 38050
rect 22542 37998 22594 38050
rect 22990 37998 23042 38050
rect 23438 37998 23490 38050
rect 31726 37998 31778 38050
rect 32510 37998 32562 38050
rect 37326 37998 37378 38050
rect 37774 37998 37826 38050
rect 39006 37998 39058 38050
rect 40014 37998 40066 38050
rect 40910 37998 40962 38050
rect 42478 37998 42530 38050
rect 42702 37998 42754 38050
rect 13470 37886 13522 37938
rect 18846 37886 18898 37938
rect 21310 37886 21362 37938
rect 23886 37886 23938 37938
rect 34638 37886 34690 37938
rect 36094 37886 36146 37938
rect 36990 37886 37042 37938
rect 38446 37886 38498 37938
rect 43710 37886 43762 37938
rect 15822 37774 15874 37826
rect 19518 37774 19570 37826
rect 19854 37774 19906 37826
rect 21646 37774 21698 37826
rect 24222 37774 24274 37826
rect 24558 37774 24610 37826
rect 24894 37774 24946 37826
rect 25230 37774 25282 37826
rect 37998 37774 38050 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 5406 37438 5458 37490
rect 13470 37438 13522 37490
rect 14702 37438 14754 37490
rect 22542 37438 22594 37490
rect 25790 37438 25842 37490
rect 29710 37438 29762 37490
rect 30046 37438 30098 37490
rect 38558 37438 38610 37490
rect 41694 37438 41746 37490
rect 16046 37326 16098 37378
rect 18958 37326 19010 37378
rect 19742 37326 19794 37378
rect 21310 37326 21362 37378
rect 24446 37326 24498 37378
rect 28366 37326 28418 37378
rect 32398 37326 32450 37378
rect 34638 37326 34690 37378
rect 40350 37326 40402 37378
rect 40910 37326 40962 37378
rect 2718 37214 2770 37266
rect 3166 37214 3218 37266
rect 10782 37214 10834 37266
rect 11230 37214 11282 37266
rect 15038 37214 15090 37266
rect 15710 37214 15762 37266
rect 17838 37214 17890 37266
rect 18734 37214 18786 37266
rect 22878 37214 22930 37266
rect 23438 37214 23490 37266
rect 23998 37214 24050 37266
rect 24558 37214 24610 37266
rect 26126 37214 26178 37266
rect 26462 37214 26514 37266
rect 28702 37214 28754 37266
rect 30382 37214 30434 37266
rect 31278 37214 31330 37266
rect 32174 37214 32226 37266
rect 34414 37214 34466 37266
rect 35422 37214 35474 37266
rect 35870 37214 35922 37266
rect 36654 37214 36706 37266
rect 37662 37214 37714 37266
rect 38894 37214 38946 37266
rect 40014 37214 40066 37266
rect 41246 37214 41298 37266
rect 43150 37214 43202 37266
rect 44158 37214 44210 37266
rect 14366 37102 14418 37154
rect 16494 37102 16546 37154
rect 17390 37102 17442 37154
rect 19518 37102 19570 37154
rect 21982 37102 22034 37154
rect 25342 37102 25394 37154
rect 29262 37102 29314 37154
rect 31614 37102 31666 37154
rect 33966 37102 34018 37154
rect 35758 37102 35810 37154
rect 37438 37102 37490 37154
rect 38110 37102 38162 37154
rect 39566 37102 39618 37154
rect 42030 37102 42082 37154
rect 6190 36990 6242 37042
rect 24334 36990 24386 37042
rect 26126 36990 26178 37042
rect 36542 36990 36594 37042
rect 42814 36990 42866 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 22318 36654 22370 36706
rect 35422 36654 35474 36706
rect 12910 36542 12962 36594
rect 13694 36542 13746 36594
rect 15486 36542 15538 36594
rect 17838 36542 17890 36594
rect 19630 36542 19682 36594
rect 28142 36542 28194 36594
rect 35982 36542 36034 36594
rect 37102 36542 37154 36594
rect 43374 36542 43426 36594
rect 9438 36430 9490 36482
rect 10110 36430 10162 36482
rect 14254 36430 14306 36482
rect 19518 36430 19570 36482
rect 21646 36430 21698 36482
rect 21870 36430 21922 36482
rect 22094 36430 22146 36482
rect 25118 36430 25170 36482
rect 25454 36430 25506 36482
rect 29486 36430 29538 36482
rect 29934 36430 29986 36482
rect 30606 36430 30658 36482
rect 31390 36430 31442 36482
rect 32286 36430 32338 36482
rect 32958 36430 33010 36482
rect 34302 36430 34354 36482
rect 36206 36430 36258 36482
rect 38558 36430 38610 36482
rect 39454 36430 39506 36482
rect 39790 36430 39842 36482
rect 43038 36430 43090 36482
rect 43262 36430 43314 36482
rect 43486 36430 43538 36482
rect 6302 36318 6354 36370
rect 6638 36318 6690 36370
rect 7086 36318 7138 36370
rect 9662 36318 9714 36370
rect 10782 36318 10834 36370
rect 15262 36318 15314 36370
rect 16494 36318 16546 36370
rect 19630 36318 19682 36370
rect 20750 36318 20802 36370
rect 23550 36318 23602 36370
rect 26574 36318 26626 36370
rect 29150 36318 29202 36370
rect 38110 36318 38162 36370
rect 39230 36318 39282 36370
rect 40686 36318 40738 36370
rect 41022 36318 41074 36370
rect 5182 36206 5234 36258
rect 5630 36206 5682 36258
rect 5966 36206 6018 36258
rect 6974 36206 7026 36258
rect 15374 36206 15426 36258
rect 22766 36206 22818 36258
rect 24894 36206 24946 36258
rect 27806 36206 27858 36258
rect 28590 36206 28642 36258
rect 30158 36206 30210 36258
rect 37550 36206 37602 36258
rect 38558 36206 38610 36258
rect 40126 36206 40178 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 6750 35870 6802 35922
rect 7534 35870 7586 35922
rect 10110 35870 10162 35922
rect 15486 35870 15538 35922
rect 16494 35870 16546 35922
rect 19630 35870 19682 35922
rect 19966 35870 20018 35922
rect 27358 35870 27410 35922
rect 31838 35870 31890 35922
rect 39118 35870 39170 35922
rect 39902 35870 39954 35922
rect 43038 35870 43090 35922
rect 15822 35758 15874 35810
rect 17614 35758 17666 35810
rect 21198 35758 21250 35810
rect 22206 35758 22258 35810
rect 26686 35758 26738 35810
rect 30942 35758 30994 35810
rect 35534 35758 35586 35810
rect 36542 35758 36594 35810
rect 41134 35758 41186 35810
rect 41470 35758 41522 35810
rect 44830 35758 44882 35810
rect 3838 35646 3890 35698
rect 4510 35646 4562 35698
rect 10670 35646 10722 35698
rect 12910 35646 12962 35698
rect 13470 35646 13522 35698
rect 16718 35646 16770 35698
rect 17502 35646 17554 35698
rect 20862 35646 20914 35698
rect 21534 35646 21586 35698
rect 21982 35646 22034 35698
rect 22878 35646 22930 35698
rect 23326 35646 23378 35698
rect 24334 35646 24386 35698
rect 25902 35646 25954 35698
rect 26350 35646 26402 35698
rect 27134 35646 27186 35698
rect 27694 35646 27746 35698
rect 28254 35646 28306 35698
rect 34190 35646 34242 35698
rect 34750 35646 34802 35698
rect 35982 35646 36034 35698
rect 36430 35646 36482 35698
rect 37214 35646 37266 35698
rect 37774 35646 37826 35698
rect 38558 35646 38610 35698
rect 39342 35646 39394 35698
rect 42702 35646 42754 35698
rect 43486 35646 43538 35698
rect 3614 35534 3666 35586
rect 7870 35534 7922 35586
rect 19182 35534 19234 35586
rect 20414 35534 20466 35586
rect 42366 35534 42418 35586
rect 44718 35534 44770 35586
rect 7758 35422 7810 35474
rect 14590 35422 14642 35474
rect 18286 35422 18338 35474
rect 18622 35422 18674 35474
rect 25566 35422 25618 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 2942 35086 2994 35138
rect 9214 35086 9266 35138
rect 28478 35086 28530 35138
rect 33182 35086 33234 35138
rect 3054 34974 3106 35026
rect 22878 34974 22930 35026
rect 26574 34974 26626 35026
rect 27134 34974 27186 35026
rect 37998 34974 38050 35026
rect 38222 34974 38274 35026
rect 41470 34974 41522 35026
rect 3502 34862 3554 34914
rect 5518 34862 5570 34914
rect 6190 34862 6242 34914
rect 14590 34862 14642 34914
rect 14926 34862 14978 34914
rect 15374 34862 15426 34914
rect 16606 34862 16658 34914
rect 17726 34862 17778 34914
rect 23214 34862 23266 34914
rect 23774 34862 23826 34914
rect 24334 34862 24386 34914
rect 24894 34862 24946 34914
rect 26014 34862 26066 34914
rect 29150 34862 29202 34914
rect 29374 34862 29426 34914
rect 29710 34862 29762 34914
rect 30158 34862 30210 34914
rect 37438 34862 37490 34914
rect 38670 34862 38722 34914
rect 39118 34862 39170 34914
rect 39454 34862 39506 34914
rect 40126 34862 40178 34914
rect 41022 34862 41074 34914
rect 41918 34862 41970 34914
rect 42702 34862 42754 34914
rect 1710 34750 1762 34802
rect 2046 34750 2098 34802
rect 4734 34750 4786 34802
rect 11118 34750 11170 34802
rect 11454 34750 11506 34802
rect 15598 34750 15650 34802
rect 16046 34750 16098 34802
rect 22542 34750 22594 34802
rect 27582 34750 27634 34802
rect 37662 34750 37714 34802
rect 39790 34750 39842 34802
rect 40462 34750 40514 34802
rect 43934 34750 43986 34802
rect 45166 34750 45218 34802
rect 2494 34638 2546 34690
rect 3726 34638 3778 34690
rect 4062 34638 4114 34690
rect 4398 34638 4450 34690
rect 5070 34638 5122 34690
rect 8430 34638 8482 34690
rect 21982 34638 22034 34690
rect 23886 34638 23938 34690
rect 37102 34638 37154 34690
rect 37214 34638 37266 34690
rect 37774 34638 37826 34690
rect 44830 34638 44882 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4734 34302 4786 34354
rect 8318 34302 8370 34354
rect 23326 34302 23378 34354
rect 23886 34302 23938 34354
rect 25566 34302 25618 34354
rect 29934 34302 29986 34354
rect 39454 34302 39506 34354
rect 41134 34302 41186 34354
rect 13694 34190 13746 34242
rect 15598 34190 15650 34242
rect 15822 34190 15874 34242
rect 16158 34190 16210 34242
rect 16830 34190 16882 34242
rect 17838 34190 17890 34242
rect 18174 34190 18226 34242
rect 22094 34190 22146 34242
rect 22430 34190 22482 34242
rect 25230 34190 25282 34242
rect 26462 34190 26514 34242
rect 37662 34190 37714 34242
rect 38334 34190 38386 34242
rect 44942 34190 44994 34242
rect 1822 34078 1874 34130
rect 2158 34078 2210 34130
rect 5630 34078 5682 34130
rect 6078 34078 6130 34130
rect 9102 34078 9154 34130
rect 9662 34078 9714 34130
rect 10782 34078 10834 34130
rect 11342 34078 11394 34130
rect 16494 34078 16546 34130
rect 23214 34078 23266 34130
rect 23438 34078 23490 34130
rect 37438 34078 37490 34130
rect 37998 34078 38050 34130
rect 39790 34078 39842 34130
rect 40238 34078 40290 34130
rect 40910 34078 40962 34130
rect 41470 34078 41522 34130
rect 41806 34078 41858 34130
rect 45390 34078 45442 34130
rect 19294 33966 19346 34018
rect 24446 33966 24498 34018
rect 36990 33966 37042 34018
rect 38894 33966 38946 34018
rect 5294 33854 5346 33906
rect 9550 33854 9602 33906
rect 14478 33854 14530 33906
rect 18398 33854 18450 33906
rect 18734 33854 18786 33906
rect 22878 33854 22930 33906
rect 22990 33854 23042 33906
rect 45950 33854 46002 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 4174 33518 4226 33570
rect 4286 33406 4338 33458
rect 4958 33406 5010 33458
rect 24670 33406 24722 33458
rect 29262 33406 29314 33458
rect 5630 33294 5682 33346
rect 6078 33294 6130 33346
rect 6638 33294 6690 33346
rect 6974 33294 7026 33346
rect 10558 33294 10610 33346
rect 13470 33294 13522 33346
rect 13918 33294 13970 33346
rect 16942 33294 16994 33346
rect 17278 33294 17330 33346
rect 21310 33294 21362 33346
rect 21758 33294 21810 33346
rect 22430 33294 22482 33346
rect 25230 33294 25282 33346
rect 29038 33294 29090 33346
rect 32062 33294 32114 33346
rect 32398 33294 32450 33346
rect 41358 33294 41410 33346
rect 41806 33294 41858 33346
rect 42702 33294 42754 33346
rect 43262 33294 43314 33346
rect 44158 33294 44210 33346
rect 3726 33182 3778 33234
rect 3838 33182 3890 33234
rect 10334 33182 10386 33234
rect 22206 33182 22258 33234
rect 28254 33182 28306 33234
rect 29598 33182 29650 33234
rect 37102 33182 37154 33234
rect 38334 33182 38386 33234
rect 40798 33182 40850 33234
rect 41022 33182 41074 33234
rect 4846 33070 4898 33122
rect 9550 33070 9602 33122
rect 10110 33070 10162 33122
rect 18062 33070 18114 33122
rect 22766 33070 22818 33122
rect 24222 33070 24274 33122
rect 25454 33070 25506 33122
rect 28702 33070 28754 33122
rect 29374 33070 29426 33122
rect 34750 33070 34802 33122
rect 35534 33070 35586 33122
rect 37662 33070 37714 33122
rect 42030 33070 42082 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4734 32734 4786 32786
rect 5406 32734 5458 32786
rect 8542 32734 8594 32786
rect 12798 32734 12850 32786
rect 38110 32734 38162 32786
rect 39118 32734 39170 32786
rect 41022 32734 41074 32786
rect 8654 32622 8706 32674
rect 12238 32622 12290 32674
rect 22206 32622 22258 32674
rect 22542 32622 22594 32674
rect 24558 32622 24610 32674
rect 25678 32622 25730 32674
rect 28702 32622 28754 32674
rect 1934 32510 1986 32562
rect 2270 32510 2322 32562
rect 12014 32510 12066 32562
rect 12574 32510 12626 32562
rect 13358 32510 13410 32562
rect 13582 32510 13634 32562
rect 17278 32510 17330 32562
rect 17950 32510 18002 32562
rect 21422 32510 21474 32562
rect 21646 32510 21698 32562
rect 24334 32510 24386 32562
rect 25902 32510 25954 32562
rect 28030 32510 28082 32562
rect 28590 32510 28642 32562
rect 29374 32510 29426 32562
rect 29822 32510 29874 32562
rect 30718 32510 30770 32562
rect 32958 32510 33010 32562
rect 33518 32510 33570 32562
rect 36430 32510 36482 32562
rect 36990 32510 37042 32562
rect 37774 32510 37826 32562
rect 38334 32510 38386 32562
rect 38782 32510 38834 32562
rect 39566 32510 39618 32562
rect 42702 32510 42754 32562
rect 43150 32510 43202 32562
rect 44046 32510 44098 32562
rect 11566 32398 11618 32450
rect 20414 32398 20466 32450
rect 25342 32398 25394 32450
rect 26462 32398 26514 32450
rect 27694 32398 27746 32450
rect 32510 32398 32562 32450
rect 41806 32398 41858 32450
rect 16606 32286 16658 32338
rect 21310 32286 21362 32338
rect 24110 32286 24162 32338
rect 45166 32286 45218 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 26910 31950 26962 32002
rect 29822 31950 29874 32002
rect 12350 31838 12402 31890
rect 16158 31838 16210 31890
rect 21310 31838 21362 31890
rect 27806 31838 27858 31890
rect 37550 31838 37602 31890
rect 6974 31726 7026 31778
rect 7422 31726 7474 31778
rect 11342 31726 11394 31778
rect 11566 31726 11618 31778
rect 13582 31726 13634 31778
rect 15038 31726 15090 31778
rect 16606 31726 16658 31778
rect 16942 31726 16994 31778
rect 17614 31726 17666 31778
rect 18174 31726 18226 31778
rect 19294 31726 19346 31778
rect 19854 31726 19906 31778
rect 21758 31726 21810 31778
rect 22094 31738 22146 31790
rect 22766 31726 22818 31778
rect 23326 31726 23378 31778
rect 24334 31726 24386 31778
rect 25230 31726 25282 31778
rect 26126 31726 26178 31778
rect 26350 31726 26402 31778
rect 28366 31726 28418 31778
rect 29262 31726 29314 31778
rect 32062 31726 32114 31778
rect 32398 31726 32450 31778
rect 34638 31726 34690 31778
rect 38894 31726 38946 31778
rect 39678 31726 39730 31778
rect 3950 31614 4002 31666
rect 9662 31614 9714 31666
rect 11902 31614 11954 31666
rect 15374 31614 15426 31666
rect 15710 31614 15762 31666
rect 17166 31614 17218 31666
rect 20414 31614 20466 31666
rect 25454 31614 25506 31666
rect 26574 31614 26626 31666
rect 36206 31614 36258 31666
rect 39454 31614 39506 31666
rect 3838 31502 3890 31554
rect 10446 31502 10498 31554
rect 12798 31502 12850 31554
rect 13806 31502 13858 31554
rect 14478 31502 14530 31554
rect 14702 31502 14754 31554
rect 20750 31502 20802 31554
rect 22318 31502 22370 31554
rect 25566 31502 25618 31554
rect 40238 31502 40290 31554
rect 44942 31502 44994 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4846 31166 4898 31218
rect 5518 31166 5570 31218
rect 8206 31166 8258 31218
rect 18958 31166 19010 31218
rect 22430 31166 22482 31218
rect 29150 31166 29202 31218
rect 34302 31166 34354 31218
rect 41582 31166 41634 31218
rect 41918 31166 41970 31218
rect 8318 31054 8370 31106
rect 14702 31054 14754 31106
rect 15038 31054 15090 31106
rect 15710 31054 15762 31106
rect 16382 31054 16434 31106
rect 21646 31054 21698 31106
rect 26238 31054 26290 31106
rect 28814 31054 28866 31106
rect 34638 31054 34690 31106
rect 35870 31054 35922 31106
rect 36878 31054 36930 31106
rect 42254 31054 42306 31106
rect 43598 31054 43650 31106
rect 2046 30942 2098 30994
rect 2494 30942 2546 30994
rect 13470 30942 13522 30994
rect 15374 30942 15426 30994
rect 16046 30942 16098 30994
rect 20190 30942 20242 30994
rect 22206 30942 22258 30994
rect 22542 30942 22594 30994
rect 23438 30942 23490 30994
rect 25566 30942 25618 30994
rect 26126 30942 26178 30994
rect 26798 30942 26850 30994
rect 27358 30942 27410 30994
rect 28366 30942 28418 30994
rect 29486 30942 29538 30994
rect 34974 30942 35026 30994
rect 36206 30942 36258 30994
rect 36654 30942 36706 30994
rect 37550 30942 37602 30994
rect 37886 30942 37938 30994
rect 39006 30942 39058 30994
rect 39566 30942 39618 30994
rect 45054 30942 45106 30994
rect 12014 30830 12066 30882
rect 16830 30830 16882 30882
rect 17614 30830 17666 30882
rect 18510 30830 18562 30882
rect 20414 30830 20466 30882
rect 24558 30830 24610 30882
rect 25230 30830 25282 30882
rect 30718 30830 30770 30882
rect 33966 30830 34018 30882
rect 35534 30830 35586 30882
rect 39902 30830 39954 30882
rect 41022 30830 41074 30882
rect 43262 30830 43314 30882
rect 45726 30830 45778 30882
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 37438 30382 37490 30434
rect 14926 30270 14978 30322
rect 20414 30270 20466 30322
rect 3726 30158 3778 30210
rect 12126 30158 12178 30210
rect 12910 30158 12962 30210
rect 13470 30158 13522 30210
rect 14030 30158 14082 30210
rect 14590 30158 14642 30210
rect 19518 30158 19570 30210
rect 20078 30158 20130 30210
rect 22094 30158 22146 30210
rect 22542 30158 22594 30210
rect 23438 30158 23490 30210
rect 24334 30158 24386 30210
rect 25230 30158 25282 30210
rect 25790 30158 25842 30210
rect 26350 30158 26402 30210
rect 27134 30158 27186 30210
rect 28030 30158 28082 30210
rect 29150 30158 29202 30210
rect 29822 30158 29874 30210
rect 35534 30158 35586 30210
rect 37886 30158 37938 30210
rect 39342 30158 39394 30210
rect 40798 30158 40850 30210
rect 41022 30158 41074 30210
rect 41694 30158 41746 30210
rect 44270 30158 44322 30210
rect 45166 30158 45218 30210
rect 45838 30158 45890 30210
rect 3838 30046 3890 30098
rect 17166 30046 17218 30098
rect 21422 30046 21474 30098
rect 23102 30046 23154 30098
rect 24894 30046 24946 30098
rect 30270 30046 30322 30098
rect 33742 30046 33794 30098
rect 34078 30046 34130 30098
rect 34414 30046 34466 30098
rect 34750 30046 34802 30098
rect 35758 30046 35810 30098
rect 36318 30046 36370 30098
rect 38222 30046 38274 30098
rect 38670 30046 38722 30098
rect 42814 30046 42866 30098
rect 44830 30046 44882 30098
rect 45502 30046 45554 30098
rect 17838 29934 17890 29986
rect 19518 29934 19570 29986
rect 21758 29934 21810 29986
rect 25902 29934 25954 29986
rect 30606 29934 30658 29986
rect 33518 29934 33570 29986
rect 35198 29934 35250 29986
rect 37102 29934 37154 29986
rect 39006 29934 39058 29986
rect 42366 29934 42418 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4846 29598 4898 29650
rect 5406 29598 5458 29650
rect 5630 29598 5682 29650
rect 16494 29598 16546 29650
rect 17390 29598 17442 29650
rect 21198 29598 21250 29650
rect 23662 29598 23714 29650
rect 24110 29598 24162 29650
rect 25230 29598 25282 29650
rect 27358 29598 27410 29650
rect 27694 29598 27746 29650
rect 33182 29598 33234 29650
rect 45502 29598 45554 29650
rect 5966 29486 6018 29538
rect 17726 29486 17778 29538
rect 19518 29486 19570 29538
rect 27806 29486 27858 29538
rect 33518 29486 33570 29538
rect 34190 29486 34242 29538
rect 34750 29486 34802 29538
rect 38222 29486 38274 29538
rect 41918 29486 41970 29538
rect 42926 29486 42978 29538
rect 1822 29374 1874 29426
rect 2270 29374 2322 29426
rect 10782 29374 10834 29426
rect 16718 29374 16770 29426
rect 19182 29374 19234 29426
rect 20526 29374 20578 29426
rect 20862 29374 20914 29426
rect 23326 29374 23378 29426
rect 25790 29374 25842 29426
rect 26798 29374 26850 29426
rect 28590 29374 28642 29426
rect 29262 29374 29314 29426
rect 31502 29374 31554 29426
rect 31838 29374 31890 29426
rect 36766 29374 36818 29426
rect 37214 29374 37266 29426
rect 41022 29374 41074 29426
rect 41470 29374 41522 29426
rect 42254 29374 42306 29426
rect 42702 29374 42754 29426
rect 43598 29374 43650 29426
rect 43934 29374 43986 29426
rect 44942 29374 44994 29426
rect 12798 29262 12850 29314
rect 20078 29262 20130 29314
rect 21982 29262 22034 29314
rect 22990 29262 23042 29314
rect 24558 29262 24610 29314
rect 25566 29262 25618 29314
rect 31166 29262 31218 29314
rect 34638 29262 34690 29314
rect 37774 29262 37826 29314
rect 45950 29262 46002 29314
rect 18398 29150 18450 29202
rect 18734 29150 18786 29202
rect 30158 29150 30210 29202
rect 31278 29150 31330 29202
rect 36094 29150 36146 29202
rect 40126 29150 40178 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 9214 28814 9266 28866
rect 12014 28814 12066 28866
rect 14926 28814 14978 28866
rect 19630 28814 19682 28866
rect 28142 28814 28194 28866
rect 43598 28814 43650 28866
rect 45390 28814 45442 28866
rect 1934 28702 1986 28754
rect 18398 28702 18450 28754
rect 22654 28702 22706 28754
rect 28366 28702 28418 28754
rect 28590 28702 28642 28754
rect 32958 28702 33010 28754
rect 36430 28702 36482 28754
rect 42702 28702 42754 28754
rect 4286 28590 4338 28642
rect 4958 28590 5010 28642
rect 5630 28590 5682 28642
rect 11678 28590 11730 28642
rect 12686 28590 12738 28642
rect 14142 28590 14194 28642
rect 14590 28590 14642 28642
rect 19182 28590 19234 28642
rect 22206 28590 22258 28642
rect 23886 28590 23938 28642
rect 24558 28590 24610 28642
rect 25006 28590 25058 28642
rect 27694 28590 27746 28642
rect 29262 28590 29314 28642
rect 29710 28590 29762 28642
rect 30158 28590 30210 28642
rect 30830 28590 30882 28642
rect 31278 28590 31330 28642
rect 32286 28590 32338 28642
rect 32846 28590 32898 28642
rect 34526 28590 34578 28642
rect 35870 28590 35922 28642
rect 38446 28590 38498 28642
rect 40686 28590 40738 28642
rect 42478 28590 42530 28642
rect 43150 28590 43202 28642
rect 45614 28590 45666 28642
rect 5742 28478 5794 28530
rect 8542 28478 8594 28530
rect 8990 28478 9042 28530
rect 10110 28478 10162 28530
rect 12798 28478 12850 28530
rect 13918 28478 13970 28530
rect 16830 28478 16882 28530
rect 19070 28478 19122 28530
rect 21310 28478 21362 28530
rect 23102 28478 23154 28530
rect 24334 28478 24386 28530
rect 25342 28478 25394 28530
rect 33630 28478 33682 28530
rect 44158 28478 44210 28530
rect 44830 28478 44882 28530
rect 44942 28478 44994 28530
rect 45054 28478 45106 28530
rect 4622 28366 4674 28418
rect 7870 28366 7922 28418
rect 9550 28366 9602 28418
rect 9998 28366 10050 28418
rect 19966 28366 20018 28418
rect 21422 28366 21474 28418
rect 21646 28366 21698 28418
rect 22094 28366 22146 28418
rect 23214 28366 23266 28418
rect 23438 28366 23490 28418
rect 23662 28366 23714 28418
rect 30270 28366 30322 28418
rect 37438 28366 37490 28418
rect 39678 28366 39730 28418
rect 41806 28366 41858 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4734 28030 4786 28082
rect 5294 28030 5346 28082
rect 10222 28030 10274 28082
rect 13470 28030 13522 28082
rect 21086 28030 21138 28082
rect 23326 28030 23378 28082
rect 23998 28030 24050 28082
rect 25342 28030 25394 28082
rect 28814 28030 28866 28082
rect 33406 28030 33458 28082
rect 34974 28030 35026 28082
rect 6638 27918 6690 27970
rect 7758 27918 7810 27970
rect 9550 27918 9602 27970
rect 15822 27918 15874 27970
rect 17614 27918 17666 27970
rect 19070 27918 19122 27970
rect 19406 27918 19458 27970
rect 20974 27918 21026 27970
rect 21870 27918 21922 27970
rect 24334 27918 24386 27970
rect 25230 27918 25282 27970
rect 26014 27918 26066 27970
rect 26126 27918 26178 27970
rect 27134 27918 27186 27970
rect 27246 27918 27298 27970
rect 32174 27918 32226 27970
rect 33070 27918 33122 27970
rect 35310 27918 35362 27970
rect 36318 27918 36370 27970
rect 1710 27806 1762 27858
rect 2270 27806 2322 27858
rect 6750 27806 6802 27858
rect 7198 27806 7250 27858
rect 9774 27806 9826 27858
rect 10446 27806 10498 27858
rect 13246 27806 13298 27858
rect 13806 27806 13858 27858
rect 14030 27806 14082 27858
rect 17502 27806 17554 27858
rect 20190 27806 20242 27858
rect 20862 27806 20914 27858
rect 21758 27806 21810 27858
rect 23662 27806 23714 27858
rect 24670 27806 24722 27858
rect 25566 27806 25618 27858
rect 26910 27806 26962 27858
rect 28590 27806 28642 27858
rect 29822 27806 29874 27858
rect 32398 27806 32450 27858
rect 34302 27806 34354 27858
rect 34750 27806 34802 27858
rect 35758 27806 35810 27858
rect 36094 27806 36146 27858
rect 36766 27806 36818 27858
rect 37438 27806 37490 27858
rect 38334 27806 38386 27858
rect 40126 27806 40178 27858
rect 41022 27806 41074 27858
rect 41918 27806 41970 27858
rect 42926 27806 42978 27858
rect 44046 27806 44098 27858
rect 22878 27694 22930 27746
rect 31502 27694 31554 27746
rect 33854 27694 33906 27746
rect 39566 27694 39618 27746
rect 40014 27694 40066 27746
rect 42814 27694 42866 27746
rect 44494 27694 44546 27746
rect 8878 27582 8930 27634
rect 16606 27582 16658 27634
rect 18286 27582 18338 27634
rect 18622 27582 18674 27634
rect 26126 27582 26178 27634
rect 39118 27582 39170 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 11566 27246 11618 27298
rect 35422 27246 35474 27298
rect 37438 27246 37490 27298
rect 38334 27246 38386 27298
rect 1934 27134 1986 27186
rect 13806 27134 13858 27186
rect 14926 27134 14978 27186
rect 16494 27134 16546 27186
rect 17614 27134 17666 27186
rect 24334 27134 24386 27186
rect 24670 27134 24722 27186
rect 30382 27134 30434 27186
rect 30718 27134 30770 27186
rect 37214 27134 37266 27186
rect 39566 27134 39618 27186
rect 4286 27022 4338 27074
rect 7870 27022 7922 27074
rect 8094 27022 8146 27074
rect 11342 27022 11394 27074
rect 11678 27022 11730 27074
rect 14478 27022 14530 27074
rect 15486 27022 15538 27074
rect 17390 27022 17442 27074
rect 18734 27022 18786 27074
rect 19406 27022 19458 27074
rect 20526 27022 20578 27074
rect 21534 27022 21586 27074
rect 22206 27022 22258 27074
rect 23102 27022 23154 27074
rect 23998 27022 24050 27074
rect 24894 27022 24946 27074
rect 25342 27022 25394 27074
rect 25454 27022 25506 27074
rect 25790 27022 25842 27074
rect 26126 27022 26178 27074
rect 26350 27022 26402 27074
rect 28590 27022 28642 27074
rect 29374 27022 29426 27074
rect 29934 27022 29986 27074
rect 31166 27022 31218 27074
rect 31502 27022 31554 27074
rect 32174 27022 32226 27074
rect 32958 27022 33010 27074
rect 33854 27022 33906 27074
rect 34526 27022 34578 27074
rect 36094 27022 36146 27074
rect 37886 27022 37938 27074
rect 38222 27022 38274 27074
rect 38558 27022 38610 27074
rect 38894 27022 38946 27074
rect 40014 27022 40066 27074
rect 40350 27022 40402 27074
rect 41358 27022 41410 27074
rect 41806 27022 41858 27074
rect 42814 27022 42866 27074
rect 4622 26910 4674 26962
rect 4734 26910 4786 26962
rect 9998 26910 10050 26962
rect 11006 26910 11058 26962
rect 11118 26910 11170 26962
rect 14254 26910 14306 26962
rect 17054 26910 17106 26962
rect 18846 26910 18898 26962
rect 19294 26910 19346 26962
rect 21422 26910 21474 26962
rect 22094 26910 22146 26962
rect 26014 26910 26066 26962
rect 27582 26910 27634 26962
rect 28254 26910 28306 26962
rect 29150 26910 29202 26962
rect 31726 26910 31778 26962
rect 34302 26910 34354 26962
rect 36206 26910 36258 26962
rect 38110 26910 38162 26962
rect 39230 26910 39282 26962
rect 10670 26798 10722 26850
rect 16270 26798 16322 26850
rect 19182 26798 19234 26850
rect 22206 26798 22258 26850
rect 25230 26798 25282 26850
rect 27918 26798 27970 26850
rect 35086 26798 35138 26850
rect 40686 26798 40738 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 9662 26462 9714 26514
rect 19742 26462 19794 26514
rect 24110 26462 24162 26514
rect 24782 26462 24834 26514
rect 27470 26462 27522 26514
rect 28030 26462 28082 26514
rect 30270 26462 30322 26514
rect 33070 26462 33122 26514
rect 35758 26462 35810 26514
rect 36430 26462 36482 26514
rect 39678 26462 39730 26514
rect 43822 26462 43874 26514
rect 44158 26462 44210 26514
rect 5406 26350 5458 26402
rect 10222 26350 10274 26402
rect 10670 26350 10722 26402
rect 21310 26350 21362 26402
rect 21982 26350 22034 26402
rect 22430 26350 22482 26402
rect 24446 26350 24498 26402
rect 24558 26350 24610 26402
rect 26350 26350 26402 26402
rect 33742 26350 33794 26402
rect 2718 26238 2770 26290
rect 3166 26238 3218 26290
rect 6414 26238 6466 26290
rect 6974 26238 7026 26290
rect 8206 26238 8258 26290
rect 9998 26238 10050 26290
rect 11678 26238 11730 26290
rect 17502 26238 17554 26290
rect 17950 26238 18002 26290
rect 18622 26238 18674 26290
rect 18846 26238 18898 26290
rect 20190 26238 20242 26290
rect 20862 26238 20914 26290
rect 21758 26238 21810 26290
rect 22542 26238 22594 26290
rect 22990 26238 23042 26290
rect 23550 26238 23602 26290
rect 25230 26238 25282 26290
rect 25678 26238 25730 26290
rect 26798 26238 26850 26290
rect 27806 26238 27858 26290
rect 28366 26238 28418 26290
rect 29710 26238 29762 26290
rect 30158 26238 30210 26290
rect 30942 26238 30994 26290
rect 31278 26238 31330 26290
rect 32398 26238 32450 26290
rect 33294 26238 33346 26290
rect 33966 26238 34018 26290
rect 34862 26238 34914 26290
rect 37102 26238 37154 26290
rect 37774 26238 37826 26290
rect 38782 26238 38834 26290
rect 8654 26126 8706 26178
rect 11342 26126 11394 26178
rect 19406 26126 19458 26178
rect 26126 26126 26178 26178
rect 28926 26126 28978 26178
rect 29262 26126 29314 26178
rect 35198 26126 35250 26178
rect 36766 26126 36818 26178
rect 38222 26126 38274 26178
rect 39118 26126 39170 26178
rect 6190 26014 6242 26066
rect 8094 26014 8146 26066
rect 18510 26014 18562 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 1934 25678 1986 25730
rect 4622 25678 4674 25730
rect 26574 25678 26626 25730
rect 5854 25566 5906 25618
rect 12126 25566 12178 25618
rect 13694 25566 13746 25618
rect 16942 25566 16994 25618
rect 25006 25566 25058 25618
rect 31278 25566 31330 25618
rect 34862 25566 34914 25618
rect 37326 25566 37378 25618
rect 40126 25566 40178 25618
rect 45278 25566 45330 25618
rect 4286 25454 4338 25506
rect 7758 25454 7810 25506
rect 9214 25454 9266 25506
rect 14030 25454 14082 25506
rect 17614 25454 17666 25506
rect 18062 25454 18114 25506
rect 18510 25454 18562 25506
rect 19070 25454 19122 25506
rect 19406 25454 19458 25506
rect 19854 25454 19906 25506
rect 20526 25454 20578 25506
rect 21310 25454 21362 25506
rect 22318 25454 22370 25506
rect 23102 25454 23154 25506
rect 23774 25454 23826 25506
rect 24110 25454 24162 25506
rect 24558 25454 24610 25506
rect 25342 25454 25394 25506
rect 25566 25454 25618 25506
rect 26238 25454 26290 25506
rect 28254 25454 28306 25506
rect 30046 25454 30098 25506
rect 36430 25454 36482 25506
rect 40910 25454 40962 25506
rect 41358 25454 41410 25506
rect 42478 25454 42530 25506
rect 43486 25454 43538 25506
rect 44830 25454 44882 25506
rect 4734 25342 4786 25394
rect 8542 25342 8594 25394
rect 8878 25342 8930 25394
rect 9998 25342 10050 25394
rect 12462 25342 12514 25394
rect 14814 25342 14866 25394
rect 17726 25342 17778 25394
rect 20414 25342 20466 25394
rect 22430 25342 22482 25394
rect 23438 25342 23490 25394
rect 25902 25342 25954 25394
rect 27918 25342 27970 25394
rect 40462 25342 40514 25394
rect 41918 25342 41970 25394
rect 12798 25230 12850 25282
rect 21198 25230 21250 25282
rect 23998 25230 24050 25282
rect 25454 25230 25506 25282
rect 26462 25230 26514 25282
rect 26910 25230 26962 25282
rect 27246 25230 27298 25282
rect 27582 25230 27634 25282
rect 28590 25230 28642 25282
rect 37774 25230 37826 25282
rect 38110 25230 38162 25282
rect 38446 25230 38498 25282
rect 38782 25230 38834 25282
rect 39118 25230 39170 25282
rect 39678 25230 39730 25282
rect 41470 25230 41522 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 6638 24894 6690 24946
rect 10110 24894 10162 24946
rect 10782 24894 10834 24946
rect 12462 24894 12514 24946
rect 19182 24894 19234 24946
rect 32286 24894 32338 24946
rect 33630 24894 33682 24946
rect 35198 24894 35250 24946
rect 5070 24782 5122 24834
rect 6974 24782 7026 24834
rect 8430 24782 8482 24834
rect 8878 24782 8930 24834
rect 9550 24782 9602 24834
rect 11342 24782 11394 24834
rect 11790 24782 11842 24834
rect 12350 24782 12402 24834
rect 13358 24782 13410 24834
rect 19742 24782 19794 24834
rect 20190 24782 20242 24834
rect 22878 24782 22930 24834
rect 26350 24782 26402 24834
rect 27470 24782 27522 24834
rect 29262 24782 29314 24834
rect 35646 24782 35698 24834
rect 39678 24782 39730 24834
rect 40238 24782 40290 24834
rect 41918 24782 41970 24834
rect 44494 24782 44546 24834
rect 2270 24670 2322 24722
rect 2718 24670 2770 24722
rect 6414 24670 6466 24722
rect 7310 24670 7362 24722
rect 7758 24670 7810 24722
rect 8094 24670 8146 24722
rect 11118 24670 11170 24722
rect 12574 24670 12626 24722
rect 13022 24670 13074 24722
rect 13246 24670 13298 24722
rect 16718 24670 16770 24722
rect 17838 24670 17890 24722
rect 18622 24670 18674 24722
rect 19518 24670 19570 24722
rect 20526 24670 20578 24722
rect 20974 24670 21026 24722
rect 21870 24670 21922 24722
rect 22542 24670 22594 24722
rect 23886 24670 23938 24722
rect 24222 24670 24274 24722
rect 25678 24670 25730 24722
rect 26126 24670 26178 24722
rect 26798 24670 26850 24722
rect 27134 24670 27186 24722
rect 30046 24670 30098 24722
rect 31726 24670 31778 24722
rect 34526 24670 34578 24722
rect 34974 24670 35026 24722
rect 36318 24670 36370 24722
rect 37214 24670 37266 24722
rect 38334 24670 38386 24722
rect 39454 24670 39506 24722
rect 41246 24670 41298 24722
rect 41806 24670 41858 24722
rect 42590 24670 42642 24722
rect 42926 24670 42978 24722
rect 44046 24670 44098 24722
rect 44718 24670 44770 24722
rect 45502 24670 45554 24722
rect 45726 24670 45778 24722
rect 1822 24558 1874 24610
rect 5854 24558 5906 24610
rect 18174 24558 18226 24610
rect 22206 24558 22258 24610
rect 22318 24558 22370 24610
rect 23998 24558 24050 24610
rect 26014 24558 26066 24610
rect 33070 24558 33122 24610
rect 34190 24558 34242 24610
rect 37886 24558 37938 24610
rect 39118 24558 39170 24610
rect 40910 24558 40962 24610
rect 1934 24446 1986 24498
rect 16830 24446 16882 24498
rect 23550 24446 23602 24498
rect 27134 24446 27186 24498
rect 44830 24446 44882 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 2830 24110 2882 24162
rect 30606 24110 30658 24162
rect 38446 24110 38498 24162
rect 14590 23998 14642 24050
rect 15374 23998 15426 24050
rect 18622 23998 18674 24050
rect 19294 23998 19346 24050
rect 27806 23998 27858 24050
rect 28366 23998 28418 24050
rect 29598 23998 29650 24050
rect 31838 23998 31890 24050
rect 37214 23998 37266 24050
rect 41918 23998 41970 24050
rect 45278 23998 45330 24050
rect 4286 23886 4338 23938
rect 4958 23886 5010 23938
rect 5630 23886 5682 23938
rect 10110 23886 10162 23938
rect 10558 23886 10610 23938
rect 11902 23886 11954 23938
rect 12798 23886 12850 23938
rect 14478 23886 14530 23938
rect 14702 23886 14754 23938
rect 15710 23886 15762 23938
rect 19630 23886 19682 23938
rect 20190 23886 20242 23938
rect 20750 23886 20802 23938
rect 21982 23886 22034 23938
rect 22654 23886 22706 23938
rect 23326 23886 23378 23938
rect 24334 23886 24386 23938
rect 25006 23886 25058 23938
rect 25342 23886 25394 23938
rect 26462 23886 26514 23938
rect 26798 23886 26850 23938
rect 27470 23886 27522 23938
rect 29822 23886 29874 23938
rect 29934 23886 29986 23938
rect 30382 23886 30434 23938
rect 31054 23886 31106 23938
rect 32286 23886 32338 23938
rect 33630 23886 33682 23938
rect 33966 23886 34018 23938
rect 34862 23886 34914 23938
rect 35422 23886 35474 23938
rect 36206 23886 36258 23938
rect 37438 23886 37490 23938
rect 37774 23886 37826 23938
rect 38782 23886 38834 23938
rect 40462 23886 40514 23938
rect 41134 23886 41186 23938
rect 42590 23886 42642 23938
rect 43038 23886 43090 23938
rect 44158 23886 44210 23938
rect 44830 23886 44882 23938
rect 45950 23886 46002 23938
rect 8654 23774 8706 23826
rect 9662 23774 9714 23826
rect 11118 23774 11170 23826
rect 14142 23774 14194 23826
rect 16494 23774 16546 23826
rect 19294 23774 19346 23826
rect 22878 23774 22930 23826
rect 23662 23774 23714 23826
rect 24558 23774 24610 23826
rect 25790 23774 25842 23826
rect 26350 23774 26402 23826
rect 32622 23774 32674 23826
rect 33182 23774 33234 23826
rect 34190 23774 34242 23826
rect 36990 23774 37042 23826
rect 39006 23774 39058 23826
rect 40798 23774 40850 23826
rect 4734 23662 4786 23714
rect 6638 23662 6690 23714
rect 8542 23662 8594 23714
rect 10670 23662 10722 23714
rect 21422 23662 21474 23714
rect 27134 23662 27186 23714
rect 27694 23662 27746 23714
rect 29374 23662 29426 23714
rect 31390 23662 31442 23714
rect 37214 23662 37266 23714
rect 41582 23662 41634 23714
rect 45726 23662 45778 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 4846 23326 4898 23378
rect 5854 23326 5906 23378
rect 7646 23326 7698 23378
rect 14926 23326 14978 23378
rect 15934 23326 15986 23378
rect 20750 23326 20802 23378
rect 23998 23326 24050 23378
rect 26462 23326 26514 23378
rect 27470 23326 27522 23378
rect 27918 23326 27970 23378
rect 31838 23326 31890 23378
rect 32286 23326 32338 23378
rect 42030 23326 42082 23378
rect 6974 23214 7026 23266
rect 8766 23214 8818 23266
rect 9662 23214 9714 23266
rect 10670 23214 10722 23266
rect 16606 23214 16658 23266
rect 23550 23214 23602 23266
rect 24558 23214 24610 23266
rect 25678 23214 25730 23266
rect 29038 23214 29090 23266
rect 30606 23214 30658 23266
rect 31054 23214 31106 23266
rect 31502 23214 31554 23266
rect 44494 23214 44546 23266
rect 1934 23102 1986 23154
rect 2382 23102 2434 23154
rect 5518 23102 5570 23154
rect 6190 23102 6242 23154
rect 6862 23102 6914 23154
rect 7982 23102 8034 23154
rect 8430 23102 8482 23154
rect 10110 23102 10162 23154
rect 10446 23102 10498 23154
rect 11118 23102 11170 23154
rect 11902 23102 11954 23154
rect 12798 23102 12850 23154
rect 14142 23102 14194 23154
rect 14814 23102 14866 23154
rect 15598 23102 15650 23154
rect 16382 23102 16434 23154
rect 17390 23102 17442 23154
rect 21198 23102 21250 23154
rect 21422 23102 21474 23154
rect 22542 23102 22594 23154
rect 23438 23102 23490 23154
rect 24222 23102 24274 23154
rect 25230 23102 25282 23154
rect 25902 23102 25954 23154
rect 26238 23102 26290 23154
rect 26798 23102 26850 23154
rect 27246 23102 27298 23154
rect 28702 23102 28754 23154
rect 33518 23102 33570 23154
rect 33854 23102 33906 23154
rect 34974 23102 35026 23154
rect 35758 23102 35810 23154
rect 36206 23102 36258 23154
rect 39006 23102 39058 23154
rect 42590 23102 42642 23154
rect 44942 23102 44994 23154
rect 45502 23102 45554 23154
rect 14478 22990 14530 23042
rect 18174 22990 18226 23042
rect 20302 22990 20354 23042
rect 21534 22990 21586 23042
rect 25790 22990 25842 23042
rect 26350 22990 26402 23042
rect 28366 22990 28418 23042
rect 33182 22990 33234 23042
rect 38558 22990 38610 23042
rect 14926 22878 14978 22930
rect 29486 22878 29538 22930
rect 30270 22878 30322 22930
rect 36430 22878 36482 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 9550 22542 9602 22594
rect 9886 22542 9938 22594
rect 13806 22542 13858 22594
rect 32398 22542 32450 22594
rect 37102 22542 37154 22594
rect 37438 22542 37490 22594
rect 2046 22430 2098 22482
rect 11678 22430 11730 22482
rect 13694 22430 13746 22482
rect 14590 22430 14642 22482
rect 15710 22430 15762 22482
rect 19294 22430 19346 22482
rect 20526 22430 20578 22482
rect 25902 22430 25954 22482
rect 30606 22430 30658 22482
rect 39790 22430 39842 22482
rect 41358 22430 41410 22482
rect 4286 22318 4338 22370
rect 4734 22318 4786 22370
rect 5966 22318 6018 22370
rect 6302 22318 6354 22370
rect 6862 22318 6914 22370
rect 7870 22318 7922 22370
rect 8430 22318 8482 22370
rect 10446 22318 10498 22370
rect 12238 22318 12290 22370
rect 15038 22318 15090 22370
rect 15374 22318 15426 22370
rect 15822 22318 15874 22370
rect 16382 22318 16434 22370
rect 19966 22318 20018 22370
rect 21422 22318 21474 22370
rect 21870 22318 21922 22370
rect 22654 22318 22706 22370
rect 23214 22318 23266 22370
rect 24222 22318 24274 22370
rect 26686 22318 26738 22370
rect 27022 22318 27074 22370
rect 27582 22318 27634 22370
rect 29262 22318 29314 22370
rect 32286 22318 32338 22370
rect 32622 22318 32674 22370
rect 33406 22318 33458 22370
rect 33518 22318 33570 22370
rect 34302 22318 34354 22370
rect 40238 22318 40290 22370
rect 42142 22318 42194 22370
rect 42478 22318 42530 22370
rect 43486 22318 43538 22370
rect 5070 22206 5122 22258
rect 7086 22206 7138 22258
rect 10558 22206 10610 22258
rect 16046 22206 16098 22258
rect 17166 22206 17218 22258
rect 23438 22206 23490 22258
rect 24334 22206 24386 22258
rect 25342 22206 25394 22258
rect 26126 22206 26178 22258
rect 27918 22206 27970 22258
rect 31166 22206 31218 22258
rect 34526 22206 34578 22258
rect 35198 22206 35250 22258
rect 37662 22206 37714 22258
rect 38222 22206 38274 22258
rect 7534 22094 7586 22146
rect 8206 22094 8258 22146
rect 11902 22094 11954 22146
rect 13022 22094 13074 22146
rect 13582 22094 13634 22146
rect 15598 22094 15650 22146
rect 21310 22094 21362 22146
rect 21534 22094 21586 22146
rect 23326 22094 23378 22146
rect 25006 22094 25058 22146
rect 25902 22094 25954 22146
rect 27134 22094 27186 22146
rect 27246 22094 27298 22146
rect 28254 22094 28306 22146
rect 28590 22094 28642 22146
rect 31278 22094 31330 22146
rect 34862 22094 34914 22146
rect 35646 22094 35698 22146
rect 40574 22094 40626 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 4846 21758 4898 21810
rect 5630 21758 5682 21810
rect 6302 21758 6354 21810
rect 8094 21758 8146 21810
rect 11566 21758 11618 21810
rect 12238 21758 12290 21810
rect 13806 21758 13858 21810
rect 15038 21758 15090 21810
rect 15150 21758 15202 21810
rect 16046 21758 16098 21810
rect 19966 21758 20018 21810
rect 20414 21758 20466 21810
rect 21982 21758 22034 21810
rect 22094 21758 22146 21810
rect 22318 21758 22370 21810
rect 22654 21758 22706 21810
rect 24334 21758 24386 21810
rect 26126 21758 26178 21810
rect 26238 21758 26290 21810
rect 26798 21758 26850 21810
rect 27806 21758 27858 21810
rect 28478 21758 28530 21810
rect 34750 21758 34802 21810
rect 36766 21758 36818 21810
rect 37998 21758 38050 21810
rect 6862 21646 6914 21698
rect 7422 21646 7474 21698
rect 11230 21646 11282 21698
rect 11902 21646 11954 21698
rect 13134 21646 13186 21698
rect 13470 21646 13522 21698
rect 16830 21646 16882 21698
rect 17614 21646 17666 21698
rect 20526 21646 20578 21698
rect 24670 21646 24722 21698
rect 28030 21646 28082 21698
rect 29262 21646 29314 21698
rect 30270 21646 30322 21698
rect 35982 21646 36034 21698
rect 41134 21646 41186 21698
rect 41470 21646 41522 21698
rect 45166 21646 45218 21698
rect 2158 21534 2210 21586
rect 2494 21534 2546 21586
rect 10670 21534 10722 21586
rect 11006 21534 11058 21586
rect 12574 21534 12626 21586
rect 14814 21534 14866 21586
rect 14926 21534 14978 21586
rect 15374 21534 15426 21586
rect 15710 21534 15762 21586
rect 15934 21534 15986 21586
rect 16158 21534 16210 21586
rect 16382 21534 16434 21586
rect 17502 21534 17554 21586
rect 19406 21534 19458 21586
rect 20302 21534 20354 21586
rect 20974 21534 21026 21586
rect 21870 21534 21922 21586
rect 23102 21534 23154 21586
rect 23438 21534 23490 21586
rect 27022 21534 27074 21586
rect 27246 21534 27298 21586
rect 29710 21534 29762 21586
rect 30046 21534 30098 21586
rect 30942 21534 30994 21586
rect 31502 21534 31554 21586
rect 32398 21534 32450 21586
rect 32958 21534 33010 21586
rect 33294 21534 33346 21586
rect 33742 21534 33794 21586
rect 35086 21534 35138 21586
rect 36206 21534 36258 21586
rect 37662 21534 37714 21586
rect 42478 21534 42530 21586
rect 43598 21534 43650 21586
rect 44718 21534 44770 21586
rect 14366 21422 14418 21474
rect 18062 21422 18114 21474
rect 23214 21422 23266 21474
rect 27134 21422 27186 21474
rect 27694 21422 27746 21474
rect 28366 21422 28418 21474
rect 35534 21422 35586 21474
rect 41918 21422 41970 21474
rect 6638 21310 6690 21362
rect 26350 21310 26402 21362
rect 28702 21310 28754 21362
rect 43374 21310 43426 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 13582 20974 13634 21026
rect 22654 20974 22706 21026
rect 27806 20974 27858 21026
rect 33742 20974 33794 21026
rect 2718 20862 2770 20914
rect 10558 20862 10610 20914
rect 11342 20862 11394 20914
rect 13918 20862 13970 20914
rect 20302 20862 20354 20914
rect 27358 20862 27410 20914
rect 28590 20862 28642 20914
rect 29710 20862 29762 20914
rect 35198 20862 35250 20914
rect 41134 20862 41186 20914
rect 4286 20750 4338 20802
rect 6302 20750 6354 20802
rect 6862 20750 6914 20802
rect 7646 20750 7698 20802
rect 12126 20750 12178 20802
rect 16830 20750 16882 20802
rect 17166 20750 17218 20802
rect 17838 20750 17890 20802
rect 20414 20750 20466 20802
rect 20862 20750 20914 20802
rect 22990 20750 23042 20802
rect 27134 20750 27186 20802
rect 27806 20750 27858 20802
rect 29262 20750 29314 20802
rect 30494 20750 30546 20802
rect 30942 20750 30994 20802
rect 32398 20750 32450 20802
rect 33294 20750 33346 20802
rect 33854 20750 33906 20802
rect 34414 20750 34466 20802
rect 34526 20750 34578 20802
rect 34638 20750 34690 20802
rect 35646 20750 35698 20802
rect 37998 20750 38050 20802
rect 39118 20750 39170 20802
rect 42702 20750 42754 20802
rect 8430 20638 8482 20690
rect 12014 20638 12066 20690
rect 12910 20638 12962 20690
rect 13470 20638 13522 20690
rect 16046 20638 16098 20690
rect 17278 20638 17330 20690
rect 23214 20638 23266 20690
rect 23774 20638 23826 20690
rect 27470 20638 27522 20690
rect 28142 20638 28194 20690
rect 30158 20638 30210 20690
rect 31166 20638 31218 20690
rect 31614 20638 31666 20690
rect 34078 20638 34130 20690
rect 35982 20638 36034 20690
rect 36318 20638 36370 20690
rect 36990 20638 37042 20690
rect 39230 20638 39282 20690
rect 42142 20638 42194 20690
rect 4734 20526 4786 20578
rect 5070 20526 5122 20578
rect 5966 20526 6018 20578
rect 6638 20526 6690 20578
rect 11006 20526 11058 20578
rect 12574 20526 12626 20578
rect 17390 20526 17442 20578
rect 20190 20526 20242 20578
rect 24334 20526 24386 20578
rect 38110 20526 38162 20578
rect 42478 20526 42530 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 6078 20190 6130 20242
rect 9550 20190 9602 20242
rect 23102 20190 23154 20242
rect 24446 20190 24498 20242
rect 30830 20190 30882 20242
rect 1710 20078 1762 20130
rect 2046 20078 2098 20130
rect 5294 20078 5346 20130
rect 8542 20078 8594 20130
rect 9886 20078 9938 20130
rect 10670 20078 10722 20130
rect 11678 20078 11730 20130
rect 12014 20078 12066 20130
rect 14030 20078 14082 20130
rect 15262 20078 15314 20130
rect 17390 20078 17442 20130
rect 22542 20078 22594 20130
rect 23774 20078 23826 20130
rect 24110 20078 24162 20130
rect 28702 20078 28754 20130
rect 29598 20078 29650 20130
rect 33518 20078 33570 20130
rect 36094 20078 36146 20130
rect 39902 20078 39954 20130
rect 41806 20078 41858 20130
rect 42814 20078 42866 20130
rect 43262 20078 43314 20130
rect 2382 19966 2434 20018
rect 2942 19966 2994 20018
rect 6414 19966 6466 20018
rect 8878 19966 8930 20018
rect 10446 19966 10498 20018
rect 11454 19966 11506 20018
rect 12798 19966 12850 20018
rect 13470 19966 13522 20018
rect 16718 19966 16770 20018
rect 17614 19966 17666 20018
rect 18174 19966 18226 20018
rect 18622 19966 18674 20018
rect 19854 19966 19906 20018
rect 28366 19966 28418 20018
rect 29262 19966 29314 20018
rect 31726 19966 31778 20018
rect 32510 19966 32562 20018
rect 33182 19966 33234 20018
rect 34526 19966 34578 20018
rect 35086 19966 35138 20018
rect 35534 19966 35586 20018
rect 35982 19966 36034 20018
rect 36766 19966 36818 20018
rect 37102 19966 37154 20018
rect 38110 19966 38162 20018
rect 39230 19966 39282 20018
rect 39566 19966 39618 20018
rect 41022 19966 41074 20018
rect 42142 19966 42194 20018
rect 42702 19966 42754 20018
rect 44046 19966 44098 20018
rect 44942 19966 44994 20018
rect 13582 19854 13634 19906
rect 19630 19854 19682 19906
rect 24558 19854 24610 19906
rect 32062 19854 32114 19906
rect 38782 19854 38834 19906
rect 40350 19854 40402 19906
rect 41358 19854 41410 19906
rect 11118 19742 11170 19794
rect 18062 19742 18114 19794
rect 18510 19742 18562 19794
rect 20302 19742 20354 19794
rect 33966 19742 34018 19794
rect 34190 19742 34242 19794
rect 34638 19742 34690 19794
rect 34750 19742 34802 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 4510 19406 4562 19458
rect 10558 19406 10610 19458
rect 10894 19406 10946 19458
rect 15710 19406 15762 19458
rect 44046 19406 44098 19458
rect 3166 19294 3218 19346
rect 4622 19294 4674 19346
rect 7982 19294 8034 19346
rect 10110 19294 10162 19346
rect 14478 19294 14530 19346
rect 15598 19294 15650 19346
rect 20078 19294 20130 19346
rect 21758 19294 21810 19346
rect 33518 19294 33570 19346
rect 36990 19294 37042 19346
rect 1822 19182 1874 19234
rect 2270 19182 2322 19234
rect 3502 19182 3554 19234
rect 5630 19182 5682 19234
rect 7198 19182 7250 19234
rect 11342 19182 11394 19234
rect 12350 19182 12402 19234
rect 13470 19182 13522 19234
rect 14030 19182 14082 19234
rect 15934 19182 15986 19234
rect 16606 19182 16658 19234
rect 17166 19182 17218 19234
rect 23214 19182 23266 19234
rect 29374 19182 29426 19234
rect 32734 19182 32786 19234
rect 35086 19182 35138 19234
rect 35646 19182 35698 19234
rect 36094 19182 36146 19234
rect 37438 19182 37490 19234
rect 37886 19182 37938 19234
rect 38894 19182 38946 19234
rect 39342 19182 39394 19234
rect 39790 19182 39842 19234
rect 2606 19070 2658 19122
rect 5070 19070 5122 19122
rect 6638 19070 6690 19122
rect 11678 19070 11730 19122
rect 16270 19070 16322 19122
rect 16718 19070 16770 19122
rect 16830 19070 16882 19122
rect 17950 19070 18002 19122
rect 24558 19070 24610 19122
rect 29710 19070 29762 19122
rect 34526 19070 34578 19122
rect 36430 19070 36482 19122
rect 42590 19070 42642 19122
rect 3838 18958 3890 19010
rect 4958 18958 5010 19010
rect 6190 18958 6242 19010
rect 12910 18958 12962 19010
rect 13806 18958 13858 19010
rect 21646 18958 21698 19010
rect 32174 18958 32226 19010
rect 33070 18958 33122 19010
rect 34078 18958 34130 19010
rect 36542 18958 36594 19010
rect 38222 18958 38274 19010
rect 38670 18958 38722 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 12798 18622 12850 18674
rect 13022 18622 13074 18674
rect 14030 18622 14082 18674
rect 14254 18622 14306 18674
rect 41582 18622 41634 18674
rect 5630 18510 5682 18562
rect 8318 18510 8370 18562
rect 8990 18510 9042 18562
rect 18398 18510 18450 18562
rect 18510 18510 18562 18562
rect 24558 18510 24610 18562
rect 29710 18510 29762 18562
rect 30382 18510 30434 18562
rect 31950 18510 32002 18562
rect 38894 18510 38946 18562
rect 41358 18510 41410 18562
rect 45054 18510 45106 18562
rect 1710 18398 1762 18450
rect 2942 18398 2994 18450
rect 3390 18398 3442 18450
rect 8094 18398 8146 18450
rect 8766 18398 8818 18450
rect 9550 18398 9602 18450
rect 10334 18398 10386 18450
rect 13358 18398 13410 18450
rect 14702 18398 14754 18450
rect 15486 18398 15538 18450
rect 15934 18398 15986 18450
rect 16382 18398 16434 18450
rect 17390 18398 17442 18450
rect 18174 18398 18226 18450
rect 19182 18398 19234 18450
rect 19742 18398 19794 18450
rect 20526 18398 20578 18450
rect 22654 18398 22706 18450
rect 23438 18398 23490 18450
rect 24222 18398 24274 18450
rect 29486 18398 29538 18450
rect 30158 18398 30210 18450
rect 34638 18398 34690 18450
rect 35422 18398 35474 18450
rect 36654 18398 36706 18450
rect 38334 18398 38386 18450
rect 39454 18398 39506 18450
rect 42030 18398 42082 18450
rect 42478 18398 42530 18450
rect 45950 18398 46002 18450
rect 2270 18286 2322 18338
rect 12462 18286 12514 18338
rect 12910 18286 12962 18338
rect 14142 18286 14194 18338
rect 15038 18286 15090 18338
rect 16830 18286 16882 18338
rect 17950 18286 18002 18338
rect 21758 18286 21810 18338
rect 25342 18286 25394 18338
rect 31726 18286 31778 18338
rect 32510 18286 32562 18338
rect 34750 18286 34802 18338
rect 35982 18286 36034 18338
rect 37438 18286 37490 18338
rect 6414 18174 6466 18226
rect 23774 18174 23826 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 4062 17838 4114 17890
rect 4958 17838 5010 17890
rect 10670 17838 10722 17890
rect 11006 17838 11058 17890
rect 23774 17838 23826 17890
rect 34414 17838 34466 17890
rect 36318 17838 36370 17890
rect 36542 17838 36594 17890
rect 42590 17838 42642 17890
rect 3278 17726 3330 17778
rect 4174 17726 4226 17778
rect 4622 17726 4674 17778
rect 5070 17726 5122 17778
rect 9662 17726 9714 17778
rect 14814 17726 14866 17778
rect 16942 17726 16994 17778
rect 17950 17726 18002 17778
rect 18622 17726 18674 17778
rect 19854 17726 19906 17778
rect 21982 17726 22034 17778
rect 29374 17726 29426 17778
rect 34974 17726 35026 17778
rect 35870 17726 35922 17778
rect 37438 17726 37490 17778
rect 37886 17726 37938 17778
rect 1710 17614 1762 17666
rect 3502 17614 3554 17666
rect 5518 17614 5570 17666
rect 6078 17614 6130 17666
rect 12462 17614 12514 17666
rect 12910 17614 12962 17666
rect 13358 17614 13410 17666
rect 13694 17614 13746 17666
rect 14030 17614 14082 17666
rect 18958 17614 19010 17666
rect 19518 17614 19570 17666
rect 20414 17614 20466 17666
rect 20638 17614 20690 17666
rect 21422 17614 21474 17666
rect 21646 17614 21698 17666
rect 23214 17614 23266 17666
rect 29822 17614 29874 17666
rect 31278 17614 31330 17666
rect 31726 17614 31778 17666
rect 34078 17614 34130 17666
rect 35422 17614 35474 17666
rect 38446 17614 38498 17666
rect 2382 17502 2434 17554
rect 3614 17502 3666 17554
rect 9214 17502 9266 17554
rect 9886 17502 9938 17554
rect 10222 17502 10274 17554
rect 11342 17502 11394 17554
rect 11566 17502 11618 17554
rect 13582 17502 13634 17554
rect 20078 17502 20130 17554
rect 21982 17502 22034 17554
rect 22206 17502 22258 17554
rect 22878 17502 22930 17554
rect 28254 17502 28306 17554
rect 28590 17502 28642 17554
rect 36430 17502 36482 17554
rect 36990 17502 37042 17554
rect 39118 17502 39170 17554
rect 2046 17390 2098 17442
rect 2718 17390 2770 17442
rect 8430 17390 8482 17442
rect 17390 17390 17442 17442
rect 20750 17390 20802 17442
rect 22542 17390 22594 17442
rect 29598 17390 29650 17442
rect 30942 17390 30994 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 4734 17054 4786 17106
rect 5294 17054 5346 17106
rect 8430 17054 8482 17106
rect 12686 17054 12738 17106
rect 13022 17054 13074 17106
rect 18062 17054 18114 17106
rect 23102 17054 23154 17106
rect 23886 17054 23938 17106
rect 24670 17054 24722 17106
rect 35982 17054 36034 17106
rect 37550 17054 37602 17106
rect 38558 17054 38610 17106
rect 40014 17054 40066 17106
rect 9662 16942 9714 16994
rect 9998 16942 10050 16994
rect 10670 16942 10722 16994
rect 12126 16942 12178 16994
rect 15710 16942 15762 16994
rect 19630 16942 19682 16994
rect 23326 16942 23378 16994
rect 28478 16942 28530 16994
rect 33294 16942 33346 16994
rect 36318 16942 36370 16994
rect 38894 16942 38946 16994
rect 39678 16942 39730 16994
rect 1710 16830 1762 16882
rect 2158 16830 2210 16882
rect 5406 16830 5458 16882
rect 5966 16830 6018 16882
rect 9102 16830 9154 16882
rect 10446 16830 10498 16882
rect 12238 16830 12290 16882
rect 16382 16830 16434 16882
rect 17502 16830 17554 16882
rect 21870 16830 21922 16882
rect 22766 16830 22818 16882
rect 26126 16830 26178 16882
rect 26350 16830 26402 16882
rect 28366 16830 28418 16882
rect 30270 16830 30322 16882
rect 33182 16830 33234 16882
rect 34750 16830 34802 16882
rect 35758 16830 35810 16882
rect 36542 16830 36594 16882
rect 39454 16830 39506 16882
rect 43486 16830 43538 16882
rect 44382 16830 44434 16882
rect 11454 16718 11506 16770
rect 13582 16718 13634 16770
rect 18734 16718 18786 16770
rect 22990 16718 23042 16770
rect 23774 16718 23826 16770
rect 26798 16718 26850 16770
rect 27246 16718 27298 16770
rect 32286 16718 32338 16770
rect 35198 16718 35250 16770
rect 45502 16718 45554 16770
rect 11118 16606 11170 16658
rect 21534 16606 21586 16658
rect 23662 16606 23714 16658
rect 25678 16606 25730 16658
rect 25902 16606 25954 16658
rect 26238 16606 26290 16658
rect 26574 16606 26626 16658
rect 31502 16606 31554 16658
rect 33966 16606 34018 16658
rect 34302 16606 34354 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 3502 16270 3554 16322
rect 14366 16270 14418 16322
rect 16606 16270 16658 16322
rect 20190 16270 20242 16322
rect 1822 16158 1874 16210
rect 2270 16158 2322 16210
rect 2718 16158 2770 16210
rect 6078 16158 6130 16210
rect 8990 16158 9042 16210
rect 11118 16158 11170 16210
rect 11902 16158 11954 16210
rect 15262 16158 15314 16210
rect 23662 16158 23714 16210
rect 25454 16158 25506 16210
rect 29262 16158 29314 16210
rect 30046 16158 30098 16210
rect 31726 16158 31778 16210
rect 35758 16158 35810 16210
rect 39006 16158 39058 16210
rect 8318 16046 8370 16098
rect 12350 16046 12402 16098
rect 13806 16046 13858 16098
rect 16270 16046 16322 16098
rect 19742 16046 19794 16098
rect 19966 16046 20018 16098
rect 20302 16046 20354 16098
rect 21646 16046 21698 16098
rect 25006 16046 25058 16098
rect 25902 16046 25954 16098
rect 26014 16046 26066 16098
rect 26910 16046 26962 16098
rect 27358 16046 27410 16098
rect 28030 16046 28082 16098
rect 28590 16046 28642 16098
rect 29710 16046 29762 16098
rect 30606 16046 30658 16098
rect 31278 16046 31330 16098
rect 32174 16046 32226 16098
rect 32510 16046 32562 16098
rect 33742 16046 33794 16098
rect 34862 16046 34914 16098
rect 35422 16046 35474 16098
rect 38222 16046 38274 16098
rect 39454 16046 39506 16098
rect 40126 16046 40178 16098
rect 40686 16046 40738 16098
rect 41246 16046 41298 16098
rect 41918 16046 41970 16098
rect 42926 16046 42978 16098
rect 43598 16046 43650 16098
rect 3614 15934 3666 15986
rect 12686 15934 12738 15986
rect 13582 15934 13634 15986
rect 15934 15934 15986 15986
rect 18622 15934 18674 15986
rect 25342 15934 25394 15986
rect 30942 15934 30994 15986
rect 32734 15934 32786 15986
rect 33182 15934 33234 15986
rect 38558 15934 38610 15986
rect 39790 15934 39842 15986
rect 43374 15934 43426 15986
rect 5966 15822 6018 15874
rect 11566 15822 11618 15874
rect 14702 15822 14754 15874
rect 20526 15822 20578 15874
rect 24334 15822 24386 15874
rect 40798 15822 40850 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 7982 15486 8034 15538
rect 9102 15486 9154 15538
rect 11566 15486 11618 15538
rect 12238 15486 12290 15538
rect 13134 15486 13186 15538
rect 16830 15486 16882 15538
rect 20302 15486 20354 15538
rect 21870 15486 21922 15538
rect 22430 15486 22482 15538
rect 23326 15486 23378 15538
rect 24110 15486 24162 15538
rect 25566 15486 25618 15538
rect 31054 15486 31106 15538
rect 32398 15486 32450 15538
rect 37326 15486 37378 15538
rect 37662 15486 37714 15538
rect 40014 15486 40066 15538
rect 4286 15374 4338 15426
rect 4622 15374 4674 15426
rect 9886 15374 9938 15426
rect 10558 15374 10610 15426
rect 10894 15374 10946 15426
rect 11230 15374 11282 15426
rect 14254 15374 14306 15426
rect 19518 15374 19570 15426
rect 21646 15374 21698 15426
rect 26014 15374 26066 15426
rect 27694 15374 27746 15426
rect 29934 15374 29986 15426
rect 33070 15374 33122 15426
rect 33406 15374 33458 15426
rect 35870 15374 35922 15426
rect 38110 15374 38162 15426
rect 39678 15374 39730 15426
rect 5070 15262 5122 15314
rect 5518 15262 5570 15314
rect 9550 15262 9602 15314
rect 10334 15262 10386 15314
rect 11790 15262 11842 15314
rect 12574 15262 12626 15314
rect 12910 15262 12962 15314
rect 14030 15262 14082 15314
rect 17502 15262 17554 15314
rect 17726 15262 17778 15314
rect 21310 15262 21362 15314
rect 22654 15262 22706 15314
rect 23662 15262 23714 15314
rect 25230 15262 25282 15314
rect 25902 15262 25954 15314
rect 27582 15262 27634 15314
rect 30046 15262 30098 15314
rect 30494 15262 30546 15314
rect 34190 15262 34242 15314
rect 34414 15262 34466 15314
rect 35086 15262 35138 15314
rect 35534 15262 35586 15314
rect 40238 15262 40290 15314
rect 41358 15262 41410 15314
rect 42254 15262 42306 15314
rect 3502 15150 3554 15202
rect 3614 15150 3666 15202
rect 8542 15150 8594 15202
rect 13246 15150 13298 15202
rect 20750 15150 20802 15202
rect 21982 15150 22034 15202
rect 22318 15150 22370 15202
rect 24670 15150 24722 15202
rect 34862 15150 34914 15202
rect 45390 15038 45442 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 21310 14702 21362 14754
rect 33854 14702 33906 14754
rect 43038 14702 43090 14754
rect 7310 14590 7362 14642
rect 9774 14590 9826 14642
rect 11902 14590 11954 14642
rect 14702 14590 14754 14642
rect 16830 14590 16882 14642
rect 18622 14590 18674 14642
rect 23662 14590 23714 14642
rect 24110 14590 24162 14642
rect 24670 14590 24722 14642
rect 25006 14590 25058 14642
rect 25342 14590 25394 14642
rect 31726 14590 31778 14642
rect 32622 14590 32674 14642
rect 4846 14478 4898 14530
rect 7982 14478 8034 14530
rect 12574 14478 12626 14530
rect 13918 14478 13970 14530
rect 19294 14478 19346 14530
rect 19742 14478 19794 14530
rect 20526 14478 20578 14530
rect 21422 14478 21474 14530
rect 21646 14478 21698 14530
rect 25790 14478 25842 14530
rect 26126 14478 26178 14530
rect 27582 14478 27634 14530
rect 28478 14478 28530 14530
rect 29150 14478 29202 14530
rect 29374 14478 29426 14530
rect 29486 14478 29538 14530
rect 29598 14478 29650 14530
rect 29822 14478 29874 14530
rect 30158 14478 30210 14530
rect 30830 14478 30882 14530
rect 32062 14478 32114 14530
rect 33182 14478 33234 14530
rect 34190 14478 34242 14530
rect 34862 14478 34914 14530
rect 35534 14478 35586 14530
rect 38670 14478 38722 14530
rect 39006 14478 39058 14530
rect 39342 14478 39394 14530
rect 8318 14366 8370 14418
rect 26350 14366 26402 14418
rect 26798 14366 26850 14418
rect 32958 14366 33010 14418
rect 34974 14366 35026 14418
rect 36990 14366 37042 14418
rect 37774 14366 37826 14418
rect 4622 14254 4674 14306
rect 7198 14254 7250 14306
rect 18174 14254 18226 14306
rect 19966 14254 20018 14306
rect 20302 14254 20354 14306
rect 30494 14254 30546 14306
rect 31166 14254 31218 14306
rect 37326 14254 37378 14306
rect 38110 14254 38162 14306
rect 38446 14254 38498 14306
rect 42366 14254 42418 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 4510 13918 4562 13970
rect 5294 13918 5346 13970
rect 8318 13918 8370 13970
rect 18734 13918 18786 13970
rect 24110 13918 24162 13970
rect 25454 13918 25506 13970
rect 27806 13918 27858 13970
rect 29038 13918 29090 13970
rect 29598 13918 29650 13970
rect 34974 13918 35026 13970
rect 38782 13918 38834 13970
rect 40910 13918 40962 13970
rect 11118 13806 11170 13858
rect 14142 13806 14194 13858
rect 15150 13806 15202 13858
rect 15822 13806 15874 13858
rect 17950 13806 18002 13858
rect 22318 13806 22370 13858
rect 25678 13806 25730 13858
rect 26014 13806 26066 13858
rect 26350 13806 26402 13858
rect 27470 13806 27522 13858
rect 28478 13806 28530 13858
rect 32062 13806 32114 13858
rect 33966 13806 34018 13858
rect 35422 13806 35474 13858
rect 37998 13806 38050 13858
rect 39342 13806 39394 13858
rect 39902 13806 39954 13858
rect 45278 13806 45330 13858
rect 1822 13694 1874 13746
rect 2158 13694 2210 13746
rect 5630 13694 5682 13746
rect 6078 13694 6130 13746
rect 10334 13694 10386 13746
rect 14478 13694 14530 13746
rect 14814 13694 14866 13746
rect 15486 13694 15538 13746
rect 18286 13694 18338 13746
rect 19630 13694 19682 13746
rect 26686 13694 26738 13746
rect 28142 13694 28194 13746
rect 29262 13694 29314 13746
rect 30494 13694 30546 13746
rect 31614 13694 31666 13746
rect 32286 13694 32338 13746
rect 33630 13694 33682 13746
rect 34414 13694 34466 13746
rect 35310 13694 35362 13746
rect 37662 13694 37714 13746
rect 38222 13694 38274 13746
rect 41134 13694 41186 13746
rect 42702 13694 42754 13746
rect 43710 13694 43762 13746
rect 13246 13582 13298 13634
rect 17614 13582 17666 13634
rect 29934 13582 29986 13634
rect 31278 13582 31330 13634
rect 33070 13582 33122 13634
rect 36318 13582 36370 13634
rect 9102 13470 9154 13522
rect 39118 13470 39170 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 16942 13134 16994 13186
rect 30046 13134 30098 13186
rect 32286 13134 32338 13186
rect 8654 13022 8706 13074
rect 18174 13022 18226 13074
rect 37326 13022 37378 13074
rect 37998 13022 38050 13074
rect 13694 12910 13746 12962
rect 14254 12910 14306 12962
rect 14590 12910 14642 12962
rect 15262 12910 15314 12962
rect 15822 12910 15874 12962
rect 17726 12910 17778 12962
rect 19070 12910 19122 12962
rect 19854 12910 19906 12962
rect 20414 12910 20466 12962
rect 23886 12910 23938 12962
rect 24446 12910 24498 12962
rect 26462 12910 26514 12962
rect 26910 12910 26962 12962
rect 27582 12910 27634 12962
rect 29822 12910 29874 12962
rect 30270 12910 30322 12962
rect 30382 12910 30434 12962
rect 31054 12910 31106 12962
rect 31390 12910 31442 12962
rect 32510 12910 32562 12962
rect 32734 12910 32786 12962
rect 33630 12910 33682 12962
rect 33966 12910 34018 12962
rect 34862 12910 34914 12962
rect 35422 12910 35474 12962
rect 36318 12910 36370 12962
rect 37550 12910 37602 12962
rect 40238 12910 40290 12962
rect 40686 12910 40738 12962
rect 42142 12910 42194 12962
rect 43038 12910 43090 12962
rect 3614 12798 3666 12850
rect 12910 12798 12962 12850
rect 13918 12798 13970 12850
rect 14926 12798 14978 12850
rect 16718 12798 16770 12850
rect 18510 12798 18562 12850
rect 19406 12798 19458 12850
rect 23326 12798 23378 12850
rect 25566 12798 25618 12850
rect 27806 12798 27858 12850
rect 31838 12798 31890 12850
rect 32062 12798 32114 12850
rect 33182 12798 33234 12850
rect 34190 12798 34242 12850
rect 38670 12798 38722 12850
rect 39678 12798 39730 12850
rect 39902 12798 39954 12850
rect 40910 12798 40962 12850
rect 41358 12798 41410 12850
rect 3502 12686 3554 12738
rect 8542 12686 8594 12738
rect 12574 12686 12626 12738
rect 17278 12686 17330 12738
rect 24558 12686 24610 12738
rect 24782 12686 24834 12738
rect 25230 12686 25282 12738
rect 27470 12686 27522 12738
rect 32174 12686 32226 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4734 12350 4786 12402
rect 5294 12350 5346 12402
rect 11790 12350 11842 12402
rect 12014 12350 12066 12402
rect 12686 12350 12738 12402
rect 18174 12350 18226 12402
rect 20302 12350 20354 12402
rect 21534 12350 21586 12402
rect 22206 12350 22258 12402
rect 26238 12350 26290 12402
rect 30270 12350 30322 12402
rect 35758 12350 35810 12402
rect 40238 12350 40290 12402
rect 41134 12350 41186 12402
rect 41806 12350 41858 12402
rect 45838 12350 45890 12402
rect 6190 12238 6242 12290
rect 12350 12238 12402 12290
rect 13022 12238 13074 12290
rect 19294 12238 19346 12290
rect 19742 12238 19794 12290
rect 21086 12238 21138 12290
rect 22542 12238 22594 12290
rect 22878 12238 22930 12290
rect 23214 12238 23266 12290
rect 33742 12238 33794 12290
rect 35646 12238 35698 12290
rect 36542 12238 36594 12290
rect 37662 12238 37714 12290
rect 1822 12126 1874 12178
rect 2158 12126 2210 12178
rect 8430 12126 8482 12178
rect 8878 12126 8930 12178
rect 13470 12126 13522 12178
rect 16494 12126 16546 12178
rect 17838 12126 17890 12178
rect 17950 12126 18002 12178
rect 18398 12126 18450 12178
rect 20750 12126 20802 12178
rect 23438 12126 23490 12178
rect 24334 12126 24386 12178
rect 25566 12126 25618 12178
rect 26126 12126 26178 12178
rect 26798 12126 26850 12178
rect 27470 12126 27522 12178
rect 28254 12126 28306 12178
rect 29598 12126 29650 12178
rect 30046 12126 30098 12178
rect 30942 12126 30994 12178
rect 31502 12126 31554 12178
rect 32398 12126 32450 12178
rect 33070 12126 33122 12178
rect 33630 12126 33682 12178
rect 34974 12126 35026 12178
rect 35534 12126 35586 12178
rect 36654 12126 36706 12178
rect 42030 12126 42082 12178
rect 42366 12126 42418 12178
rect 42814 12126 42866 12178
rect 9662 12014 9714 12066
rect 10110 12014 10162 12066
rect 13918 12014 13970 12066
rect 15374 12014 15426 12066
rect 23886 12014 23938 12066
rect 25230 12014 25282 12066
rect 29262 12014 29314 12066
rect 34078 12014 34130 12066
rect 5406 11902 5458 11954
rect 9550 11902 9602 11954
rect 9998 11902 10050 11954
rect 18286 11902 18338 11954
rect 19966 11902 20018 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 4062 11566 4114 11618
rect 11006 11566 11058 11618
rect 42478 11566 42530 11618
rect 3726 11454 3778 11506
rect 6190 11454 6242 11506
rect 19854 11454 19906 11506
rect 26126 11454 26178 11506
rect 29598 11454 29650 11506
rect 30606 11454 30658 11506
rect 32174 11454 32226 11506
rect 33966 11454 34018 11506
rect 34638 11454 34690 11506
rect 3614 11342 3666 11394
rect 5630 11342 5682 11394
rect 7310 11342 7362 11394
rect 7982 11342 8034 11394
rect 11342 11342 11394 11394
rect 12014 11342 12066 11394
rect 12686 11342 12738 11394
rect 14702 11342 14754 11394
rect 15038 11342 15090 11394
rect 16382 11342 16434 11394
rect 16830 11342 16882 11394
rect 18062 11342 18114 11394
rect 19182 11342 19234 11394
rect 19630 11342 19682 11394
rect 20078 11342 20130 11394
rect 21310 11342 21362 11394
rect 22654 11342 22706 11394
rect 23102 11342 23154 11394
rect 23886 11342 23938 11394
rect 24222 11342 24274 11394
rect 26014 11342 26066 11394
rect 26350 11342 26402 11394
rect 27806 11342 27858 11394
rect 30158 11342 30210 11394
rect 31726 11342 31778 11394
rect 33518 11342 33570 11394
rect 34526 11342 34578 11394
rect 37214 11342 37266 11394
rect 37774 11342 37826 11394
rect 37998 11342 38050 11394
rect 38334 11342 38386 11394
rect 38670 11342 38722 11394
rect 4174 11230 4226 11282
rect 11566 11230 11618 11282
rect 12910 11230 12962 11282
rect 15710 11230 15762 11282
rect 16046 11230 16098 11282
rect 17054 11230 17106 11282
rect 17502 11230 17554 11282
rect 27358 11230 27410 11282
rect 36990 11230 37042 11282
rect 41582 11230 41634 11282
rect 10334 11118 10386 11170
rect 12238 11118 12290 11170
rect 21422 11118 21474 11170
rect 29150 11118 29202 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4734 10782 4786 10834
rect 5294 10782 5346 10834
rect 6078 10782 6130 10834
rect 12462 10782 12514 10834
rect 19518 10782 19570 10834
rect 23662 10782 23714 10834
rect 24446 10782 24498 10834
rect 24558 10782 24610 10834
rect 24670 10782 24722 10834
rect 33182 10782 33234 10834
rect 33294 10782 33346 10834
rect 33406 10782 33458 10834
rect 14814 10670 14866 10722
rect 22542 10670 22594 10722
rect 23102 10670 23154 10722
rect 26238 10670 26290 10722
rect 28254 10670 28306 10722
rect 1822 10558 1874 10610
rect 2158 10558 2210 10610
rect 8430 10558 8482 10610
rect 9102 10558 9154 10610
rect 9662 10558 9714 10610
rect 9998 10558 10050 10610
rect 13470 10558 13522 10610
rect 13918 10558 13970 10610
rect 14366 10558 14418 10610
rect 16046 10558 16098 10610
rect 17390 10558 17442 10610
rect 17614 10558 17666 10610
rect 17726 10558 17778 10610
rect 18958 10558 19010 10610
rect 19294 10558 19346 10610
rect 19966 10558 20018 10610
rect 20750 10558 20802 10610
rect 21646 10558 21698 10610
rect 23998 10558 24050 10610
rect 27022 10558 27074 10610
rect 29934 10558 29986 10610
rect 30382 10558 30434 10610
rect 31502 10558 31554 10610
rect 16606 10446 16658 10498
rect 18174 10446 18226 10498
rect 18510 10446 18562 10498
rect 25678 10446 25730 10498
rect 29598 10446 29650 10498
rect 33630 10446 33682 10498
rect 33854 10446 33906 10498
rect 5406 10334 5458 10386
rect 13134 10334 13186 10386
rect 23326 10334 23378 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 6078 9998 6130 10050
rect 11454 9998 11506 10050
rect 13918 9998 13970 10050
rect 14030 9998 14082 10050
rect 14254 9998 14306 10050
rect 21870 9998 21922 10050
rect 23214 9998 23266 10050
rect 5966 9886 6018 9938
rect 19294 9886 19346 9938
rect 30270 9886 30322 9938
rect 32622 9886 32674 9938
rect 7982 9774 8034 9826
rect 8430 9774 8482 9826
rect 12910 9774 12962 9826
rect 15486 9774 15538 9826
rect 15934 9774 15986 9826
rect 16830 9774 16882 9826
rect 17278 9774 17330 9826
rect 18286 9774 18338 9826
rect 20190 9774 20242 9826
rect 21310 9774 21362 9826
rect 22990 9774 23042 9826
rect 24446 9774 24498 9826
rect 24782 9774 24834 9826
rect 26126 9774 26178 9826
rect 27134 9774 27186 9826
rect 29598 9774 29650 9826
rect 31166 9774 31218 9826
rect 32062 9774 32114 9826
rect 33294 9774 33346 9826
rect 33742 9774 33794 9826
rect 34638 9774 34690 9826
rect 35086 9774 35138 9826
rect 35982 9774 36034 9826
rect 38782 9774 38834 9826
rect 39342 9774 39394 9826
rect 39902 9774 39954 9826
rect 40686 9774 40738 9826
rect 41582 9774 41634 9826
rect 4286 9662 4338 9714
rect 4958 9662 5010 9714
rect 10670 9662 10722 9714
rect 12574 9662 12626 9714
rect 14814 9662 14866 9714
rect 15150 9662 15202 9714
rect 19966 9662 20018 9714
rect 23550 9662 23602 9714
rect 23998 9662 24050 9714
rect 25006 9662 25058 9714
rect 25454 9662 25506 9714
rect 29822 9662 29874 9714
rect 31390 9662 31442 9714
rect 31726 9662 31778 9714
rect 32958 9662 33010 9714
rect 33966 9662 34018 9714
rect 38446 9662 38498 9714
rect 39454 9662 39506 9714
rect 4174 9550 4226 9602
rect 4846 9550 4898 9602
rect 16158 9550 16210 9602
rect 20638 9550 20690 9602
rect 30718 9550 30770 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 2942 9214 2994 9266
rect 3726 9214 3778 9266
rect 9886 9214 9938 9266
rect 18174 9214 18226 9266
rect 30942 9214 30994 9266
rect 31726 9214 31778 9266
rect 32062 9214 32114 9266
rect 32398 9214 32450 9266
rect 33406 9214 33458 9266
rect 38558 9214 38610 9266
rect 43374 9214 43426 9266
rect 13582 9102 13634 9154
rect 15598 9102 15650 9154
rect 18622 9102 18674 9154
rect 19070 9102 19122 9154
rect 23326 9102 23378 9154
rect 26126 9102 26178 9154
rect 29598 9102 29650 9154
rect 37550 9102 37602 9154
rect 41246 9102 41298 9154
rect 41806 9102 41858 9154
rect 5966 8990 6018 9042
rect 6638 8990 6690 9042
rect 9998 8990 10050 9042
rect 13470 8990 13522 9042
rect 14366 8990 14418 9042
rect 20638 8990 20690 9042
rect 22990 8990 23042 9042
rect 23662 8990 23714 9042
rect 24110 8990 24162 9042
rect 25230 8990 25282 9042
rect 26238 8990 26290 9042
rect 29822 8990 29874 9042
rect 33182 8990 33234 9042
rect 34862 8990 34914 9042
rect 35422 8990 35474 9042
rect 14478 8878 14530 8930
rect 20190 8878 20242 8930
rect 25678 8878 25730 8930
rect 31278 8878 31330 8930
rect 41582 8878 41634 8930
rect 19294 8766 19346 8818
rect 19630 8766 19682 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 13582 8318 13634 8370
rect 15822 8318 15874 8370
rect 23326 8318 23378 8370
rect 35086 8318 35138 8370
rect 13694 8206 13746 8258
rect 15038 8206 15090 8258
rect 18734 8206 18786 8258
rect 19182 8206 19234 8258
rect 19742 8206 19794 8258
rect 20302 8206 20354 8258
rect 21646 8206 21698 8258
rect 22990 8206 23042 8258
rect 24894 8206 24946 8258
rect 26910 8206 26962 8258
rect 30830 8206 30882 8258
rect 31278 8206 31330 8258
rect 31838 8206 31890 8258
rect 35758 8206 35810 8258
rect 37886 8206 37938 8258
rect 38446 8206 38498 8258
rect 40910 8206 40962 8258
rect 19966 8094 20018 8146
rect 22318 8094 22370 8146
rect 22766 8094 22818 8146
rect 24670 8094 24722 8146
rect 25118 8094 25170 8146
rect 26686 8094 26738 8146
rect 27022 8094 27074 8146
rect 27582 8094 27634 8146
rect 30606 8094 30658 8146
rect 34078 8094 34130 8146
rect 18958 7982 19010 8034
rect 20638 7982 20690 8034
rect 21310 7982 21362 8034
rect 23886 7982 23938 8034
rect 24222 7982 24274 8034
rect 25902 7982 25954 8034
rect 36094 7982 36146 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4958 7646 5010 7698
rect 5518 7646 5570 7698
rect 21982 7646 22034 7698
rect 26798 7646 26850 7698
rect 32398 7646 32450 7698
rect 35534 7646 35586 7698
rect 38558 7646 38610 7698
rect 19070 7534 19122 7586
rect 19854 7534 19906 7586
rect 21310 7534 21362 7586
rect 25790 7534 25842 7586
rect 27246 7534 27298 7586
rect 30158 7534 30210 7586
rect 2046 7422 2098 7474
rect 2494 7422 2546 7474
rect 18846 7422 18898 7474
rect 22878 7422 22930 7474
rect 24110 7422 24162 7474
rect 24670 7422 24722 7474
rect 26126 7422 26178 7474
rect 26686 7422 26738 7474
rect 28030 7422 28082 7474
rect 28814 7422 28866 7474
rect 29486 7422 29538 7474
rect 33630 7422 33682 7474
rect 33966 7422 34018 7474
rect 34302 7422 34354 7474
rect 35646 7422 35698 7474
rect 36206 7422 36258 7474
rect 19518 7310 19570 7362
rect 21646 7310 21698 7362
rect 22430 7310 22482 7362
rect 23438 7310 23490 7362
rect 39342 7198 39394 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 28030 6862 28082 6914
rect 33742 6862 33794 6914
rect 19294 6750 19346 6802
rect 15486 6638 15538 6690
rect 21646 6638 21698 6690
rect 22094 6638 22146 6690
rect 22878 6638 22930 6690
rect 23326 6638 23378 6690
rect 24446 6638 24498 6690
rect 24894 6638 24946 6690
rect 25454 6638 25506 6690
rect 28366 6638 28418 6690
rect 29486 6638 29538 6690
rect 30158 6638 30210 6690
rect 30606 6638 30658 6690
rect 32846 6638 32898 6690
rect 19854 6526 19906 6578
rect 20638 6526 20690 6578
rect 21310 6526 21362 6578
rect 22318 6526 22370 6578
rect 29150 6526 29202 6578
rect 18286 6414 18338 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 5070 6078 5122 6130
rect 5854 6078 5906 6130
rect 22430 6078 22482 6130
rect 25342 6078 25394 6130
rect 15934 5966 15986 6018
rect 16158 5966 16210 6018
rect 17502 5966 17554 6018
rect 18510 5966 18562 6018
rect 19854 5966 19906 6018
rect 2158 5854 2210 5906
rect 2718 5854 2770 5906
rect 15598 5854 15650 5906
rect 16382 5854 16434 5906
rect 18622 5854 18674 5906
rect 21198 5854 21250 5906
rect 21758 5854 21810 5906
rect 22206 5854 22258 5906
rect 22878 5854 22930 5906
rect 23662 5854 23714 5906
rect 24558 5854 24610 5906
rect 25230 5854 25282 5906
rect 25678 5854 25730 5906
rect 27582 5854 27634 5906
rect 21422 5742 21474 5794
rect 28814 5742 28866 5794
rect 16718 5630 16770 5682
rect 25454 5630 25506 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 27582 5294 27634 5346
rect 21422 5182 21474 5234
rect 22990 5182 23042 5234
rect 24558 5182 24610 5234
rect 15262 5070 15314 5122
rect 20414 5070 20466 5122
rect 21534 5070 21586 5122
rect 23550 5070 23602 5122
rect 25006 5070 25058 5122
rect 28590 5070 28642 5122
rect 20750 4958 20802 5010
rect 23886 4958 23938 5010
rect 24894 4958 24946 5010
rect 1710 4846 1762 4898
rect 18510 4846 18562 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 19630 4510 19682 4562
rect 22094 4510 22146 4562
rect 23662 4510 23714 4562
rect 19182 4398 19234 4450
rect 20638 4398 20690 4450
rect 20974 4398 21026 4450
rect 23102 4398 23154 4450
rect 24670 4398 24722 4450
rect 17502 4286 17554 4338
rect 18510 4286 18562 4338
rect 19742 4286 19794 4338
rect 20302 4286 20354 4338
rect 21422 4286 21474 4338
rect 21646 4286 21698 4338
rect 23550 4286 23602 4338
rect 24110 4286 24162 4338
rect 21198 4062 21250 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 19854 3502 19906 3554
rect 19518 3390 19570 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 1708 43764 1764 43802
rect 1708 43698 1764 43708
rect 28364 43762 28420 43774
rect 28364 43710 28366 43762
rect 28418 43710 28420 43762
rect 13244 43650 13300 43662
rect 13244 43598 13246 43650
rect 13298 43598 13300 43650
rect 13020 43538 13076 43550
rect 13020 43486 13022 43538
rect 13074 43486 13076 43538
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 1708 42532 1764 42542
rect 1708 42438 1764 42476
rect 12796 41970 12852 41982
rect 12796 41918 12798 41970
rect 12850 41918 12852 41970
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 12572 40962 12628 40974
rect 12572 40910 12574 40962
rect 12626 40910 12628 40962
rect 11900 40628 11956 40638
rect 11452 40514 11508 40526
rect 11452 40462 11454 40514
rect 11506 40462 11508 40514
rect 11228 40402 11284 40414
rect 11228 40350 11230 40402
rect 11282 40350 11284 40402
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 9212 39506 9268 39518
rect 9212 39454 9214 39506
rect 9266 39454 9268 39506
rect 7644 39396 7700 39406
rect 4844 39060 4900 39070
rect 4844 39058 5012 39060
rect 4844 39006 4846 39058
rect 4898 39006 5012 39058
rect 4844 39004 5012 39006
rect 4844 38994 4900 39004
rect 1932 38836 1988 38846
rect 1932 38834 2212 38836
rect 1932 38782 1934 38834
rect 1986 38782 2212 38834
rect 1932 38780 2212 38782
rect 1932 38770 1988 38780
rect 2044 36372 2100 36382
rect 1708 34802 1764 34814
rect 1708 34750 1710 34802
rect 1762 34750 1764 34802
rect 1708 34356 1764 34750
rect 2044 34802 2100 36316
rect 2044 34750 2046 34802
rect 2098 34750 2100 34802
rect 2044 34738 2100 34750
rect 1708 34290 1764 34300
rect 1820 34132 1876 34142
rect 1820 34130 2100 34132
rect 1820 34078 1822 34130
rect 1874 34078 2100 34130
rect 1820 34076 2100 34078
rect 1820 34066 1876 34076
rect 2044 33236 2100 34076
rect 2156 34130 2212 38780
rect 2380 38834 2436 38846
rect 2380 38782 2382 38834
rect 2434 38782 2436 38834
rect 2380 37268 2436 38782
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4956 37604 5012 39004
rect 5404 38612 5460 38622
rect 5404 38610 5572 38612
rect 5404 38558 5406 38610
rect 5458 38558 5572 38610
rect 5404 38556 5572 38558
rect 5404 38546 5460 38556
rect 4844 37548 5460 37604
rect 2716 37268 2772 37278
rect 2380 37266 2772 37268
rect 2380 37214 2718 37266
rect 2770 37214 2772 37266
rect 2380 37212 2772 37214
rect 2716 35140 2772 37212
rect 3164 37266 3220 37278
rect 3164 37214 3166 37266
rect 3218 37214 3220 37266
rect 3164 35700 3220 37214
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4844 35924 4900 37548
rect 5404 37490 5460 37548
rect 5404 37438 5406 37490
rect 5458 37438 5460 37490
rect 5404 37426 5460 37438
rect 5516 36484 5572 38556
rect 6188 37044 6244 37054
rect 5404 36428 5572 36484
rect 6076 37042 6244 37044
rect 6076 36990 6190 37042
rect 6242 36990 6244 37042
rect 6076 36988 6244 36990
rect 5180 36258 5236 36270
rect 5180 36206 5182 36258
rect 5234 36206 5236 36258
rect 5180 36148 5236 36206
rect 5180 36082 5236 36092
rect 3164 35634 3220 35644
rect 3836 35700 3892 35710
rect 3612 35586 3668 35598
rect 3612 35534 3614 35586
rect 3666 35534 3668 35586
rect 3500 35476 3556 35486
rect 3612 35476 3668 35534
rect 3556 35420 3668 35476
rect 2940 35140 2996 35150
rect 2716 35138 2996 35140
rect 2716 35086 2942 35138
rect 2994 35086 2996 35138
rect 2716 35084 2996 35086
rect 2940 35074 2996 35084
rect 3052 35028 3108 35038
rect 3052 34934 3108 34972
rect 3500 34914 3556 35420
rect 3836 35364 3892 35644
rect 4508 35700 4564 35710
rect 4508 35606 4564 35644
rect 3500 34862 3502 34914
rect 3554 34862 3556 34914
rect 3500 34850 3556 34862
rect 3612 35308 3892 35364
rect 4476 35308 4740 35318
rect 2492 34690 2548 34702
rect 2492 34638 2494 34690
rect 2546 34638 2548 34690
rect 2492 34356 2548 34638
rect 2492 34290 2548 34300
rect 2156 34078 2158 34130
rect 2210 34078 2212 34130
rect 2156 33572 2212 34078
rect 2156 33506 2212 33516
rect 1932 32562 1988 32574
rect 1932 32510 1934 32562
rect 1986 32510 1988 32562
rect 1932 31948 1988 32510
rect 2044 32564 2100 33180
rect 3612 33012 3668 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4732 34804 4788 34814
rect 4844 34804 4900 35868
rect 4732 34802 4900 34804
rect 4732 34750 4734 34802
rect 4786 34750 4900 34802
rect 4732 34748 4900 34750
rect 4956 35140 5012 35150
rect 4732 34738 4788 34748
rect 3724 34692 3780 34702
rect 4060 34692 4116 34702
rect 3724 34690 4116 34692
rect 3724 34638 3726 34690
rect 3778 34638 4062 34690
rect 4114 34638 4116 34690
rect 3724 34636 4116 34638
rect 3724 34626 3780 34636
rect 4060 33460 4116 34636
rect 4396 34692 4452 34702
rect 4396 34598 4452 34636
rect 4732 34356 4788 34366
rect 4732 34354 4900 34356
rect 4732 34302 4734 34354
rect 4786 34302 4900 34354
rect 4732 34300 4900 34302
rect 4732 34290 4788 34300
rect 4284 33908 4340 33918
rect 4172 33572 4228 33582
rect 4172 33478 4228 33516
rect 4060 33394 4116 33404
rect 4284 33458 4340 33852
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4284 33406 4286 33458
rect 4338 33406 4340 33458
rect 4284 33394 4340 33406
rect 4844 33348 4900 34300
rect 4956 33458 5012 35084
rect 5404 35028 5460 36428
rect 5404 34962 5460 34972
rect 5516 36260 5572 36270
rect 5516 35700 5572 36204
rect 5516 34914 5572 35644
rect 5628 36258 5684 36270
rect 5628 36206 5630 36258
rect 5682 36206 5684 36258
rect 5628 35588 5684 36206
rect 5964 36258 6020 36270
rect 5964 36206 5966 36258
rect 6018 36206 6020 36258
rect 5964 36148 6020 36206
rect 5964 36082 6020 36092
rect 5628 35522 5684 35532
rect 6076 35140 6132 36988
rect 6188 36978 6244 36988
rect 6300 36372 6356 36382
rect 6300 36278 6356 36316
rect 6636 36372 6692 36382
rect 7084 36372 7140 36382
rect 6636 36370 6804 36372
rect 6636 36318 6638 36370
rect 6690 36318 6804 36370
rect 6636 36316 6804 36318
rect 6636 36306 6692 36316
rect 6748 36148 6804 36316
rect 7084 36370 7588 36372
rect 7084 36318 7086 36370
rect 7138 36318 7588 36370
rect 7084 36316 7588 36318
rect 7084 36306 7140 36316
rect 6972 36260 7028 36270
rect 6972 36166 7028 36204
rect 6748 36082 6804 36092
rect 6748 35924 6804 35934
rect 6748 35830 6804 35868
rect 7532 35922 7588 36316
rect 7532 35870 7534 35922
rect 7586 35870 7588 35922
rect 7532 35858 7588 35870
rect 7644 35700 7700 39340
rect 9212 38948 9268 39454
rect 11228 39060 11284 40350
rect 11452 40292 11508 40462
rect 11900 40402 11956 40572
rect 11900 40350 11902 40402
rect 11954 40350 11956 40402
rect 11900 40338 11956 40350
rect 12124 40514 12180 40526
rect 12124 40462 12126 40514
rect 12178 40462 12180 40514
rect 11452 40226 11508 40236
rect 12124 40180 12180 40462
rect 12124 40114 12180 40124
rect 12572 40514 12628 40910
rect 12572 40462 12574 40514
rect 12626 40462 12628 40514
rect 9212 38882 9268 38892
rect 11116 39004 11228 39060
rect 10780 37268 10836 37278
rect 10780 37266 10948 37268
rect 10780 37214 10782 37266
rect 10834 37214 10948 37266
rect 10780 37212 10948 37214
rect 10780 37202 10836 37212
rect 9436 36484 9492 36494
rect 9436 36390 9492 36428
rect 10108 36482 10164 36494
rect 10108 36430 10110 36482
rect 10162 36430 10164 36482
rect 9660 36372 9716 36382
rect 9660 36278 9716 36316
rect 10108 36372 10164 36430
rect 7308 35644 7700 35700
rect 7980 36148 8036 36158
rect 6076 35074 6132 35084
rect 6188 35476 6244 35486
rect 6188 34916 6244 35420
rect 5516 34862 5518 34914
rect 5570 34862 5572 34914
rect 5516 34850 5572 34862
rect 5628 34914 6244 34916
rect 5628 34862 6190 34914
rect 6242 34862 6244 34914
rect 5628 34860 6244 34862
rect 5068 34692 5124 34702
rect 5068 34598 5124 34636
rect 5628 34130 5684 34860
rect 6188 34850 6244 34860
rect 5628 34078 5630 34130
rect 5682 34078 5684 34130
rect 5628 34066 5684 34078
rect 5964 34692 6020 34702
rect 5292 33908 5348 33918
rect 5292 33814 5348 33852
rect 4956 33406 4958 33458
rect 5010 33406 5012 33458
rect 4956 33394 5012 33406
rect 4732 33292 4844 33348
rect 3724 33236 3780 33246
rect 3724 33142 3780 33180
rect 3836 33234 3892 33246
rect 3836 33182 3838 33234
rect 3890 33182 3892 33234
rect 3724 33012 3780 33022
rect 3612 32956 3724 33012
rect 3724 32946 3780 32956
rect 3836 32788 3892 33182
rect 3836 32722 3892 32732
rect 4732 32788 4788 33292
rect 4844 33282 4900 33292
rect 5628 33348 5684 33358
rect 5964 33348 6020 34636
rect 6076 34130 6132 34142
rect 6076 34078 6078 34130
rect 6130 34078 6132 34130
rect 6076 33908 6132 34078
rect 6076 33842 6132 33852
rect 6636 33908 6692 33918
rect 6188 33460 6244 33470
rect 6076 33348 6132 33358
rect 5964 33346 6132 33348
rect 5964 33294 6078 33346
rect 6130 33294 6132 33346
rect 5964 33292 6132 33294
rect 5628 33254 5684 33292
rect 6076 33282 6132 33292
rect 4844 33122 4900 33134
rect 4844 33070 4846 33122
rect 4898 33070 4900 33122
rect 4844 33012 4900 33070
rect 4844 32946 4900 32956
rect 5404 32788 5460 32798
rect 4732 32786 4900 32788
rect 4732 32734 4734 32786
rect 4786 32734 4900 32786
rect 4732 32732 4900 32734
rect 4732 32722 4788 32732
rect 2268 32564 2324 32574
rect 2044 32562 2324 32564
rect 2044 32510 2270 32562
rect 2322 32510 2324 32562
rect 2044 32508 2324 32510
rect 2268 32498 2324 32508
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 1932 31892 2548 31948
rect 2492 31556 2548 31892
rect 3948 31668 4004 31678
rect 3948 31574 4004 31612
rect 2044 30996 2100 31006
rect 2044 30994 2324 30996
rect 2044 30942 2046 30994
rect 2098 30942 2324 30994
rect 2044 30940 2324 30942
rect 2044 30930 2100 30940
rect 2268 30212 2324 30940
rect 2492 30994 2548 31500
rect 3836 31556 3892 31566
rect 3836 31462 3892 31500
rect 2492 30942 2494 30994
rect 2546 30942 2548 30994
rect 2492 30930 2548 30942
rect 4844 31218 4900 32732
rect 5404 32694 5460 32732
rect 6188 31948 6244 33404
rect 6636 33346 6692 33852
rect 6636 33294 6638 33346
rect 6690 33294 6692 33346
rect 6636 33282 6692 33294
rect 6972 33346 7028 33358
rect 6972 33294 6974 33346
rect 7026 33294 7028 33346
rect 5964 31892 6244 31948
rect 6972 32788 7028 33294
rect 4844 31166 4846 31218
rect 4898 31166 4900 31218
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 1820 29426 1876 29438
rect 1820 29374 1822 29426
rect 1874 29374 1876 29426
rect 1820 28644 1876 29374
rect 2268 29426 2324 30156
rect 3724 30212 3780 30222
rect 3724 30118 3780 30156
rect 3836 30100 3892 30110
rect 3836 30006 3892 30044
rect 4844 29650 4900 31166
rect 5516 31668 5572 31678
rect 5516 31218 5572 31612
rect 5516 31166 5518 31218
rect 5570 31166 5572 31218
rect 5516 31154 5572 31166
rect 5404 30100 5460 30110
rect 4844 29598 4846 29650
rect 4898 29598 4900 29650
rect 4844 29586 4900 29598
rect 5068 29652 5124 29662
rect 2268 29374 2270 29426
rect 2322 29374 2324 29426
rect 2268 29362 2324 29374
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 1820 28578 1876 28588
rect 1932 28754 1988 28766
rect 1932 28702 1934 28754
rect 1986 28702 1988 28754
rect 1708 27858 1764 27870
rect 1708 27806 1710 27858
rect 1762 27806 1764 27858
rect 1708 21812 1764 27806
rect 1932 27636 1988 28702
rect 2268 28644 2324 28654
rect 2268 27858 2324 28588
rect 4284 28642 4340 28654
rect 4284 28590 4286 28642
rect 4338 28590 4340 28642
rect 4284 28084 4340 28590
rect 4956 28644 5012 28654
rect 5068 28644 5124 29596
rect 5404 29650 5460 30044
rect 5404 29598 5406 29650
rect 5458 29598 5460 29650
rect 5404 29586 5460 29598
rect 5628 29652 5684 29662
rect 5628 29558 5684 29596
rect 5964 29538 6020 31892
rect 6972 31778 7028 32732
rect 6972 31726 6974 31778
rect 7026 31726 7028 31778
rect 6972 31714 7028 31726
rect 5964 29486 5966 29538
rect 6018 29486 6020 29538
rect 5964 29474 6020 29486
rect 4956 28642 5124 28644
rect 4956 28590 4958 28642
rect 5010 28590 5124 28642
rect 4956 28588 5124 28590
rect 4956 28578 5012 28588
rect 4620 28420 4676 28430
rect 4620 28418 4788 28420
rect 4620 28366 4622 28418
rect 4674 28366 4788 28418
rect 4620 28364 4788 28366
rect 4620 28354 4676 28364
rect 4284 28018 4340 28028
rect 4732 28082 4788 28364
rect 4732 28030 4734 28082
rect 4786 28030 4788 28082
rect 4732 27972 4788 28030
rect 4732 27906 4788 27916
rect 2268 27806 2270 27858
rect 2322 27806 2324 27858
rect 2268 27794 2324 27806
rect 1932 27570 1988 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 1932 27188 1988 27198
rect 1932 27094 1988 27132
rect 4284 27076 4340 27086
rect 4284 26982 4340 27020
rect 2380 26964 2436 26974
rect 2268 26852 2436 26908
rect 3164 26964 3220 26974
rect 1932 26292 1988 26302
rect 1932 25730 1988 26236
rect 1932 25678 1934 25730
rect 1986 25678 1988 25730
rect 1932 25666 1988 25678
rect 2268 24722 2324 26852
rect 2716 26290 2772 26302
rect 2716 26238 2718 26290
rect 2770 26238 2772 26290
rect 2716 25732 2772 26238
rect 3164 26290 3220 26908
rect 4620 26964 4676 26974
rect 4620 26870 4676 26908
rect 4732 26964 4788 26974
rect 4732 26962 4900 26964
rect 4732 26910 4734 26962
rect 4786 26910 4900 26962
rect 4732 26908 4900 26910
rect 4732 26898 4788 26908
rect 3164 26238 3166 26290
rect 3218 26238 3220 26290
rect 3164 26226 3220 26238
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4844 25844 4900 26908
rect 5068 26068 5124 28588
rect 5628 28644 5684 28654
rect 5628 28550 5684 28588
rect 5740 28530 5796 28542
rect 5740 28478 5742 28530
rect 5794 28478 5796 28530
rect 5740 28196 5796 28478
rect 5292 28140 5796 28196
rect 5292 28082 5348 28140
rect 5292 28030 5294 28082
rect 5346 28030 5348 28082
rect 5292 28018 5348 28030
rect 6636 27972 6692 27982
rect 6636 27878 6692 27916
rect 6748 27860 6804 27870
rect 7196 27860 7252 27870
rect 6748 27858 7252 27860
rect 6748 27806 6750 27858
rect 6802 27806 7198 27858
rect 7250 27806 7252 27858
rect 6748 27804 7252 27806
rect 6748 27794 6804 27804
rect 7196 27794 7252 27804
rect 5068 26002 5124 26012
rect 5404 26402 5460 26414
rect 5404 26350 5406 26402
rect 5458 26350 5460 26402
rect 5404 26292 5460 26350
rect 6412 26292 6468 26302
rect 5404 26290 6468 26292
rect 5404 26238 6414 26290
rect 6466 26238 6468 26290
rect 5404 26236 6468 26238
rect 4844 25778 4900 25788
rect 2716 25666 2772 25676
rect 4620 25732 4676 25742
rect 4620 25638 4676 25676
rect 2828 25620 2884 25630
rect 2268 24670 2270 24722
rect 2322 24670 2324 24722
rect 2268 24658 2324 24670
rect 2716 24722 2772 24734
rect 2716 24670 2718 24722
rect 2770 24670 2772 24722
rect 1820 24612 1876 24622
rect 1820 24518 1876 24556
rect 1932 24500 1988 24510
rect 2716 24500 2772 24670
rect 1932 24498 2772 24500
rect 1932 24446 1934 24498
rect 1986 24446 2772 24498
rect 1932 24444 2772 24446
rect 1932 23154 1988 24444
rect 1932 23102 1934 23154
rect 1986 23102 1988 23154
rect 1932 23090 1988 23102
rect 2044 24276 2100 24286
rect 2044 22482 2100 24220
rect 2828 24162 2884 25564
rect 4284 25620 4340 25630
rect 4284 25506 4340 25564
rect 4284 25454 4286 25506
rect 4338 25454 4340 25506
rect 4284 25442 4340 25454
rect 4732 25396 4788 25406
rect 4732 25302 4788 25340
rect 2828 24110 2830 24162
rect 2882 24110 2884 24162
rect 2828 24098 2884 24110
rect 4284 24836 4340 24846
rect 5068 24836 5124 24846
rect 5404 24836 5460 26236
rect 6412 26226 6468 26236
rect 6972 26290 7028 26302
rect 6972 26238 6974 26290
rect 7026 26238 7028 26290
rect 6188 26066 6244 26078
rect 6188 26014 6190 26066
rect 6242 26014 6244 26066
rect 6188 25844 6244 26014
rect 6972 26068 7028 26238
rect 6972 26002 7028 26012
rect 6188 25778 6244 25788
rect 5852 25618 5908 25630
rect 5852 25566 5854 25618
rect 5906 25566 5908 25618
rect 5852 25284 5908 25566
rect 5852 25218 5908 25228
rect 6636 25508 6692 25518
rect 6636 24946 6692 25452
rect 7308 24948 7364 35644
rect 7868 35586 7924 35598
rect 7868 35534 7870 35586
rect 7922 35534 7924 35586
rect 7756 35476 7812 35486
rect 7756 35382 7812 35420
rect 7868 35140 7924 35534
rect 7868 35074 7924 35084
rect 7980 31948 8036 36092
rect 10108 35922 10164 36316
rect 10780 36370 10836 36382
rect 10780 36318 10782 36370
rect 10834 36318 10836 36370
rect 10780 36260 10836 36318
rect 10892 36372 10948 37212
rect 10892 36306 10948 36316
rect 11116 36484 11172 39004
rect 11228 38994 11284 39004
rect 11676 38948 11732 38958
rect 11676 38854 11732 38892
rect 12572 38948 12628 40462
rect 12796 40292 12852 41918
rect 12908 40962 12964 40974
rect 12908 40910 12910 40962
rect 12962 40910 12964 40962
rect 12908 40404 12964 40910
rect 12908 40338 12964 40348
rect 12796 40180 12852 40236
rect 12796 40124 12964 40180
rect 12572 38882 12628 38892
rect 12796 39394 12852 39406
rect 12796 39342 12798 39394
rect 12850 39342 12852 39394
rect 12796 38052 12852 39342
rect 12908 39284 12964 40124
rect 12908 39218 12964 39228
rect 12796 37986 12852 37996
rect 13020 37492 13076 43486
rect 13244 42756 13300 43598
rect 28252 43650 28308 43662
rect 28252 43598 28254 43650
rect 28306 43598 28308 43650
rect 19180 43540 19236 43550
rect 22876 43540 22932 43550
rect 19180 43538 19572 43540
rect 19180 43486 19182 43538
rect 19234 43486 19572 43538
rect 19180 43484 19572 43486
rect 19180 43474 19236 43484
rect 13580 42756 13636 42766
rect 13244 42754 13636 42756
rect 13244 42702 13582 42754
rect 13634 42702 13636 42754
rect 13244 42700 13636 42702
rect 13580 42084 13636 42700
rect 14924 42756 14980 42766
rect 14924 42754 15092 42756
rect 14924 42702 14926 42754
rect 14978 42702 15092 42754
rect 14924 42700 15092 42702
rect 14924 42690 14980 42700
rect 13580 42018 13636 42028
rect 14140 41970 14196 41982
rect 14140 41918 14142 41970
rect 14194 41918 14196 41970
rect 13692 41188 13748 41198
rect 13692 41094 13748 41132
rect 14140 41188 14196 41918
rect 14140 41186 14420 41188
rect 14140 41134 14142 41186
rect 14194 41134 14420 41186
rect 14140 41132 14420 41134
rect 14140 41122 14196 41132
rect 13468 40962 13524 40974
rect 13468 40910 13470 40962
rect 13522 40910 13524 40962
rect 13468 40292 13524 40910
rect 13804 40460 14308 40516
rect 13468 40226 13524 40236
rect 13692 40404 13748 40414
rect 13692 39730 13748 40348
rect 13692 39678 13694 39730
rect 13746 39678 13748 39730
rect 13692 39666 13748 39678
rect 13804 39508 13860 40460
rect 14252 40402 14308 40460
rect 14252 40350 14254 40402
rect 14306 40350 14308 40402
rect 14252 40338 14308 40350
rect 13916 40292 13972 40302
rect 13916 40290 14196 40292
rect 13916 40238 13918 40290
rect 13970 40238 14196 40290
rect 13916 40236 14196 40238
rect 13916 40226 13972 40236
rect 13580 39452 13860 39508
rect 13468 38948 13524 38958
rect 13468 37938 13524 38892
rect 13468 37886 13470 37938
rect 13522 37886 13524 37938
rect 13468 37874 13524 37886
rect 13020 37426 13076 37436
rect 13468 37492 13524 37502
rect 13580 37492 13636 39452
rect 13692 39284 13748 39294
rect 13692 38050 13748 39228
rect 14140 39172 14196 40236
rect 14364 40180 14420 41132
rect 14588 41186 14644 41198
rect 14588 41134 14590 41186
rect 14642 41134 14644 41186
rect 14588 40404 14644 41134
rect 15036 40516 15092 42700
rect 17948 42642 18004 42654
rect 17948 42590 17950 42642
rect 18002 42590 18004 42642
rect 17388 42084 17444 42094
rect 16044 41860 16100 41870
rect 16044 41766 16100 41804
rect 17388 40964 17444 42028
rect 17948 41860 18004 42590
rect 19516 42196 19572 43484
rect 19852 43426 19908 43438
rect 19852 43374 19854 43426
rect 19906 43374 19908 43426
rect 19740 42644 19796 42654
rect 19852 42644 19908 43374
rect 22316 43426 22372 43438
rect 22316 43374 22318 43426
rect 22370 43374 22372 43426
rect 20076 42756 20132 42766
rect 21980 42756 22036 42766
rect 20076 42754 20356 42756
rect 20076 42702 20078 42754
rect 20130 42702 20356 42754
rect 20076 42700 20356 42702
rect 20076 42690 20132 42700
rect 19740 42642 19852 42644
rect 19740 42590 19742 42642
rect 19794 42590 19852 42642
rect 19740 42588 19852 42590
rect 19740 42578 19796 42588
rect 19852 42550 19908 42588
rect 20188 42532 20244 42542
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19516 41970 19572 42140
rect 19516 41918 19518 41970
rect 19570 41918 19572 41970
rect 17388 40962 17556 40964
rect 17388 40910 17390 40962
rect 17442 40910 17556 40962
rect 17388 40908 17556 40910
rect 17388 40898 17444 40908
rect 16044 40628 16100 40638
rect 15148 40516 15204 40526
rect 15036 40460 15148 40516
rect 14588 40338 14644 40348
rect 15148 40402 15204 40460
rect 15148 40350 15150 40402
rect 15202 40350 15204 40402
rect 15148 40338 15204 40350
rect 15932 40514 15988 40526
rect 15932 40462 15934 40514
rect 15986 40462 15988 40514
rect 14364 39620 14420 40124
rect 14364 39526 14420 39564
rect 15036 40292 15092 40302
rect 15036 39618 15092 40236
rect 15932 40292 15988 40462
rect 15932 40226 15988 40236
rect 15036 39566 15038 39618
rect 15090 39566 15092 39618
rect 15036 39554 15092 39566
rect 15484 40178 15540 40190
rect 15484 40126 15486 40178
rect 15538 40126 15540 40178
rect 15372 39508 15428 39518
rect 14812 39396 14868 39406
rect 15260 39396 15316 39406
rect 14812 39394 14980 39396
rect 14812 39342 14814 39394
rect 14866 39342 14980 39394
rect 14812 39340 14980 39342
rect 14812 39330 14868 39340
rect 14140 39116 14868 39172
rect 14364 38948 14420 38958
rect 14364 38834 14420 38892
rect 14364 38782 14366 38834
rect 14418 38782 14420 38834
rect 14364 38770 14420 38782
rect 13804 38724 13860 38734
rect 13804 38630 13860 38668
rect 14812 38162 14868 39116
rect 14924 38836 14980 39340
rect 15260 39302 15316 39340
rect 15372 39172 15428 39452
rect 15260 39116 15428 39172
rect 15036 38836 15092 38846
rect 14924 38780 15036 38836
rect 15036 38770 15092 38780
rect 15260 38834 15316 39116
rect 15260 38782 15262 38834
rect 15314 38782 15316 38834
rect 14812 38110 14814 38162
rect 14866 38110 14868 38162
rect 14812 38098 14868 38110
rect 13692 37998 13694 38050
rect 13746 37998 13748 38050
rect 13692 37986 13748 37998
rect 15148 38050 15204 38062
rect 15148 37998 15150 38050
rect 15202 37998 15204 38050
rect 14252 37492 14308 37502
rect 13468 37490 13748 37492
rect 13468 37438 13470 37490
rect 13522 37438 13748 37490
rect 13468 37436 13748 37438
rect 13468 37426 13524 37436
rect 10108 35870 10110 35922
rect 10162 35870 10164 35922
rect 10108 35858 10164 35870
rect 10668 36204 10780 36260
rect 10668 35698 10724 36204
rect 10780 36194 10836 36204
rect 10668 35646 10670 35698
rect 10722 35646 10724 35698
rect 10668 35634 10724 35646
rect 8540 35588 8596 35598
rect 8204 35364 8260 35374
rect 8204 34804 8260 35308
rect 8204 34738 8260 34748
rect 8540 34804 8596 35532
rect 9212 35140 9268 35150
rect 9212 35046 9268 35084
rect 8540 34738 8596 34748
rect 9884 34804 9940 34814
rect 8316 34692 8372 34702
rect 8428 34692 8484 34702
rect 8372 34690 8484 34692
rect 8372 34638 8430 34690
rect 8482 34638 8484 34690
rect 8372 34636 8484 34638
rect 8316 34354 8372 34636
rect 8428 34626 8484 34636
rect 8316 34302 8318 34354
rect 8370 34302 8372 34354
rect 8316 34290 8372 34302
rect 9100 34132 9156 34142
rect 9660 34132 9716 34142
rect 9100 34130 9716 34132
rect 9100 34078 9102 34130
rect 9154 34078 9662 34130
rect 9714 34078 9716 34130
rect 9100 34076 9716 34078
rect 9100 34066 9156 34076
rect 9660 34066 9716 34076
rect 9548 33908 9604 33918
rect 9548 33814 9604 33852
rect 9548 33236 9604 33246
rect 8652 33124 8708 33134
rect 8540 32788 8596 32798
rect 8540 32694 8596 32732
rect 8652 32674 8708 33068
rect 8652 32622 8654 32674
rect 8706 32622 8708 32674
rect 8652 32610 8708 32622
rect 9548 33122 9604 33180
rect 9548 33070 9550 33122
rect 9602 33070 9604 33122
rect 7644 31892 8036 31948
rect 9548 31948 9604 33070
rect 9548 31892 9716 31948
rect 7420 31778 7476 31790
rect 7420 31726 7422 31778
rect 7474 31726 7476 31778
rect 7420 31220 7476 31726
rect 7420 31154 7476 31164
rect 6636 24894 6638 24946
rect 6690 24894 6692 24946
rect 6636 24882 6692 24894
rect 7196 24892 7364 24948
rect 7644 24948 7700 31892
rect 9660 31666 9716 31892
rect 9660 31614 9662 31666
rect 9714 31614 9716 31666
rect 9660 31602 9716 31614
rect 8316 31556 8372 31566
rect 8204 31220 8260 31230
rect 8204 31126 8260 31164
rect 8316 31106 8372 31500
rect 8316 31054 8318 31106
rect 8370 31054 8372 31106
rect 8316 31042 8372 31054
rect 9212 31556 9268 31566
rect 9212 28866 9268 31500
rect 9212 28814 9214 28866
rect 9266 28814 9268 28866
rect 9212 28802 9268 28814
rect 8540 28530 8596 28542
rect 8540 28478 8542 28530
rect 8594 28478 8596 28530
rect 7868 28418 7924 28430
rect 7868 28366 7870 28418
rect 7922 28366 7924 28418
rect 7756 27970 7812 27982
rect 7756 27918 7758 27970
rect 7810 27918 7812 27970
rect 7756 26292 7812 27918
rect 7868 27074 7924 28366
rect 7868 27022 7870 27074
rect 7922 27022 7924 27074
rect 7868 27010 7924 27022
rect 8092 27074 8148 27086
rect 8092 27022 8094 27074
rect 8146 27022 8148 27074
rect 7756 26226 7812 26236
rect 8092 26066 8148 27022
rect 8092 26014 8094 26066
rect 8146 26014 8148 26066
rect 8092 26002 8148 26014
rect 8204 26292 8260 26302
rect 8092 25844 8148 25854
rect 7756 25508 7812 25518
rect 7756 25414 7812 25452
rect 7644 24892 7924 24948
rect 4284 23938 4340 24780
rect 4844 24834 5460 24836
rect 4844 24782 5070 24834
rect 5122 24782 5460 24834
rect 4844 24780 5460 24782
rect 6972 24836 7028 24846
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 23886 4286 23938
rect 4338 23886 4340 23938
rect 4284 23874 4340 23886
rect 4732 23716 4788 23726
rect 4284 23714 4788 23716
rect 4284 23662 4734 23714
rect 4786 23662 4788 23714
rect 4284 23660 4788 23662
rect 2044 22430 2046 22482
rect 2098 22430 2100 22482
rect 2044 22418 2100 22430
rect 2380 23154 2436 23166
rect 2380 23102 2382 23154
rect 2434 23102 2436 23154
rect 2380 23044 2436 23102
rect 1708 21756 2100 21812
rect 1708 21588 1764 21598
rect 1708 20132 1764 21532
rect 1708 20038 1764 20076
rect 1820 20916 1876 20926
rect 1820 19460 1876 20860
rect 2044 20356 2100 21756
rect 2156 21588 2212 21598
rect 2380 21588 2436 22988
rect 2716 22932 2772 22942
rect 2156 21586 2436 21588
rect 2156 21534 2158 21586
rect 2210 21534 2436 21586
rect 2156 21532 2436 21534
rect 2492 21586 2548 21598
rect 2492 21534 2494 21586
rect 2546 21534 2548 21586
rect 2156 21522 2212 21532
rect 2044 20300 2212 20356
rect 1708 19404 1876 19460
rect 1932 20244 1988 20254
rect 1708 18564 1764 19404
rect 1708 18450 1764 18508
rect 1708 18398 1710 18450
rect 1762 18398 1764 18450
rect 1708 18386 1764 18398
rect 1820 19234 1876 19246
rect 1820 19182 1822 19234
rect 1874 19182 1876 19234
rect 1820 18900 1876 19182
rect 1932 19124 1988 20188
rect 2044 20130 2100 20142
rect 2044 20078 2046 20130
rect 2098 20078 2100 20130
rect 2044 19796 2100 20078
rect 2044 19730 2100 19740
rect 1932 19058 1988 19068
rect 1708 18228 1764 18238
rect 1708 17780 1764 18172
rect 1708 17666 1764 17724
rect 1708 17614 1710 17666
rect 1762 17614 1764 17666
rect 1708 17602 1764 17614
rect 1708 17444 1764 17454
rect 1708 16882 1764 17388
rect 1708 16830 1710 16882
rect 1762 16830 1764 16882
rect 1708 16818 1764 16830
rect 1820 16210 1876 18844
rect 2156 18788 2212 20300
rect 2380 20020 2436 20030
rect 2492 20020 2548 21534
rect 2716 20914 2772 22876
rect 4284 22370 4340 23660
rect 4732 23650 4788 23660
rect 4844 23378 4900 24780
rect 5068 24770 5124 24780
rect 6972 24742 7028 24780
rect 6412 24722 6468 24734
rect 6412 24670 6414 24722
rect 6466 24670 6468 24722
rect 5852 24612 5908 24622
rect 5852 24518 5908 24556
rect 4844 23326 4846 23378
rect 4898 23326 4900 23378
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4284 22318 4286 22370
rect 4338 22318 4340 22370
rect 4284 22306 4340 22318
rect 4732 22372 4788 22382
rect 4732 22278 4788 22316
rect 2716 20862 2718 20914
rect 2770 20862 2772 20914
rect 2716 20850 2772 20862
rect 4284 22148 4340 22158
rect 4284 20802 4340 22092
rect 4844 21810 4900 23326
rect 4956 23938 5012 23950
rect 5628 23940 5684 23950
rect 4956 23886 4958 23938
rect 5010 23886 5012 23938
rect 4956 23380 5012 23886
rect 4956 23314 5012 23324
rect 5068 23938 5684 23940
rect 5068 23886 5630 23938
rect 5682 23886 5684 23938
rect 5068 23884 5684 23886
rect 5068 22258 5124 23884
rect 5628 23874 5684 23884
rect 6188 23828 6244 23838
rect 5852 23380 5908 23390
rect 5852 23286 5908 23324
rect 5516 23156 5572 23166
rect 6188 23156 6244 23772
rect 6412 23380 6468 24670
rect 6636 23716 6692 23726
rect 6636 23622 6692 23660
rect 6412 23314 6468 23324
rect 6972 23492 7028 23502
rect 5516 23154 6244 23156
rect 5516 23102 5518 23154
rect 5570 23102 6190 23154
rect 6242 23102 6244 23154
rect 5516 23100 6244 23102
rect 5516 23090 5572 23100
rect 6188 23090 6244 23100
rect 6860 23268 6916 23278
rect 6860 23154 6916 23212
rect 6972 23266 7028 23436
rect 6972 23214 6974 23266
rect 7026 23214 7028 23266
rect 6972 23202 7028 23214
rect 6860 23102 6862 23154
rect 6914 23102 6916 23154
rect 5964 22372 6020 22382
rect 6300 22372 6356 22382
rect 5964 22278 6020 22316
rect 6076 22370 6356 22372
rect 6076 22318 6302 22370
rect 6354 22318 6356 22370
rect 6076 22316 6356 22318
rect 5068 22206 5070 22258
rect 5122 22206 5124 22258
rect 5068 22194 5124 22206
rect 6076 21924 6132 22316
rect 6300 22306 6356 22316
rect 6412 22372 6468 22382
rect 4844 21758 4846 21810
rect 4898 21758 4900 21810
rect 4844 21746 4900 21758
rect 5628 21868 6132 21924
rect 5628 21810 5684 21868
rect 5628 21758 5630 21810
rect 5682 21758 5684 21810
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4284 20750 4286 20802
rect 4338 20750 4340 20802
rect 4284 20738 4340 20750
rect 4732 20578 4788 20590
rect 4732 20526 4734 20578
rect 4786 20526 4788 20578
rect 4284 20468 4340 20478
rect 3164 20244 3220 20254
rect 2380 20018 2548 20020
rect 2380 19966 2382 20018
rect 2434 19966 2548 20018
rect 2380 19964 2548 19966
rect 2940 20018 2996 20030
rect 2940 19966 2942 20018
rect 2994 19966 2996 20018
rect 2268 19236 2324 19246
rect 2268 19142 2324 19180
rect 2044 18732 2156 18788
rect 2044 18004 2100 18732
rect 2156 18722 2212 18732
rect 2156 18564 2212 18574
rect 2156 18116 2212 18508
rect 2268 18340 2324 18350
rect 2268 18246 2324 18284
rect 2156 18060 2324 18116
rect 2044 17948 2212 18004
rect 2044 17444 2100 17454
rect 2044 17350 2100 17388
rect 2156 16882 2212 17948
rect 2156 16830 2158 16882
rect 2210 16830 2212 16882
rect 2156 16818 2212 16830
rect 1820 16158 1822 16210
rect 1874 16158 1876 16210
rect 1820 16146 1876 16158
rect 2156 16324 2212 16334
rect 1820 15204 1876 15214
rect 1820 13748 1876 15148
rect 1820 13746 2100 13748
rect 1820 13694 1822 13746
rect 1874 13694 2100 13746
rect 1820 13692 2100 13694
rect 1820 13682 1876 13692
rect 2044 13524 2100 13692
rect 2156 13746 2212 16268
rect 2268 16210 2324 18060
rect 2380 17892 2436 19964
rect 2940 19460 2996 19966
rect 2604 19124 2660 19134
rect 2604 19030 2660 19068
rect 2940 18450 2996 19404
rect 3164 19346 3220 20188
rect 4172 19908 4228 19918
rect 3164 19294 3166 19346
rect 3218 19294 3220 19346
rect 3164 19282 3220 19294
rect 3500 19572 3556 19582
rect 3500 19236 3556 19516
rect 2940 18398 2942 18450
rect 2994 18398 2996 18450
rect 2940 18386 2996 18398
rect 3276 19234 3556 19236
rect 3276 19182 3502 19234
rect 3554 19182 3556 19234
rect 3276 19180 3556 19182
rect 2380 17826 2436 17836
rect 3276 17778 3332 19180
rect 3500 19170 3556 19180
rect 3836 19012 3892 19022
rect 3836 18918 3892 18956
rect 3388 18452 3444 18462
rect 3388 18358 3444 18396
rect 4060 17892 4116 17902
rect 4060 17798 4116 17836
rect 3276 17726 3278 17778
rect 3330 17726 3332 17778
rect 3276 17714 3332 17726
rect 4172 17778 4228 19852
rect 4172 17726 4174 17778
rect 4226 17726 4228 17778
rect 4172 17714 4228 17726
rect 3500 17668 3556 17678
rect 3500 17574 3556 17612
rect 2380 17554 2436 17566
rect 2380 17502 2382 17554
rect 2434 17502 2436 17554
rect 2380 16884 2436 17502
rect 3612 17556 3668 17566
rect 3612 17462 3668 17500
rect 2716 17444 2772 17454
rect 2716 17350 2772 17388
rect 4172 17220 4228 17230
rect 2436 16828 2772 16884
rect 2380 16818 2436 16828
rect 2268 16158 2270 16210
rect 2322 16158 2324 16210
rect 2268 16146 2324 16158
rect 2716 16210 2772 16828
rect 3500 16324 3556 16334
rect 3500 16230 3556 16268
rect 2716 16158 2718 16210
rect 2770 16158 2772 16210
rect 2716 16146 2772 16158
rect 3612 15988 3668 15998
rect 3612 15986 3780 15988
rect 3612 15934 3614 15986
rect 3666 15934 3780 15986
rect 3612 15932 3780 15934
rect 3612 15922 3668 15932
rect 3500 15204 3556 15214
rect 3500 15110 3556 15148
rect 3612 15202 3668 15214
rect 3612 15150 3614 15202
rect 3666 15150 3668 15202
rect 2156 13694 2158 13746
rect 2210 13694 2212 13746
rect 2156 13682 2212 13694
rect 3612 13524 3668 15150
rect 3724 13972 3780 15932
rect 4172 13972 4228 17164
rect 4284 15426 4340 20412
rect 4732 20188 4788 20526
rect 5068 20580 5124 20590
rect 5068 20486 5124 20524
rect 4732 20132 4900 20188
rect 5292 20132 5348 20142
rect 4844 20130 5348 20132
rect 4844 20078 5294 20130
rect 5346 20078 5348 20130
rect 4844 20076 5348 20078
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4508 19460 4564 19470
rect 4508 19366 4564 19404
rect 4844 19460 4900 20076
rect 5292 20066 5348 20076
rect 5628 19908 5684 21758
rect 6300 21812 6356 21822
rect 6412 21812 6468 22316
rect 6300 21810 6468 21812
rect 6300 21758 6302 21810
rect 6354 21758 6468 21810
rect 6300 21756 6468 21758
rect 6860 22370 6916 23102
rect 6860 22318 6862 22370
rect 6914 22318 6916 22370
rect 6300 21746 6356 21756
rect 6860 21698 6916 22318
rect 7084 22260 7140 22270
rect 7084 22166 7140 22204
rect 6860 21646 6862 21698
rect 6914 21646 6916 21698
rect 6860 21634 6916 21646
rect 6636 21364 6692 21374
rect 6412 21362 6692 21364
rect 6412 21310 6638 21362
rect 6690 21310 6692 21362
rect 6412 21308 6692 21310
rect 6300 20804 6356 20814
rect 6300 20710 6356 20748
rect 5964 20578 6020 20590
rect 5964 20526 5966 20578
rect 6018 20526 6020 20578
rect 5964 20468 6020 20526
rect 6412 20468 6468 21308
rect 6636 21298 6692 21308
rect 6860 20802 6916 20814
rect 6860 20750 6862 20802
rect 6914 20750 6916 20802
rect 5964 20402 6020 20412
rect 6076 20412 6468 20468
rect 6636 20580 6692 20590
rect 5628 19842 5684 19852
rect 6076 20242 6132 20412
rect 6076 20190 6078 20242
rect 6130 20190 6132 20242
rect 4620 19348 4676 19358
rect 4620 19254 4676 19292
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4620 17780 4676 17790
rect 4620 17686 4676 17724
rect 4732 17108 4788 17118
rect 4844 17108 4900 19404
rect 6076 19348 6132 20190
rect 6636 20188 6692 20524
rect 6860 20468 6916 20750
rect 6860 20402 6916 20412
rect 6076 19282 6132 19292
rect 6188 20132 6692 20188
rect 7196 20188 7252 24892
rect 7308 24724 7364 24734
rect 7756 24724 7812 24734
rect 7308 24722 7812 24724
rect 7308 24670 7310 24722
rect 7362 24670 7758 24722
rect 7810 24670 7812 24722
rect 7308 24668 7812 24670
rect 7308 24658 7364 24668
rect 7756 24658 7812 24668
rect 7644 23380 7700 23390
rect 7644 23286 7700 23324
rect 7868 22372 7924 24892
rect 8092 24722 8148 25788
rect 8204 25396 8260 26236
rect 8540 26180 8596 28478
rect 8988 28532 9044 28542
rect 8988 28530 9492 28532
rect 8988 28478 8990 28530
rect 9042 28478 9492 28530
rect 8988 28476 9492 28478
rect 8988 28466 9044 28476
rect 8876 27636 8932 27646
rect 8540 26114 8596 26124
rect 8652 27634 8932 27636
rect 8652 27582 8878 27634
rect 8930 27582 8932 27634
rect 8652 27580 8932 27582
rect 8652 26292 8708 27580
rect 8876 27570 8932 27580
rect 8652 26178 8708 26236
rect 8652 26126 8654 26178
rect 8706 26126 8708 26178
rect 8652 26114 8708 26126
rect 9212 26068 9268 26078
rect 9212 25506 9268 26012
rect 9212 25454 9214 25506
rect 9266 25454 9268 25506
rect 9212 25442 9268 25454
rect 8540 25396 8596 25406
rect 8204 25394 8596 25396
rect 8204 25342 8542 25394
rect 8594 25342 8596 25394
rect 8204 25340 8596 25342
rect 8540 25330 8596 25340
rect 8876 25396 8932 25406
rect 8876 25394 9156 25396
rect 8876 25342 8878 25394
rect 8930 25342 9156 25394
rect 8876 25340 9156 25342
rect 8876 25330 8932 25340
rect 8092 24670 8094 24722
rect 8146 24670 8148 24722
rect 8092 24658 8148 24670
rect 8428 24836 8484 24846
rect 7980 24612 8036 24622
rect 7980 23154 8036 24556
rect 7980 23102 7982 23154
rect 8034 23102 8036 23154
rect 7980 23090 8036 23102
rect 8428 23154 8484 24780
rect 8876 24834 8932 24846
rect 8876 24782 8878 24834
rect 8930 24782 8932 24834
rect 8876 24612 8932 24782
rect 8876 24546 8932 24556
rect 8652 23828 8708 23838
rect 8988 23828 9044 23838
rect 8652 23734 8708 23772
rect 8764 23772 8988 23828
rect 8428 23102 8430 23154
rect 8482 23102 8484 23154
rect 8428 23090 8484 23102
rect 8540 23714 8596 23726
rect 8540 23662 8542 23714
rect 8594 23662 8596 23714
rect 8540 23044 8596 23662
rect 8764 23266 8820 23772
rect 8988 23762 9044 23772
rect 9100 23604 9156 25340
rect 9436 24836 9492 28476
rect 9548 28420 9604 28430
rect 9548 28326 9604 28364
rect 9548 27970 9604 27982
rect 9548 27918 9550 27970
rect 9602 27918 9604 27970
rect 9548 27076 9604 27918
rect 9548 27010 9604 27020
rect 9772 27858 9828 27870
rect 9772 27806 9774 27858
rect 9826 27806 9828 27858
rect 9660 26516 9716 26526
rect 9772 26516 9828 27806
rect 9884 27412 9940 34748
rect 11116 34802 11172 36428
rect 11228 37266 11284 37278
rect 11228 37214 11230 37266
rect 11282 37214 11284 37266
rect 11228 36260 11284 37214
rect 12908 36596 12964 36606
rect 13692 36596 13748 37436
rect 12908 36594 13076 36596
rect 12908 36542 12910 36594
rect 12962 36542 13076 36594
rect 12908 36540 13076 36542
rect 12908 36530 12964 36540
rect 11228 36194 11284 36204
rect 12908 36148 12964 36158
rect 12908 35698 12964 36092
rect 12908 35646 12910 35698
rect 12962 35646 12964 35698
rect 12908 35634 12964 35646
rect 13020 35028 13076 36540
rect 13468 36540 13692 36596
rect 13468 35698 13524 36540
rect 13692 36502 13748 36540
rect 14252 36482 14308 37436
rect 14700 37492 14756 37502
rect 15148 37492 15204 37998
rect 14700 37398 14756 37436
rect 14924 37436 15204 37492
rect 14588 37268 14644 37278
rect 14476 37212 14588 37268
rect 14252 36430 14254 36482
rect 14306 36430 14308 36482
rect 14252 36418 14308 36430
rect 14364 37154 14420 37166
rect 14364 37102 14366 37154
rect 14418 37102 14420 37154
rect 14364 36036 14420 37102
rect 14364 35970 14420 35980
rect 13468 35646 13470 35698
rect 13522 35646 13524 35698
rect 13468 35634 13524 35646
rect 14476 35252 14532 37212
rect 14588 37202 14644 37212
rect 13020 34962 13076 34972
rect 14364 35196 14532 35252
rect 14588 35474 14644 35486
rect 14588 35422 14590 35474
rect 14642 35422 14644 35474
rect 11116 34750 11118 34802
rect 11170 34750 11172 34802
rect 11116 34738 11172 34750
rect 11452 34802 11508 34814
rect 11452 34750 11454 34802
rect 11506 34750 11508 34802
rect 10780 34130 10836 34142
rect 10780 34078 10782 34130
rect 10834 34078 10836 34130
rect 10556 33460 10612 33470
rect 10556 33346 10612 33404
rect 10556 33294 10558 33346
rect 10610 33294 10612 33346
rect 10556 33282 10612 33294
rect 10332 33236 10388 33246
rect 10332 33142 10388 33180
rect 10108 33124 10164 33134
rect 10108 33030 10164 33068
rect 10556 32452 10612 32462
rect 10444 31556 10500 31566
rect 10444 31462 10500 31500
rect 10108 28532 10164 28542
rect 10108 28438 10164 28476
rect 9884 27346 9940 27356
rect 9996 28418 10052 28430
rect 9996 28366 9998 28418
rect 10050 28366 10052 28418
rect 9996 26964 10052 28366
rect 10444 28420 10500 28430
rect 10220 28084 10276 28094
rect 10220 27990 10276 28028
rect 10444 27858 10500 28364
rect 10444 27806 10446 27858
rect 10498 27806 10500 27858
rect 10444 27794 10500 27806
rect 9996 26870 10052 26908
rect 10556 26628 10612 32396
rect 10780 30212 10836 34078
rect 11340 34130 11396 34142
rect 11340 34078 11342 34130
rect 11394 34078 11396 34130
rect 11340 33460 11396 34078
rect 11340 33394 11396 33404
rect 11452 31948 11508 34750
rect 13692 34242 13748 34254
rect 13692 34190 13694 34242
rect 13746 34190 13748 34242
rect 12796 33572 12852 33582
rect 12796 32786 12852 33516
rect 12796 32734 12798 32786
rect 12850 32734 12852 32786
rect 12796 32722 12852 32734
rect 13356 33460 13412 33470
rect 11676 32676 11732 32686
rect 11564 32452 11620 32462
rect 11564 32358 11620 32396
rect 11228 31892 11508 31948
rect 11228 31668 11284 31892
rect 11340 31780 11396 31790
rect 11564 31780 11620 31790
rect 11340 31778 11564 31780
rect 11340 31726 11342 31778
rect 11394 31726 11564 31778
rect 11340 31724 11564 31726
rect 11340 31714 11396 31724
rect 11564 31686 11620 31724
rect 11228 31602 11284 31612
rect 10780 29426 10836 30156
rect 10780 29374 10782 29426
rect 10834 29374 10836 29426
rect 10780 29362 10836 29374
rect 11676 29092 11732 32620
rect 12236 32674 12292 32686
rect 12236 32622 12238 32674
rect 12290 32622 12292 32674
rect 12012 32562 12068 32574
rect 12012 32510 12014 32562
rect 12066 32510 12068 32562
rect 12012 32452 12068 32510
rect 12012 32386 12068 32396
rect 12236 31780 12292 32622
rect 12572 32564 12628 32574
rect 12572 32470 12628 32508
rect 13356 32562 13412 33404
rect 13356 32510 13358 32562
rect 13410 32510 13412 32562
rect 13356 32498 13412 32510
rect 13468 33346 13524 33358
rect 13468 33294 13470 33346
rect 13522 33294 13524 33346
rect 12908 32228 12964 32238
rect 12348 31892 12404 31902
rect 12908 31892 12964 32172
rect 12348 31890 12964 31892
rect 12348 31838 12350 31890
rect 12402 31838 12964 31890
rect 12348 31836 12964 31838
rect 12348 31826 12404 31836
rect 11900 31668 11956 31678
rect 11900 31574 11956 31612
rect 12236 31220 12292 31724
rect 12796 31554 12852 31566
rect 12796 31502 12798 31554
rect 12850 31502 12852 31554
rect 12236 31164 12404 31220
rect 12236 30996 12292 31006
rect 11676 29026 11732 29036
rect 12012 30882 12068 30894
rect 12012 30830 12014 30882
rect 12066 30830 12068 30882
rect 12012 28866 12068 30830
rect 12124 30212 12180 30222
rect 12124 30118 12180 30156
rect 12012 28814 12014 28866
rect 12066 28814 12068 28866
rect 12012 28802 12068 28814
rect 11676 28644 11732 28654
rect 11676 28642 11844 28644
rect 11676 28590 11678 28642
rect 11730 28590 11844 28642
rect 11676 28588 11844 28590
rect 11676 28578 11732 28588
rect 11452 28532 11508 28542
rect 11452 27300 11508 28476
rect 11564 27300 11620 27310
rect 11452 27298 11620 27300
rect 11452 27246 11566 27298
rect 11618 27246 11620 27298
rect 11452 27244 11620 27246
rect 11564 27234 11620 27244
rect 11340 27076 11396 27086
rect 11676 27076 11732 27086
rect 11340 27074 11732 27076
rect 11340 27022 11342 27074
rect 11394 27022 11678 27074
rect 11730 27022 11732 27074
rect 11340 27020 11732 27022
rect 11340 27010 11396 27020
rect 11676 27010 11732 27020
rect 11788 27076 11844 28588
rect 11788 27010 11844 27020
rect 11004 26962 11060 26974
rect 11004 26910 11006 26962
rect 11058 26910 11060 26962
rect 10668 26852 10724 26862
rect 10668 26850 10948 26852
rect 10668 26798 10670 26850
rect 10722 26798 10948 26850
rect 10668 26796 10948 26798
rect 10668 26786 10724 26796
rect 9660 26514 9828 26516
rect 9660 26462 9662 26514
rect 9714 26462 9828 26514
rect 9660 26460 9828 26462
rect 10332 26572 10612 26628
rect 9660 26450 9716 26460
rect 10220 26404 10276 26414
rect 10108 26348 10220 26404
rect 9996 26292 10052 26302
rect 9996 26198 10052 26236
rect 9996 26068 10052 26078
rect 9884 26012 9996 26068
rect 9548 24836 9604 24846
rect 9436 24834 9604 24836
rect 9436 24782 9550 24834
rect 9602 24782 9604 24834
rect 9436 24780 9604 24782
rect 9100 23548 9380 23604
rect 8764 23214 8766 23266
rect 8818 23214 8820 23266
rect 8764 23202 8820 23214
rect 8540 22978 8596 22988
rect 9324 22596 9380 23548
rect 9436 23268 9492 24780
rect 9548 24770 9604 24780
rect 9660 23828 9716 23838
rect 9660 23734 9716 23772
rect 9884 23492 9940 26012
rect 9996 26002 10052 26012
rect 9996 25394 10052 25406
rect 9996 25342 9998 25394
rect 10050 25342 10052 25394
rect 9996 24724 10052 25342
rect 10108 24946 10164 26348
rect 10220 26310 10276 26348
rect 10108 24894 10110 24946
rect 10162 24894 10164 24946
rect 10108 24882 10164 24894
rect 9996 24658 10052 24668
rect 9436 23202 9492 23212
rect 9660 23436 9940 23492
rect 10108 23938 10164 23950
rect 10108 23886 10110 23938
rect 10162 23886 10164 23938
rect 9660 23266 9716 23436
rect 9660 23214 9662 23266
rect 9714 23214 9716 23266
rect 9660 23202 9716 23214
rect 9884 23268 9940 23278
rect 9548 22596 9604 22606
rect 9324 22594 9604 22596
rect 9324 22542 9550 22594
rect 9602 22542 9604 22594
rect 9324 22540 9604 22542
rect 9548 22530 9604 22540
rect 9884 22594 9940 23212
rect 10108 23156 10164 23886
rect 10108 23154 10276 23156
rect 10108 23102 10110 23154
rect 10162 23102 10276 23154
rect 10108 23100 10276 23102
rect 10108 23090 10164 23100
rect 9884 22542 9886 22594
rect 9938 22542 9940 22594
rect 9884 22530 9940 22542
rect 8428 22372 8484 22382
rect 7868 22370 8148 22372
rect 7868 22318 7870 22370
rect 7922 22318 8148 22370
rect 7868 22316 8148 22318
rect 7868 22306 7924 22316
rect 7532 22146 7588 22158
rect 7532 22094 7534 22146
rect 7586 22094 7588 22146
rect 7420 21700 7476 21710
rect 7420 21606 7476 21644
rect 7532 21588 7588 22094
rect 8092 21812 8148 22316
rect 8428 22278 8484 22316
rect 8204 22148 8260 22158
rect 8204 22054 8260 22092
rect 10220 22036 10276 23100
rect 8092 21718 8148 21756
rect 10108 21980 10276 22036
rect 7532 20804 7588 21532
rect 7532 20738 7588 20748
rect 7644 20802 7700 20814
rect 7644 20750 7646 20802
rect 7698 20750 7700 20802
rect 7644 20468 7700 20750
rect 8428 20692 8484 20702
rect 8428 20690 9604 20692
rect 8428 20638 8430 20690
rect 8482 20638 9604 20690
rect 8428 20636 9604 20638
rect 8428 20626 8484 20636
rect 7644 20402 7700 20412
rect 9548 20242 9604 20636
rect 9548 20190 9550 20242
rect 9602 20190 9604 20242
rect 7196 20132 7364 20188
rect 9548 20178 9604 20190
rect 9884 20580 9940 20590
rect 8540 20132 8596 20142
rect 5628 19234 5684 19246
rect 5628 19182 5630 19234
rect 5682 19182 5684 19234
rect 5068 19124 5124 19134
rect 5068 19122 5348 19124
rect 5068 19070 5070 19122
rect 5122 19070 5348 19122
rect 5068 19068 5348 19070
rect 5068 19058 5124 19068
rect 4956 19010 5012 19022
rect 4956 18958 4958 19010
rect 5010 18958 5012 19010
rect 4956 18788 5012 18958
rect 4956 18722 5012 18732
rect 4732 17106 4900 17108
rect 4732 17054 4734 17106
rect 4786 17054 4900 17106
rect 4732 17052 4900 17054
rect 4956 18452 5012 18462
rect 4956 17890 5012 18396
rect 5180 18228 5236 18238
rect 4956 17838 4958 17890
rect 5010 17838 5012 17890
rect 4732 17042 4788 17052
rect 4956 16996 5012 17838
rect 5068 18172 5180 18228
rect 5068 17778 5124 18172
rect 5180 18162 5236 18172
rect 5068 17726 5070 17778
rect 5122 17726 5124 17778
rect 5068 17714 5124 17726
rect 5292 17106 5348 19068
rect 5628 18562 5684 19182
rect 5628 18510 5630 18562
rect 5682 18510 5684 18562
rect 5292 17054 5294 17106
rect 5346 17054 5348 17106
rect 5292 17042 5348 17054
rect 5516 17666 5572 17678
rect 5516 17614 5518 17666
rect 5570 17614 5572 17666
rect 4956 16940 5236 16996
rect 5180 16884 5236 16940
rect 5404 16884 5460 16894
rect 5180 16882 5460 16884
rect 5180 16830 5406 16882
rect 5458 16830 5460 16882
rect 5180 16828 5460 16830
rect 5404 16818 5460 16828
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 5516 16324 5572 17614
rect 5628 17220 5684 18510
rect 6188 19010 6244 20132
rect 6412 20020 6468 20030
rect 6412 19926 6468 19964
rect 7196 19460 7252 19470
rect 6748 19348 6804 19358
rect 6636 19124 6692 19134
rect 6636 19030 6692 19068
rect 6188 18958 6190 19010
rect 6242 18958 6244 19010
rect 6076 17668 6132 17678
rect 6076 17574 6132 17612
rect 5628 17154 5684 17164
rect 6188 17220 6244 18958
rect 6748 18340 6804 19292
rect 7196 19234 7252 19404
rect 7196 19182 7198 19234
rect 7250 19182 7252 19234
rect 7196 19170 7252 19182
rect 6748 18274 6804 18284
rect 6412 18228 6468 18238
rect 6412 18134 6468 18172
rect 7308 18228 7364 20132
rect 7980 20130 8596 20132
rect 7980 20078 8542 20130
rect 8594 20078 8596 20130
rect 7980 20076 8596 20078
rect 7980 19346 8036 20076
rect 8540 20066 8596 20076
rect 9884 20130 9940 20524
rect 9884 20078 9886 20130
rect 9938 20078 9940 20130
rect 9884 20066 9940 20078
rect 8876 20020 8932 20030
rect 8876 19926 8932 19964
rect 7980 19294 7982 19346
rect 8034 19294 8036 19346
rect 7980 19282 8036 19294
rect 8764 19796 8820 19806
rect 8316 18562 8372 18574
rect 8316 18510 8318 18562
rect 8370 18510 8372 18562
rect 7308 18162 7364 18172
rect 8092 18450 8148 18462
rect 8092 18398 8094 18450
rect 8146 18398 8148 18450
rect 8092 17892 8148 18398
rect 8092 17826 8148 17836
rect 6188 17154 6244 17164
rect 8316 16996 8372 18510
rect 8764 18450 8820 19740
rect 10108 19572 10164 21980
rect 10220 21812 10276 21822
rect 10220 21364 10276 21756
rect 10220 21298 10276 21308
rect 10332 20188 10388 26572
rect 10668 26402 10724 26414
rect 10668 26350 10670 26402
rect 10722 26350 10724 26402
rect 10556 25172 10612 25182
rect 10556 23940 10612 25116
rect 10668 24388 10724 26350
rect 10892 25396 10948 26796
rect 11004 26404 11060 26910
rect 11116 26964 11172 26974
rect 11116 26870 11172 26908
rect 11004 26338 11060 26348
rect 11676 26404 11732 26414
rect 11676 26292 11732 26348
rect 11676 26290 12180 26292
rect 11676 26238 11678 26290
rect 11730 26238 12180 26290
rect 11676 26236 12180 26238
rect 11676 26226 11732 26236
rect 10780 25284 10836 25294
rect 10780 24946 10836 25228
rect 10780 24894 10782 24946
rect 10834 24894 10836 24946
rect 10780 24882 10836 24894
rect 10892 24724 10948 25340
rect 11340 26178 11396 26190
rect 11340 26126 11342 26178
rect 11394 26126 11396 26178
rect 11340 24836 11396 26126
rect 12124 25618 12180 26236
rect 12124 25566 12126 25618
rect 12178 25566 12180 25618
rect 12124 25554 12180 25566
rect 11340 24742 11396 24780
rect 11788 24834 11844 24846
rect 11788 24782 11790 24834
rect 11842 24782 11844 24834
rect 11116 24724 11172 24734
rect 10892 24722 11172 24724
rect 10892 24670 11118 24722
rect 11170 24670 11172 24722
rect 10892 24668 11172 24670
rect 11116 24658 11172 24668
rect 10780 24388 10836 24398
rect 10668 24332 10780 24388
rect 10444 23938 10612 23940
rect 10444 23886 10558 23938
rect 10610 23886 10612 23938
rect 10444 23884 10612 23886
rect 10444 23492 10500 23884
rect 10556 23874 10612 23884
rect 10668 23716 10724 23726
rect 10444 23426 10500 23436
rect 10556 23714 10724 23716
rect 10556 23662 10670 23714
rect 10722 23662 10724 23714
rect 10556 23660 10724 23662
rect 10444 23156 10500 23166
rect 10444 23062 10500 23100
rect 10444 22370 10500 22382
rect 10444 22318 10446 22370
rect 10498 22318 10500 22370
rect 10444 20916 10500 22318
rect 10556 22258 10612 23660
rect 10668 23650 10724 23660
rect 10668 23268 10724 23278
rect 10668 23174 10724 23212
rect 10780 23156 10836 24332
rect 10780 23090 10836 23100
rect 11116 23826 11172 23838
rect 11116 23774 11118 23826
rect 11170 23774 11172 23826
rect 11116 23154 11172 23774
rect 11788 23604 11844 24782
rect 11900 24612 11956 24622
rect 11900 23938 11956 24556
rect 11900 23886 11902 23938
rect 11954 23886 11956 23938
rect 11900 23874 11956 23886
rect 12012 24164 12068 24174
rect 11900 23604 11956 23614
rect 11788 23548 11900 23604
rect 11900 23538 11956 23548
rect 11900 23156 11956 23166
rect 12012 23156 12068 24108
rect 11116 23102 11118 23154
rect 11170 23102 11172 23154
rect 10556 22206 10558 22258
rect 10610 22206 10612 22258
rect 10556 22194 10612 22206
rect 10668 21588 10724 21598
rect 11004 21588 11060 21598
rect 10668 21586 11004 21588
rect 10668 21534 10670 21586
rect 10722 21534 11004 21586
rect 10668 21532 11004 21534
rect 10668 21522 10724 21532
rect 11004 21494 11060 21532
rect 10556 20916 10612 20926
rect 10444 20860 10556 20916
rect 10556 20822 10612 20860
rect 11004 20580 11060 20590
rect 11004 20486 11060 20524
rect 11116 20188 11172 23102
rect 11788 23154 12068 23156
rect 11788 23102 11902 23154
rect 11954 23102 12068 23154
rect 11788 23100 12068 23102
rect 11676 22596 11732 22606
rect 11676 22484 11732 22540
rect 11564 22482 11732 22484
rect 11564 22430 11678 22482
rect 11730 22430 11732 22482
rect 11564 22428 11732 22430
rect 11564 21810 11620 22428
rect 11676 22418 11732 22428
rect 11788 22260 11844 23100
rect 11900 23090 11956 23100
rect 12236 22820 12292 30940
rect 12348 27524 12404 31164
rect 12796 30100 12852 31502
rect 12908 30210 12964 31836
rect 13468 31780 13524 33294
rect 13580 32562 13636 32574
rect 13580 32510 13582 32562
rect 13634 32510 13636 32562
rect 13580 32228 13636 32510
rect 13692 32564 13748 34190
rect 13916 33460 13972 33470
rect 13916 33346 13972 33404
rect 13916 33294 13918 33346
rect 13970 33294 13972 33346
rect 13916 33282 13972 33294
rect 13692 32498 13748 32508
rect 13580 32162 13636 32172
rect 13692 32004 13748 32014
rect 13356 31724 13524 31780
rect 13580 31778 13636 31790
rect 13580 31726 13582 31778
rect 13634 31726 13636 31778
rect 13356 31444 13412 31724
rect 13580 31668 13636 31726
rect 13580 31602 13636 31612
rect 13356 31388 13524 31444
rect 13468 30994 13524 31388
rect 13468 30942 13470 30994
rect 13522 30942 13524 30994
rect 13468 30436 13524 30942
rect 12908 30158 12910 30210
rect 12962 30158 12964 30210
rect 12908 30146 12964 30158
rect 13356 30380 13524 30436
rect 13356 30212 13412 30380
rect 13356 30146 13412 30156
rect 13468 30210 13524 30222
rect 13468 30158 13470 30210
rect 13522 30158 13524 30210
rect 12796 30034 12852 30044
rect 13468 30100 13524 30158
rect 13468 30034 13524 30044
rect 12796 29314 12852 29326
rect 12796 29262 12798 29314
rect 12850 29262 12852 29314
rect 12348 27458 12404 27468
rect 12684 28642 12740 28654
rect 12684 28590 12686 28642
rect 12738 28590 12740 28642
rect 12684 27188 12740 28590
rect 12796 28530 12852 29262
rect 12796 28478 12798 28530
rect 12850 28478 12852 28530
rect 12796 28466 12852 28478
rect 13468 28084 13524 28094
rect 13692 28084 13748 31948
rect 13804 31554 13860 31566
rect 13804 31502 13806 31554
rect 13858 31502 13860 31554
rect 13804 30212 13860 31502
rect 14364 31108 14420 35196
rect 14588 35140 14644 35422
rect 14588 35074 14644 35084
rect 14476 35028 14532 35038
rect 14476 34916 14532 34972
rect 14588 34916 14644 34926
rect 14476 34914 14644 34916
rect 14476 34862 14590 34914
rect 14642 34862 14644 34914
rect 14476 34860 14644 34862
rect 14588 34850 14644 34860
rect 14924 34914 14980 37436
rect 15148 37380 15204 37436
rect 15148 37314 15204 37324
rect 15036 37266 15092 37278
rect 15036 37214 15038 37266
rect 15090 37214 15092 37266
rect 15036 37044 15092 37214
rect 15036 36978 15092 36988
rect 15260 37044 15316 38782
rect 15260 36978 15316 36988
rect 15372 38948 15428 38958
rect 14924 34862 14926 34914
rect 14978 34862 14980 34914
rect 14924 34850 14980 34862
rect 15148 36932 15204 36942
rect 15372 36932 15428 38892
rect 15484 38836 15540 40126
rect 15596 39620 15652 39630
rect 15596 39526 15652 39564
rect 15484 38770 15540 38780
rect 15596 38052 15652 38062
rect 15596 37958 15652 37996
rect 15820 37826 15876 37838
rect 15820 37774 15822 37826
rect 15874 37774 15876 37826
rect 15708 37268 15764 37278
rect 15708 37174 15764 37212
rect 15372 36876 15764 36932
rect 14476 33906 14532 33918
rect 14476 33854 14478 33906
rect 14530 33854 14532 33906
rect 14476 32900 14532 33854
rect 14476 32834 14532 32844
rect 14924 33460 14980 33470
rect 14700 32564 14756 32574
rect 14476 31556 14532 31566
rect 14476 31462 14532 31500
rect 14700 31556 14756 32508
rect 14700 31554 14868 31556
rect 14700 31502 14702 31554
rect 14754 31502 14868 31554
rect 14700 31500 14868 31502
rect 14700 31490 14756 31500
rect 14700 31108 14756 31118
rect 14364 31106 14756 31108
rect 14364 31054 14702 31106
rect 14754 31054 14756 31106
rect 14364 31052 14756 31054
rect 14028 30212 14084 30222
rect 13804 30210 14196 30212
rect 13804 30158 14030 30210
rect 14082 30158 14196 30210
rect 13804 30156 14196 30158
rect 14028 30146 14084 30156
rect 13916 29540 13972 29550
rect 13916 28530 13972 29484
rect 14140 29316 14196 30156
rect 14140 29250 14196 29260
rect 14140 29092 14196 29102
rect 14140 28644 14196 29036
rect 14140 28642 14308 28644
rect 14140 28590 14142 28642
rect 14194 28590 14308 28642
rect 14140 28588 14308 28590
rect 14140 28578 14196 28588
rect 13916 28478 13918 28530
rect 13970 28478 13972 28530
rect 13468 28082 13860 28084
rect 13468 28030 13470 28082
rect 13522 28030 13860 28082
rect 13468 28028 13860 28030
rect 13468 28018 13524 28028
rect 13244 27858 13300 27870
rect 13244 27806 13246 27858
rect 13298 27806 13300 27858
rect 13244 27300 13300 27806
rect 13804 27858 13860 28028
rect 13804 27806 13806 27858
rect 13858 27806 13860 27858
rect 13804 27794 13860 27806
rect 13916 27860 13972 28478
rect 14028 27860 14084 27870
rect 13916 27858 14084 27860
rect 13916 27806 14030 27858
rect 14082 27806 14084 27858
rect 13916 27804 14084 27806
rect 14028 27794 14084 27804
rect 13244 27234 13300 27244
rect 13692 27412 13748 27422
rect 12684 27122 12740 27132
rect 12460 25620 12516 25630
rect 12460 25394 12516 25564
rect 13692 25620 13748 27356
rect 13804 27300 13860 27310
rect 13804 27186 13860 27244
rect 13804 27134 13806 27186
rect 13858 27134 13860 27186
rect 13804 27122 13860 27134
rect 14252 26962 14308 28588
rect 14476 27074 14532 31052
rect 14700 31042 14756 31052
rect 14588 30212 14644 30222
rect 14812 30212 14868 31500
rect 14588 30210 14868 30212
rect 14588 30158 14590 30210
rect 14642 30158 14868 30210
rect 14588 30156 14868 30158
rect 14924 30322 14980 33404
rect 15036 33348 15092 33358
rect 15036 32004 15092 33292
rect 15036 31778 15092 31948
rect 15148 31892 15204 36876
rect 15484 36596 15540 36606
rect 15484 36502 15540 36540
rect 15260 36372 15316 36382
rect 15260 36278 15316 36316
rect 15372 36260 15428 36270
rect 15428 36204 15540 36260
rect 15372 36166 15428 36204
rect 15484 35922 15540 36204
rect 15484 35870 15486 35922
rect 15538 35870 15540 35922
rect 15484 35858 15540 35870
rect 15596 35476 15652 35486
rect 15372 34916 15428 34926
rect 15372 34822 15428 34860
rect 15596 34802 15652 35420
rect 15596 34750 15598 34802
rect 15650 34750 15652 34802
rect 15596 34738 15652 34750
rect 15596 34244 15652 34254
rect 15596 34150 15652 34188
rect 15148 31836 15540 31892
rect 15036 31726 15038 31778
rect 15090 31726 15092 31778
rect 15036 31714 15092 31726
rect 15372 31668 15428 31678
rect 15148 31612 15372 31668
rect 15036 31108 15092 31118
rect 15036 31014 15092 31052
rect 15148 30772 15204 31612
rect 15372 31574 15428 31612
rect 14924 30270 14926 30322
rect 14978 30270 14980 30322
rect 14588 28642 14644 30156
rect 14924 29652 14980 30270
rect 14924 29586 14980 29596
rect 15036 30716 15204 30772
rect 15372 31332 15428 31342
rect 15372 30994 15428 31276
rect 15372 30942 15374 30994
rect 15426 30942 15428 30994
rect 14924 29092 14980 29102
rect 14588 28590 14590 28642
rect 14642 28590 14644 28642
rect 14588 28578 14644 28590
rect 14812 29036 14924 29092
rect 14812 27300 14868 29036
rect 14924 29026 14980 29036
rect 14924 28868 14980 28878
rect 15036 28868 15092 30716
rect 14924 28866 15092 28868
rect 14924 28814 14926 28866
rect 14978 28814 15092 28866
rect 14924 28812 15092 28814
rect 14924 28802 14980 28812
rect 14812 27188 14868 27244
rect 14924 27188 14980 27198
rect 14812 27186 14980 27188
rect 14812 27134 14926 27186
rect 14978 27134 14980 27186
rect 14812 27132 14980 27134
rect 14924 27122 14980 27132
rect 14476 27022 14478 27074
rect 14530 27022 14532 27074
rect 14476 27010 14532 27022
rect 14252 26910 14254 26962
rect 14306 26910 14308 26962
rect 14252 26898 14308 26910
rect 15372 26908 15428 30942
rect 15484 30212 15540 31836
rect 15708 31792 15764 36876
rect 15820 36820 15876 37774
rect 15820 36754 15876 36764
rect 16044 37378 16100 40572
rect 16492 40516 16548 40526
rect 16548 40460 16660 40516
rect 16492 40450 16548 40460
rect 16268 40404 16324 40414
rect 16268 40402 16436 40404
rect 16268 40350 16270 40402
rect 16322 40350 16436 40402
rect 16268 40348 16436 40350
rect 16268 40338 16324 40348
rect 16156 40292 16212 40302
rect 16156 39618 16212 40236
rect 16156 39566 16158 39618
rect 16210 39566 16212 39618
rect 16156 39554 16212 39566
rect 16268 38836 16324 38846
rect 16268 38742 16324 38780
rect 16044 37326 16046 37378
rect 16098 37326 16100 37378
rect 15820 35812 15876 35822
rect 16044 35812 16100 37326
rect 16380 37268 16436 40348
rect 16492 38276 16548 38286
rect 16492 38050 16548 38220
rect 16492 37998 16494 38050
rect 16546 37998 16548 38050
rect 16492 37986 16548 37998
rect 16380 35924 16436 37212
rect 16492 37154 16548 37166
rect 16492 37102 16494 37154
rect 16546 37102 16548 37154
rect 16492 37044 16548 37102
rect 16492 36978 16548 36988
rect 16604 37156 16660 40460
rect 17388 40404 17444 40414
rect 17388 40310 17444 40348
rect 17500 39620 17556 40908
rect 17948 40740 18004 41804
rect 18508 41858 18564 41870
rect 18508 41806 18510 41858
rect 18562 41806 18564 41858
rect 18508 41188 18564 41806
rect 18508 41122 18564 41132
rect 19404 41188 19460 41198
rect 19292 41074 19348 41086
rect 19292 41022 19294 41074
rect 19346 41022 19348 41074
rect 17948 40674 18004 40684
rect 18060 40962 18116 40974
rect 18060 40910 18062 40962
rect 18114 40910 18116 40962
rect 17500 39554 17556 39564
rect 16716 38948 16772 38958
rect 16716 38854 16772 38892
rect 16828 38836 16884 38846
rect 16828 38050 16884 38780
rect 17724 38834 17780 38846
rect 17724 38782 17726 38834
rect 17778 38782 17780 38834
rect 17388 38724 17444 38734
rect 17388 38630 17444 38668
rect 16828 37998 16830 38050
rect 16882 37998 16884 38050
rect 16828 37986 16884 37998
rect 17724 37380 17780 38782
rect 17724 37314 17780 37324
rect 17836 38836 17892 38846
rect 17836 37268 17892 38780
rect 18060 38668 18116 40910
rect 19068 40964 19124 40974
rect 19292 40964 19348 41022
rect 19068 40962 19348 40964
rect 19068 40910 19070 40962
rect 19122 40910 19348 40962
rect 19068 40908 19348 40910
rect 18284 40290 18340 40302
rect 18284 40238 18286 40290
rect 18338 40238 18340 40290
rect 18284 38834 18340 40238
rect 19068 39732 19124 40908
rect 19404 40628 19460 41132
rect 18620 39676 19124 39732
rect 19180 40572 19460 40628
rect 19180 39732 19236 40572
rect 19404 40404 19460 40414
rect 19516 40404 19572 41918
rect 20188 41970 20244 42476
rect 20188 41918 20190 41970
rect 20242 41918 20244 41970
rect 19628 41188 19684 41198
rect 19628 41074 19684 41132
rect 19628 41022 19630 41074
rect 19682 41022 19684 41074
rect 19628 41010 19684 41022
rect 19836 40796 20100 40806
rect 19404 40402 19572 40404
rect 19404 40350 19406 40402
rect 19458 40350 19572 40402
rect 19404 40348 19572 40350
rect 19628 40740 19684 40750
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19404 40338 19460 40348
rect 18396 38948 18452 38958
rect 18396 38946 18564 38948
rect 18396 38894 18398 38946
rect 18450 38894 18564 38946
rect 18396 38892 18564 38894
rect 18396 38882 18452 38892
rect 18284 38782 18286 38834
rect 18338 38782 18340 38834
rect 18284 38770 18340 38782
rect 17948 38612 18116 38668
rect 17948 38050 18004 38612
rect 17948 37998 17950 38050
rect 18002 37998 18004 38050
rect 17948 37986 18004 37998
rect 17836 37174 17892 37212
rect 16492 36372 16548 36382
rect 16604 36372 16660 37100
rect 17388 37156 17444 37166
rect 17388 37062 17444 37100
rect 16492 36370 16660 36372
rect 16492 36318 16494 36370
rect 16546 36318 16660 36370
rect 16492 36316 16660 36318
rect 17612 36820 17668 36830
rect 16492 36148 16548 36316
rect 16492 36082 16548 36092
rect 16604 36036 16660 36046
rect 16492 35924 16548 35934
rect 16380 35922 16548 35924
rect 16380 35870 16494 35922
rect 16546 35870 16548 35922
rect 16380 35868 16548 35870
rect 16492 35858 16548 35868
rect 15820 35810 16100 35812
rect 15820 35758 15822 35810
rect 15874 35758 16100 35810
rect 15820 35756 16100 35758
rect 15820 35746 15876 35756
rect 16604 34914 16660 35980
rect 17612 35810 17668 36764
rect 17836 36596 17892 36606
rect 17612 35758 17614 35810
rect 17666 35758 17668 35810
rect 17612 35746 17668 35758
rect 17724 36594 17892 36596
rect 17724 36542 17838 36594
rect 17890 36542 17892 36594
rect 17724 36540 17892 36542
rect 16604 34862 16606 34914
rect 16658 34862 16660 34914
rect 16604 34850 16660 34862
rect 16716 35698 16772 35710
rect 16716 35646 16718 35698
rect 16770 35646 16772 35698
rect 16044 34802 16100 34814
rect 16044 34750 16046 34802
rect 16098 34750 16100 34802
rect 15820 34242 15876 34254
rect 15820 34190 15822 34242
rect 15874 34190 15876 34242
rect 15820 33572 15876 34190
rect 16044 33684 16100 34750
rect 16156 34244 16212 34254
rect 16156 34150 16212 34188
rect 16492 34132 16548 34142
rect 16044 33618 16100 33628
rect 16268 34130 16548 34132
rect 16268 34078 16494 34130
rect 16546 34078 16548 34130
rect 16268 34076 16548 34078
rect 15820 33506 15876 33516
rect 16156 32900 16212 32910
rect 16156 31890 16212 32844
rect 16156 31838 16158 31890
rect 16210 31838 16212 31890
rect 16156 31826 16212 31838
rect 15484 27074 15540 30156
rect 15484 27022 15486 27074
rect 15538 27022 15540 27074
rect 15484 27010 15540 27022
rect 15596 31736 15764 31792
rect 15260 26852 15428 26908
rect 13692 25618 14084 25620
rect 13692 25566 13694 25618
rect 13746 25566 14084 25618
rect 13692 25564 14084 25566
rect 13692 25554 13748 25564
rect 12460 25342 12462 25394
rect 12514 25342 12516 25394
rect 12460 25330 12516 25342
rect 14028 25506 14084 25564
rect 14028 25454 14030 25506
rect 14082 25454 14084 25506
rect 12796 25284 12852 25294
rect 12796 25190 12852 25228
rect 14028 25172 14084 25454
rect 14812 25396 14868 25406
rect 14028 25106 14084 25116
rect 14588 25394 14868 25396
rect 14588 25342 14814 25394
rect 14866 25342 14868 25394
rect 14588 25340 14868 25342
rect 12460 24948 12516 24958
rect 14476 24948 14532 24958
rect 12460 24946 13412 24948
rect 12460 24894 12462 24946
rect 12514 24894 13412 24946
rect 12460 24892 13412 24894
rect 12460 24882 12516 24892
rect 12348 24836 12404 24846
rect 12348 24742 12404 24780
rect 13356 24834 13412 24892
rect 13356 24782 13358 24834
rect 13410 24782 13412 24834
rect 13356 24770 13412 24782
rect 12572 24722 12628 24734
rect 12572 24670 12574 24722
rect 12626 24670 12628 24722
rect 12572 23492 12628 24670
rect 13020 24722 13076 24734
rect 13020 24670 13022 24722
rect 13074 24670 13076 24722
rect 12796 23938 12852 23950
rect 12796 23886 12798 23938
rect 12850 23886 12852 23938
rect 12796 23604 12852 23886
rect 13020 23940 13076 24670
rect 13244 24724 13300 24734
rect 13244 24630 13300 24668
rect 13020 23874 13076 23884
rect 14252 23940 14308 23950
rect 14140 23828 14196 23838
rect 12796 23538 12852 23548
rect 13692 23826 14196 23828
rect 13692 23774 14142 23826
rect 14194 23774 14196 23826
rect 13692 23772 14196 23774
rect 12572 23426 12628 23436
rect 12908 23492 12964 23502
rect 12796 23154 12852 23166
rect 12796 23102 12798 23154
rect 12850 23102 12852 23154
rect 12236 22764 12404 22820
rect 12236 22596 12292 22606
rect 12236 22370 12292 22540
rect 12236 22318 12238 22370
rect 12290 22318 12292 22370
rect 12236 22306 12292 22318
rect 11564 21758 11566 21810
rect 11618 21758 11620 21810
rect 11564 21746 11620 21758
rect 11676 22204 11844 22260
rect 11676 21812 11732 22204
rect 11900 22148 11956 22158
rect 11676 21746 11732 21756
rect 11788 22146 11956 22148
rect 11788 22094 11902 22146
rect 11954 22094 11956 22146
rect 11788 22092 11956 22094
rect 10108 19346 10164 19516
rect 10108 19294 10110 19346
rect 10162 19294 10164 19346
rect 10108 19282 10164 19294
rect 10220 20132 10388 20188
rect 10444 20132 10500 20142
rect 8764 18398 8766 18450
rect 8818 18398 8820 18450
rect 8764 18386 8820 18398
rect 8988 18562 9044 18574
rect 8988 18510 8990 18562
rect 9042 18510 9044 18562
rect 8988 18452 9044 18510
rect 8988 18386 9044 18396
rect 9548 18450 9604 18462
rect 9548 18398 9550 18450
rect 9602 18398 9604 18450
rect 9212 17556 9268 17566
rect 9212 17462 9268 17500
rect 8428 17442 8484 17454
rect 8428 17390 8430 17442
rect 8482 17390 8484 17442
rect 8428 17108 8484 17390
rect 8428 17014 8484 17052
rect 8540 17220 8596 17230
rect 8204 16940 8372 16996
rect 5516 16258 5572 16268
rect 5964 16882 6020 16894
rect 5964 16830 5966 16882
rect 6018 16830 6020 16882
rect 5964 15874 6020 16830
rect 6076 16884 6132 16894
rect 6076 16210 6132 16828
rect 8204 16772 8260 16940
rect 8540 16884 8596 17164
rect 9548 17220 9604 18398
rect 9660 18004 9716 18014
rect 9660 17778 9716 17948
rect 9660 17726 9662 17778
rect 9714 17726 9716 17778
rect 9660 17714 9716 17726
rect 9884 17556 9940 17566
rect 9548 17154 9604 17164
rect 9772 17554 9940 17556
rect 9772 17502 9886 17554
rect 9938 17502 9940 17554
rect 9772 17500 9940 17502
rect 9660 16994 9716 17006
rect 9660 16942 9662 16994
rect 9714 16942 9716 16994
rect 8204 16706 8260 16716
rect 8316 16828 8596 16884
rect 9100 16884 9156 16894
rect 6076 16158 6078 16210
rect 6130 16158 6132 16210
rect 6076 16146 6132 16158
rect 8316 16098 8372 16828
rect 9100 16790 9156 16828
rect 8988 16772 9044 16782
rect 8988 16210 9044 16716
rect 8988 16158 8990 16210
rect 9042 16158 9044 16210
rect 8988 16146 9044 16158
rect 9660 16772 9716 16942
rect 8316 16046 8318 16098
rect 8370 16046 8372 16098
rect 8316 16034 8372 16046
rect 5964 15822 5966 15874
rect 6018 15822 6020 15874
rect 4284 15374 4286 15426
rect 4338 15374 4340 15426
rect 4284 15362 4340 15374
rect 4620 15428 4676 15438
rect 4620 15426 4900 15428
rect 4620 15374 4622 15426
rect 4674 15374 4900 15426
rect 4620 15372 4900 15374
rect 4620 15362 4676 15372
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4844 14532 4900 15372
rect 5068 15316 5124 15326
rect 5068 15222 5124 15260
rect 5516 15316 5572 15326
rect 5964 15316 6020 15822
rect 7980 15540 8036 15550
rect 9100 15540 9156 15550
rect 7980 15538 8372 15540
rect 7980 15486 7982 15538
rect 8034 15486 8372 15538
rect 7980 15484 8372 15486
rect 7980 15474 8036 15484
rect 5516 15314 5684 15316
rect 5516 15262 5518 15314
rect 5570 15262 5684 15314
rect 5516 15260 5684 15262
rect 5516 15250 5572 15260
rect 4844 14438 4900 14476
rect 4620 14308 4676 14318
rect 5628 14308 5684 15260
rect 5964 15250 6020 15260
rect 7308 15204 7364 15214
rect 7308 14642 7364 15148
rect 7308 14590 7310 14642
rect 7362 14590 7364 14642
rect 7308 14578 7364 14590
rect 7980 14532 8036 14542
rect 7980 14438 8036 14476
rect 8316 14418 8372 15484
rect 9100 15446 9156 15484
rect 9548 15314 9604 15326
rect 9548 15262 9550 15314
rect 9602 15262 9604 15314
rect 8540 15204 8596 15214
rect 8540 15110 8596 15148
rect 9548 14532 9604 15262
rect 9660 15204 9716 16716
rect 9660 15138 9716 15148
rect 9772 14642 9828 17500
rect 9884 17490 9940 17500
rect 10220 17554 10276 20132
rect 10444 20018 10500 20076
rect 10668 20130 10724 20142
rect 10668 20078 10670 20130
rect 10722 20078 10724 20130
rect 10444 19966 10446 20018
rect 10498 19966 10500 20018
rect 10444 19954 10500 19966
rect 10556 20020 10612 20030
rect 10556 19458 10612 19964
rect 10556 19406 10558 19458
rect 10610 19406 10612 19458
rect 10556 19394 10612 19406
rect 10668 19460 10724 20078
rect 11004 20132 11172 20188
rect 11228 21698 11284 21710
rect 11228 21646 11230 21698
rect 11282 21646 11284 21698
rect 11228 20188 11284 21646
rect 11788 21588 11844 22092
rect 11900 22082 11956 22092
rect 12236 21812 12292 21822
rect 12348 21812 12404 22764
rect 12796 22260 12852 23102
rect 12796 22194 12852 22204
rect 11900 21810 12404 21812
rect 11900 21758 12238 21810
rect 12290 21758 12404 21810
rect 11900 21756 12404 21758
rect 12460 22148 12516 22158
rect 11900 21698 11956 21756
rect 12236 21746 12292 21756
rect 12460 21700 12516 22092
rect 11900 21646 11902 21698
rect 11954 21646 11956 21698
rect 11900 21634 11956 21646
rect 12348 21644 12516 21700
rect 11340 20916 11396 20926
rect 11340 20822 11396 20860
rect 11228 20132 11508 20188
rect 10780 19572 10836 19582
rect 10836 19516 10948 19572
rect 10780 19506 10836 19516
rect 10668 19394 10724 19404
rect 10892 19458 10948 19516
rect 10892 19406 10894 19458
rect 10946 19406 10948 19458
rect 10892 19394 10948 19406
rect 10332 18452 10388 18462
rect 10332 18358 10388 18396
rect 10220 17502 10222 17554
rect 10274 17502 10276 17554
rect 9996 16994 10052 17006
rect 9996 16942 9998 16994
rect 10050 16942 10052 16994
rect 9996 16660 10052 16942
rect 9996 16594 10052 16604
rect 10220 15540 10276 17502
rect 10444 18004 10500 18014
rect 10444 16882 10500 17948
rect 10668 17892 10724 17902
rect 10668 17798 10724 17836
rect 11004 17892 11060 20132
rect 11452 20020 11508 20132
rect 11676 20132 11732 20142
rect 11676 20038 11732 20076
rect 11452 19926 11508 19964
rect 11116 19796 11172 19806
rect 11116 19702 11172 19740
rect 11340 19796 11396 19806
rect 11340 19234 11396 19740
rect 11340 19182 11342 19234
rect 11394 19182 11396 19234
rect 11004 17890 11172 17892
rect 11004 17838 11006 17890
rect 11058 17838 11172 17890
rect 11004 17836 11172 17838
rect 11004 17826 11060 17836
rect 10444 16830 10446 16882
rect 10498 16830 10500 16882
rect 10444 16818 10500 16830
rect 10668 16994 10724 17006
rect 10668 16942 10670 16994
rect 10722 16942 10724 16994
rect 10668 16884 10724 16942
rect 11116 16884 11172 17836
rect 11340 17554 11396 19182
rect 11788 19572 11844 21532
rect 12348 21028 12404 21644
rect 12572 21588 12628 21598
rect 12012 20972 12404 21028
rect 12460 21586 12628 21588
rect 12460 21534 12574 21586
rect 12626 21534 12628 21586
rect 12460 21532 12628 21534
rect 12012 20690 12068 20972
rect 12012 20638 12014 20690
rect 12066 20638 12068 20690
rect 12012 20130 12068 20638
rect 12124 20802 12180 20814
rect 12124 20750 12126 20802
rect 12178 20750 12180 20802
rect 12124 20188 12180 20750
rect 12124 20132 12292 20188
rect 12012 20078 12014 20130
rect 12066 20078 12068 20130
rect 12012 19908 12068 20078
rect 12012 19842 12068 19852
rect 12236 19908 12292 20132
rect 12236 19842 12292 19852
rect 12348 20020 12404 20030
rect 11676 19122 11732 19134
rect 11676 19070 11678 19122
rect 11730 19070 11732 19122
rect 11564 18004 11620 18014
rect 11340 17502 11342 17554
rect 11394 17502 11396 17554
rect 11340 17490 11396 17502
rect 11452 17948 11564 18004
rect 11452 16996 11508 17948
rect 11564 17938 11620 17948
rect 11676 17668 11732 19070
rect 11564 17554 11620 17566
rect 11564 17502 11566 17554
rect 11618 17502 11620 17554
rect 11564 17444 11620 17502
rect 11564 17378 11620 17388
rect 11676 17332 11732 17612
rect 11676 17266 11732 17276
rect 11452 16940 11620 16996
rect 11116 16828 11284 16884
rect 10668 16818 10724 16828
rect 11116 16660 11172 16670
rect 10220 15474 10276 15484
rect 10332 16658 11172 16660
rect 10332 16606 11118 16658
rect 11170 16606 11172 16658
rect 10332 16604 11172 16606
rect 9884 15426 9940 15438
rect 9884 15374 9886 15426
rect 9938 15374 9940 15426
rect 9884 14756 9940 15374
rect 10332 15314 10388 16604
rect 11116 16594 11172 16604
rect 11116 16212 11172 16222
rect 11228 16212 11284 16828
rect 11452 16772 11508 16782
rect 11452 16678 11508 16716
rect 11116 16210 11284 16212
rect 11116 16158 11118 16210
rect 11170 16158 11284 16210
rect 11116 16156 11284 16158
rect 11116 16146 11172 16156
rect 11564 16100 11620 16940
rect 11564 16044 11732 16100
rect 11564 15876 11620 15886
rect 11228 15874 11620 15876
rect 11228 15822 11566 15874
rect 11618 15822 11620 15874
rect 11228 15820 11620 15822
rect 10332 15262 10334 15314
rect 10386 15262 10388 15314
rect 10332 15250 10388 15262
rect 10556 15426 10612 15438
rect 10556 15374 10558 15426
rect 10610 15374 10612 15426
rect 9884 14690 9940 14700
rect 9772 14590 9774 14642
rect 9826 14590 9828 14642
rect 9772 14578 9828 14590
rect 10556 14644 10612 15374
rect 10892 15428 10948 15438
rect 10892 15426 11172 15428
rect 10892 15374 10894 15426
rect 10946 15374 11172 15426
rect 10892 15372 11172 15374
rect 10892 15362 10948 15372
rect 10556 14578 10612 14588
rect 9548 14466 9604 14476
rect 8316 14366 8318 14418
rect 8370 14366 8372 14418
rect 4620 14306 4900 14308
rect 4620 14254 4622 14306
rect 4674 14254 4900 14306
rect 4620 14252 4900 14254
rect 4620 14242 4676 14252
rect 4508 13972 4564 13982
rect 4172 13970 4564 13972
rect 4172 13918 4510 13970
rect 4562 13918 4564 13970
rect 4172 13916 4564 13918
rect 3724 13906 3780 13916
rect 4508 13906 4564 13916
rect 2044 13468 2212 13524
rect 1820 12740 1876 12750
rect 1820 12180 1876 12684
rect 1820 12178 2100 12180
rect 1820 12126 1822 12178
rect 1874 12126 2100 12178
rect 1820 12124 2100 12126
rect 1820 12114 1876 12124
rect 1820 11508 1876 11518
rect 1820 10610 1876 11452
rect 1820 10558 1822 10610
rect 1874 10558 1876 10610
rect 1820 10546 1876 10558
rect 2044 10612 2100 12124
rect 2156 12178 2212 13468
rect 3612 13458 3668 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 3612 12850 3668 12862
rect 3612 12798 3614 12850
rect 3666 12798 3668 12850
rect 3500 12740 3556 12750
rect 3500 12646 3556 12684
rect 2156 12126 2158 12178
rect 2210 12126 2212 12178
rect 2156 12114 2212 12126
rect 3612 11620 3668 12798
rect 4732 12404 4788 12414
rect 4844 12404 4900 14252
rect 5292 13972 5348 13982
rect 5292 13878 5348 13916
rect 5628 13746 5684 14252
rect 7196 14308 7252 14318
rect 7196 14214 7252 14252
rect 8316 13970 8372 14366
rect 8316 13918 8318 13970
rect 8370 13918 8372 13970
rect 5628 13694 5630 13746
rect 5682 13694 5684 13746
rect 5628 13682 5684 13694
rect 6076 13746 6132 13758
rect 6076 13694 6078 13746
rect 6130 13694 6132 13746
rect 5068 13524 5124 13534
rect 5124 13468 5236 13524
rect 5068 13458 5124 13468
rect 4732 12402 4900 12404
rect 4732 12350 4734 12402
rect 4786 12350 4900 12402
rect 4732 12348 4900 12350
rect 5180 12404 5236 13468
rect 6076 12740 6132 13694
rect 8316 13748 8372 13918
rect 11116 13858 11172 15372
rect 11228 15426 11284 15820
rect 11564 15810 11620 15820
rect 11564 15540 11620 15550
rect 11676 15540 11732 16044
rect 11788 15764 11844 19516
rect 12348 19460 12404 19964
rect 12236 19404 12404 19460
rect 12236 17780 12292 19404
rect 12348 19234 12404 19246
rect 12348 19182 12350 19234
rect 12402 19182 12404 19234
rect 12348 18900 12404 19182
rect 12348 18834 12404 18844
rect 12460 18338 12516 21532
rect 12572 21522 12628 21532
rect 12908 20690 12964 23436
rect 13692 22482 13748 23772
rect 14140 23762 14196 23772
rect 14252 23380 14308 23884
rect 14476 23938 14532 24892
rect 14588 24050 14644 25340
rect 14812 25330 14868 25340
rect 14588 23998 14590 24050
rect 14642 23998 14644 24050
rect 14588 23986 14644 23998
rect 15148 24724 15204 24734
rect 14476 23886 14478 23938
rect 14530 23886 14532 23938
rect 14476 23874 14532 23886
rect 14700 23940 14756 23950
rect 14700 23846 14756 23884
rect 14364 23492 14420 23502
rect 14924 23492 14980 23502
rect 14420 23436 14924 23492
rect 14364 23426 14420 23436
rect 13692 22430 13694 22482
rect 13746 22430 13748 22482
rect 13692 22418 13748 22430
rect 13804 23324 14308 23380
rect 14924 23378 14980 23436
rect 14924 23326 14926 23378
rect 14978 23326 14980 23378
rect 13804 22594 13860 23324
rect 14924 23314 14980 23326
rect 14476 23268 14532 23278
rect 14140 23212 14476 23268
rect 13804 22542 13806 22594
rect 13858 22542 13860 22594
rect 13020 22146 13076 22158
rect 13020 22094 13022 22146
rect 13074 22094 13076 22146
rect 13020 21924 13076 22094
rect 13580 22148 13636 22158
rect 13804 22148 13860 22542
rect 13580 22054 13636 22092
rect 13692 22092 13860 22148
rect 13916 23156 13972 23166
rect 13020 21858 13076 21868
rect 13132 21700 13188 21710
rect 13132 21606 13188 21644
rect 13468 21698 13524 21710
rect 13468 21646 13470 21698
rect 13522 21646 13524 21698
rect 13468 20916 13524 21646
rect 13692 21588 13748 22092
rect 13804 21924 13860 21934
rect 13804 21810 13860 21868
rect 13804 21758 13806 21810
rect 13858 21758 13860 21810
rect 13804 21746 13860 21758
rect 13692 21532 13860 21588
rect 13580 21028 13636 21038
rect 13580 20934 13636 20972
rect 13468 20850 13524 20860
rect 12908 20638 12910 20690
rect 12962 20638 12964 20690
rect 12908 20626 12964 20638
rect 13468 20690 13524 20702
rect 13468 20638 13470 20690
rect 13522 20638 13524 20690
rect 12460 18286 12462 18338
rect 12514 18286 12516 18338
rect 12460 18274 12516 18286
rect 12572 20578 12628 20590
rect 12572 20526 12574 20578
rect 12626 20526 12628 20578
rect 12572 20132 12628 20526
rect 13468 20188 13524 20638
rect 13468 20132 13748 20188
rect 12236 17724 12404 17780
rect 12124 17668 12180 17678
rect 12124 16996 12180 17612
rect 12124 16902 12180 16940
rect 12236 17556 12292 17566
rect 12236 16884 12292 17500
rect 12348 16996 12404 17724
rect 12460 17668 12516 17678
rect 12572 17668 12628 20076
rect 12796 20020 12852 20030
rect 12796 19926 12852 19964
rect 13468 20018 13524 20030
rect 13468 19966 13470 20018
rect 13522 19966 13524 20018
rect 13468 19684 13524 19966
rect 13692 20020 13748 20132
rect 13580 19908 13636 19918
rect 13580 19814 13636 19852
rect 13580 19684 13636 19694
rect 13468 19628 13580 19684
rect 12796 19460 12852 19470
rect 12684 19236 12740 19246
rect 12684 18452 12740 19180
rect 12796 18676 12852 19404
rect 13468 19460 13524 19470
rect 13468 19234 13524 19404
rect 13468 19182 13470 19234
rect 13522 19182 13524 19234
rect 13356 19124 13412 19134
rect 12796 18582 12852 18620
rect 12908 19010 12964 19022
rect 12908 18958 12910 19010
rect 12962 18958 12964 19010
rect 12908 18564 12964 18958
rect 13020 18788 13076 18798
rect 13356 18788 13412 19068
rect 13020 18674 13076 18732
rect 13020 18622 13022 18674
rect 13074 18622 13076 18674
rect 13020 18610 13076 18622
rect 13132 18732 13412 18788
rect 12908 18498 12964 18508
rect 13132 18452 13188 18732
rect 13468 18564 13524 19182
rect 13580 19012 13636 19628
rect 13692 19348 13748 19964
rect 13692 19282 13748 19292
rect 13804 19908 13860 21532
rect 13916 20914 13972 23100
rect 14140 23154 14196 23212
rect 14476 23202 14532 23212
rect 15036 23268 15092 23278
rect 14140 23102 14142 23154
rect 14194 23102 14196 23154
rect 14140 23090 14196 23102
rect 14812 23154 14868 23166
rect 14812 23102 14814 23154
rect 14866 23102 14868 23154
rect 14476 23044 14532 23054
rect 14812 23044 14868 23102
rect 14476 23042 14868 23044
rect 14476 22990 14478 23042
rect 14530 22990 14868 23042
rect 14476 22988 14868 22990
rect 13916 20862 13918 20914
rect 13970 20862 13972 20914
rect 13916 20850 13972 20862
rect 14028 21700 14084 21710
rect 14028 20692 14084 21644
rect 14364 21476 14420 21486
rect 14476 21476 14532 22988
rect 14924 22930 14980 22942
rect 14924 22878 14926 22930
rect 14978 22878 14980 22930
rect 14588 22482 14644 22494
rect 14588 22430 14590 22482
rect 14642 22430 14644 22482
rect 14588 21924 14644 22430
rect 14700 21924 14756 21934
rect 14588 21868 14700 21924
rect 14420 21420 14532 21476
rect 14364 21382 14420 21420
rect 13804 19236 13860 19852
rect 13804 19170 13860 19180
rect 13916 20636 14084 20692
rect 14140 20804 14196 20814
rect 13580 18946 13636 18956
rect 13804 19012 13860 19022
rect 13804 18918 13860 18956
rect 13468 18508 13860 18564
rect 12684 18396 12852 18452
rect 12460 17666 12740 17668
rect 12460 17614 12462 17666
rect 12514 17614 12740 17666
rect 12460 17612 12740 17614
rect 12460 17602 12516 17612
rect 12684 17106 12740 17612
rect 12684 17054 12686 17106
rect 12738 17054 12740 17106
rect 12684 17042 12740 17054
rect 12348 16940 12628 16996
rect 12236 16882 12404 16884
rect 12236 16830 12238 16882
rect 12290 16830 12404 16882
rect 12236 16828 12404 16830
rect 12236 16818 12292 16828
rect 12236 16548 12292 16558
rect 11900 16212 11956 16222
rect 12236 16212 12292 16492
rect 11900 16210 12292 16212
rect 11900 16158 11902 16210
rect 11954 16158 12292 16210
rect 11900 16156 12292 16158
rect 11900 16146 11956 16156
rect 11788 15708 11956 15764
rect 11564 15538 11732 15540
rect 11564 15486 11566 15538
rect 11618 15486 11732 15538
rect 11564 15484 11732 15486
rect 11788 15540 11844 15550
rect 11564 15474 11620 15484
rect 11228 15374 11230 15426
rect 11282 15374 11284 15426
rect 11228 15362 11284 15374
rect 11788 15314 11844 15484
rect 11788 15262 11790 15314
rect 11842 15262 11844 15314
rect 11788 15250 11844 15262
rect 11900 15092 11956 15708
rect 12236 15538 12292 16156
rect 12348 16098 12404 16828
rect 12572 16660 12628 16940
rect 12572 16594 12628 16604
rect 12684 16884 12740 16894
rect 12348 16046 12350 16098
rect 12402 16046 12404 16098
rect 12348 16034 12404 16046
rect 12684 15988 12740 16828
rect 12684 15894 12740 15932
rect 12236 15486 12238 15538
rect 12290 15486 12292 15538
rect 12236 15474 12292 15486
rect 12572 15316 12628 15326
rect 12628 15260 12740 15316
rect 12572 15222 12628 15260
rect 11116 13806 11118 13858
rect 11170 13806 11172 13858
rect 11116 13794 11172 13806
rect 11788 15036 11956 15092
rect 8316 13682 8372 13692
rect 10332 13748 10388 13758
rect 10332 13654 10388 13692
rect 9100 13524 9156 13534
rect 8652 13522 9156 13524
rect 8652 13470 9102 13522
rect 9154 13470 9156 13522
rect 8652 13468 9156 13470
rect 8652 13074 8708 13468
rect 9100 13458 9156 13468
rect 8652 13022 8654 13074
rect 8706 13022 8708 13074
rect 8652 13010 8708 13022
rect 6076 12674 6132 12684
rect 7308 12740 7364 12750
rect 5292 12404 5348 12414
rect 5180 12402 5348 12404
rect 5180 12350 5294 12402
rect 5346 12350 5348 12402
rect 5180 12348 5348 12350
rect 4732 12338 4788 12348
rect 4060 12180 4116 12190
rect 3612 11554 3668 11564
rect 3724 11956 3780 11966
rect 3500 11508 3556 11518
rect 3500 11396 3556 11452
rect 3724 11506 3780 11900
rect 3724 11454 3726 11506
rect 3778 11454 3780 11506
rect 3724 11442 3780 11454
rect 4060 11618 4116 12124
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4060 11566 4062 11618
rect 4114 11566 4116 11618
rect 3612 11396 3668 11406
rect 3500 11394 3668 11396
rect 3500 11342 3614 11394
rect 3666 11342 3668 11394
rect 3500 11340 3668 11342
rect 3612 11330 3668 11340
rect 2156 10612 2212 10622
rect 2044 10610 2212 10612
rect 2044 10558 2158 10610
rect 2210 10558 2212 10610
rect 2044 10556 2212 10558
rect 2156 10546 2212 10556
rect 3724 10388 3780 10398
rect 2492 10052 2548 10062
rect 2044 9604 2100 9614
rect 1932 9044 1988 9054
rect 1932 5908 1988 8988
rect 2044 7474 2100 9548
rect 2044 7422 2046 7474
rect 2098 7422 2100 7474
rect 2044 7252 2100 7422
rect 2492 7474 2548 9996
rect 2940 9716 2996 9726
rect 2940 9266 2996 9660
rect 2940 9214 2942 9266
rect 2994 9214 2996 9266
rect 2940 9202 2996 9214
rect 3724 9266 3780 10332
rect 4060 10052 4116 11566
rect 4844 11396 4900 12348
rect 5292 12338 5348 12348
rect 6188 12290 6244 12302
rect 6188 12238 6190 12290
rect 6242 12238 6244 12290
rect 5404 11956 5460 11966
rect 5404 11862 5460 11900
rect 4060 9986 4116 9996
rect 4172 11282 4228 11294
rect 4172 11230 4174 11282
rect 4226 11230 4228 11282
rect 4172 9828 4228 11230
rect 4732 10836 4788 10846
rect 4844 10836 4900 11340
rect 4732 10834 4900 10836
rect 4732 10782 4734 10834
rect 4786 10782 4900 10834
rect 4732 10780 4900 10782
rect 5292 11620 5348 11630
rect 5292 10834 5348 11564
rect 6188 11506 6244 12238
rect 6188 11454 6190 11506
rect 6242 11454 6244 11506
rect 5628 11396 5684 11406
rect 5628 11302 5684 11340
rect 6076 11396 6132 11406
rect 5292 10782 5294 10834
rect 5346 10782 5348 10834
rect 4732 10770 4788 10780
rect 5292 10770 5348 10782
rect 6076 10834 6132 11340
rect 6076 10782 6078 10834
rect 6130 10782 6132 10834
rect 6076 10770 6132 10782
rect 6076 10612 6132 10622
rect 5180 10388 5236 10398
rect 5068 10332 5180 10388
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4172 9762 4228 9772
rect 4284 9714 4340 9726
rect 4284 9662 4286 9714
rect 4338 9662 4340 9714
rect 4172 9604 4228 9614
rect 4172 9510 4228 9548
rect 3724 9214 3726 9266
rect 3778 9214 3780 9266
rect 3724 9202 3780 9214
rect 2492 7422 2494 7474
rect 2546 7422 2548 7474
rect 2492 7410 2548 7422
rect 2044 7196 2324 7252
rect 2156 5908 2212 5918
rect 1932 5906 2212 5908
rect 1932 5854 2158 5906
rect 2210 5854 2212 5906
rect 1932 5852 2212 5854
rect 2268 5908 2324 7196
rect 4284 6916 4340 9662
rect 4956 9716 5012 9726
rect 4956 9622 5012 9660
rect 4844 9602 4900 9614
rect 4844 9550 4846 9602
rect 4898 9550 4900 9602
rect 4844 9044 4900 9550
rect 5068 9492 5124 10332
rect 5180 10322 5236 10332
rect 5404 10388 5460 10398
rect 5404 10386 6020 10388
rect 5404 10334 5406 10386
rect 5458 10334 6020 10386
rect 5404 10332 6020 10334
rect 5404 10322 5460 10332
rect 5964 9938 6020 10332
rect 6076 10050 6132 10556
rect 6188 10388 6244 11454
rect 7308 11394 7364 12684
rect 8540 12740 8596 12750
rect 8540 12646 8596 12684
rect 11788 12404 11844 15036
rect 12572 14756 12628 14766
rect 11900 14644 11956 14654
rect 11900 14550 11956 14588
rect 12572 14532 12628 14700
rect 12460 14530 12628 14532
rect 12460 14478 12574 14530
rect 12626 14478 12628 14530
rect 12460 14476 12628 14478
rect 12012 12404 12068 12414
rect 11788 12402 12068 12404
rect 11788 12350 11790 12402
rect 11842 12350 12014 12402
rect 12066 12350 12068 12402
rect 11788 12348 12068 12350
rect 11788 12338 11844 12348
rect 12012 12338 12068 12348
rect 11564 12292 11620 12302
rect 8428 12178 8484 12190
rect 8428 12126 8430 12178
rect 8482 12126 8484 12178
rect 7308 11342 7310 11394
rect 7362 11342 7364 11394
rect 7308 11330 7364 11342
rect 7980 11956 8036 11966
rect 7980 11394 8036 11900
rect 8428 11508 8484 12126
rect 8876 12180 8932 12190
rect 8876 12086 8932 12124
rect 9660 12066 9716 12078
rect 9660 12014 9662 12066
rect 9714 12014 9716 12066
rect 9548 11956 9604 11966
rect 9548 11862 9604 11900
rect 9660 11620 9716 12014
rect 10108 12068 10164 12078
rect 10108 12066 11508 12068
rect 10108 12014 10110 12066
rect 10162 12014 11508 12066
rect 10108 12012 11508 12014
rect 10108 12002 10164 12012
rect 9996 11956 10052 11966
rect 9660 11554 9716 11564
rect 9772 11954 10052 11956
rect 9772 11902 9998 11954
rect 10050 11902 10052 11954
rect 9772 11900 10052 11902
rect 8428 11442 8484 11452
rect 7980 11342 7982 11394
rect 8034 11342 8036 11394
rect 6188 10322 6244 10332
rect 6636 10612 6692 10622
rect 6076 9998 6078 10050
rect 6130 9998 6132 10050
rect 6076 9986 6132 9998
rect 5964 9886 5966 9938
rect 6018 9886 6020 9938
rect 5964 9874 6020 9886
rect 4844 8978 4900 8988
rect 4956 9436 5124 9492
rect 5516 9828 5572 9838
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4956 7698 5012 9436
rect 4956 7646 4958 7698
rect 5010 7646 5012 7698
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4284 6850 4340 6860
rect 4956 6132 5012 7646
rect 5516 7698 5572 9772
rect 5964 9044 6020 9054
rect 5964 8950 6020 8988
rect 6636 9042 6692 10556
rect 7980 9826 8036 11342
rect 8428 10612 8484 10622
rect 8428 10518 8484 10556
rect 9100 10612 9156 10622
rect 9660 10612 9716 10622
rect 9772 10612 9828 11900
rect 9996 11890 10052 11900
rect 11340 11732 11396 11742
rect 11004 11620 11060 11630
rect 11004 11526 11060 11564
rect 11340 11394 11396 11676
rect 11340 11342 11342 11394
rect 11394 11342 11396 11394
rect 11340 11330 11396 11342
rect 10332 11172 10388 11182
rect 10332 11078 10388 11116
rect 10668 11172 10724 11182
rect 9100 10518 9156 10556
rect 9212 10610 9828 10612
rect 9212 10558 9662 10610
rect 9714 10558 9828 10610
rect 9212 10556 9828 10558
rect 9996 10612 10052 10622
rect 7980 9774 7982 9826
rect 8034 9774 8036 9826
rect 7980 9762 8036 9774
rect 8428 9828 8484 9838
rect 9212 9828 9268 10556
rect 9660 10546 9716 10556
rect 9884 10388 9940 10398
rect 8428 9826 9268 9828
rect 8428 9774 8430 9826
rect 8482 9774 9268 9826
rect 8428 9772 9268 9774
rect 9772 10332 9884 10388
rect 8428 9762 8484 9772
rect 6636 8990 6638 9042
rect 6690 8990 6692 9042
rect 6636 8978 6692 8990
rect 9772 9044 9828 10332
rect 9884 10322 9940 10332
rect 9884 9268 9940 9278
rect 9996 9268 10052 10556
rect 10668 9714 10724 11116
rect 11452 10050 11508 12012
rect 11564 11282 11620 12236
rect 12348 12290 12404 12302
rect 12348 12238 12350 12290
rect 12402 12238 12404 12290
rect 12348 12180 12404 12238
rect 12348 11732 12404 12124
rect 12348 11666 12404 11676
rect 12012 11396 12068 11406
rect 12012 11302 12068 11340
rect 11564 11230 11566 11282
rect 11618 11230 11620 11282
rect 11564 11218 11620 11230
rect 12236 11170 12292 11182
rect 12236 11118 12238 11170
rect 12290 11118 12292 11170
rect 12236 10836 12292 11118
rect 12236 10770 12292 10780
rect 12460 11172 12516 14476
rect 12572 14466 12628 14476
rect 12460 10834 12516 11116
rect 12460 10782 12462 10834
rect 12514 10782 12516 10834
rect 12460 10770 12516 10782
rect 12572 12738 12628 12750
rect 12572 12686 12574 12738
rect 12626 12686 12628 12738
rect 11452 9998 11454 10050
rect 11506 9998 11508 10050
rect 11452 9986 11508 9998
rect 10668 9662 10670 9714
rect 10722 9662 10724 9714
rect 10668 9650 10724 9662
rect 12572 9716 12628 12686
rect 12684 12402 12740 15260
rect 12796 15092 12852 18396
rect 13020 18396 13188 18452
rect 13244 18452 13300 18462
rect 12908 18340 12964 18350
rect 12908 18246 12964 18284
rect 12908 17666 12964 17678
rect 12908 17614 12910 17666
rect 12962 17614 12964 17666
rect 12908 17556 12964 17614
rect 12908 17490 12964 17500
rect 13020 17106 13076 18396
rect 13244 17332 13300 18396
rect 13356 18450 13412 18462
rect 13356 18398 13358 18450
rect 13410 18398 13412 18450
rect 13356 17666 13412 18398
rect 13356 17614 13358 17666
rect 13410 17614 13412 17666
rect 13356 17602 13412 17614
rect 13692 17668 13748 17678
rect 13692 17574 13748 17612
rect 13580 17556 13636 17566
rect 13580 17462 13636 17500
rect 13244 17276 13636 17332
rect 13020 17054 13022 17106
rect 13074 17054 13076 17106
rect 13020 17042 13076 17054
rect 13132 17108 13188 17118
rect 12908 16996 12964 17006
rect 12908 15314 12964 16940
rect 13132 15538 13188 17052
rect 13580 16770 13636 17276
rect 13580 16718 13582 16770
rect 13634 16718 13636 16770
rect 13580 16706 13636 16718
rect 13804 16098 13860 18508
rect 13916 17668 13972 20636
rect 14028 20130 14084 20142
rect 14028 20078 14030 20130
rect 14082 20078 14084 20130
rect 14028 19234 14084 20078
rect 14028 19182 14030 19234
rect 14082 19182 14084 19234
rect 14028 19124 14084 19182
rect 14028 19058 14084 19068
rect 14028 18676 14084 18686
rect 14140 18676 14196 20748
rect 14700 20188 14756 21868
rect 14924 21812 14980 22878
rect 15036 22370 15092 23212
rect 15036 22318 15038 22370
rect 15090 22318 15092 22370
rect 15036 22306 15092 22318
rect 14924 21746 14980 21756
rect 15036 21924 15092 21934
rect 15036 21810 15092 21868
rect 15036 21758 15038 21810
rect 15090 21758 15092 21810
rect 15036 21746 15092 21758
rect 15148 21810 15204 24668
rect 15148 21758 15150 21810
rect 15202 21758 15204 21810
rect 15148 21746 15204 21758
rect 14812 21586 14868 21598
rect 14812 21534 14814 21586
rect 14866 21534 14868 21586
rect 14812 20804 14868 21534
rect 14812 20738 14868 20748
rect 14924 21586 14980 21598
rect 14924 21534 14926 21586
rect 14978 21534 14980 21586
rect 14924 21028 14980 21534
rect 15260 21028 15316 26852
rect 15372 25172 15428 25182
rect 15372 24050 15428 25116
rect 15372 23998 15374 24050
rect 15426 23998 15428 24050
rect 15372 23940 15428 23998
rect 15372 23874 15428 23884
rect 15596 23548 15652 31736
rect 15708 31668 15764 31678
rect 15708 31666 15988 31668
rect 15708 31614 15710 31666
rect 15762 31614 15988 31666
rect 15708 31612 15988 31614
rect 15708 31602 15764 31612
rect 15708 31108 15764 31118
rect 15708 31014 15764 31052
rect 15820 30100 15876 30110
rect 15820 28532 15876 30044
rect 15932 29540 15988 31612
rect 16044 30996 16100 31006
rect 16044 30902 16100 30940
rect 16268 30548 16324 34076
rect 16492 34066 16548 34076
rect 16716 33572 16772 35646
rect 17500 35698 17556 35710
rect 17500 35646 17502 35698
rect 17554 35646 17556 35698
rect 16828 34244 16884 34254
rect 16884 34188 17108 34244
rect 16828 34150 16884 34188
rect 16940 33572 16996 33582
rect 16716 33516 16940 33572
rect 16940 33346 16996 33516
rect 16940 33294 16942 33346
rect 16994 33294 16996 33346
rect 16604 32340 16660 32350
rect 16940 32340 16996 33294
rect 16604 32338 16772 32340
rect 16604 32286 16606 32338
rect 16658 32286 16772 32338
rect 16604 32284 16772 32286
rect 16604 32274 16660 32284
rect 16604 31892 16660 31902
rect 16604 31778 16660 31836
rect 16604 31726 16606 31778
rect 16658 31726 16660 31778
rect 16604 31714 16660 31726
rect 16716 31780 16772 32284
rect 16940 32274 16996 32284
rect 16940 31780 16996 31790
rect 16716 31778 16996 31780
rect 16716 31726 16942 31778
rect 16994 31726 16996 31778
rect 16716 31724 16996 31726
rect 16940 31714 16996 31724
rect 16380 31106 16436 31118
rect 16380 31054 16382 31106
rect 16434 31054 16436 31106
rect 16380 30884 16436 31054
rect 16380 30818 16436 30828
rect 16828 31108 16884 31118
rect 16828 30884 16884 31052
rect 16828 30882 16996 30884
rect 16828 30830 16830 30882
rect 16882 30830 16996 30882
rect 16828 30828 16996 30830
rect 16828 30818 16884 30828
rect 16268 30492 16436 30548
rect 15932 29474 15988 29484
rect 15820 27970 15876 28476
rect 15820 27918 15822 27970
rect 15874 27918 15876 27970
rect 15820 27906 15876 27918
rect 16268 26964 16324 26974
rect 16268 26850 16324 26908
rect 16268 26798 16270 26850
rect 16322 26798 16324 26850
rect 16268 26786 16324 26798
rect 15708 23940 15764 23978
rect 15764 23884 15876 23940
rect 15708 23874 15764 23884
rect 15372 23492 15428 23502
rect 15372 22370 15428 23436
rect 15372 22318 15374 22370
rect 15426 22318 15428 22370
rect 15372 22036 15428 22318
rect 15372 21970 15428 21980
rect 15484 23492 15652 23548
rect 15708 23716 15764 23726
rect 15708 23492 15764 23660
rect 14924 20692 14980 20972
rect 14924 20626 14980 20636
rect 15148 20972 15316 21028
rect 15372 21586 15428 21598
rect 15372 21534 15374 21586
rect 15426 21534 15428 21586
rect 14700 20132 14980 20188
rect 14084 18620 14196 18676
rect 14252 19796 14308 19806
rect 14252 18674 14308 19740
rect 14476 19460 14532 19470
rect 14476 19346 14532 19404
rect 14476 19294 14478 19346
rect 14530 19294 14532 19346
rect 14476 19282 14532 19294
rect 14252 18622 14254 18674
rect 14306 18622 14308 18674
rect 14028 18582 14084 18620
rect 14252 18610 14308 18622
rect 14700 18452 14756 18462
rect 14700 18358 14756 18396
rect 14140 18338 14196 18350
rect 14140 18286 14142 18338
rect 14194 18286 14196 18338
rect 14140 17892 14196 18286
rect 14140 17836 14868 17892
rect 14812 17778 14868 17836
rect 14812 17726 14814 17778
rect 14866 17726 14868 17778
rect 14812 17714 14868 17726
rect 14028 17668 14084 17678
rect 13916 17666 14084 17668
rect 13916 17614 14030 17666
rect 14082 17614 14084 17666
rect 13916 17612 14084 17614
rect 14028 17602 14084 17612
rect 13804 16046 13806 16098
rect 13858 16046 13860 16098
rect 13804 16034 13860 16046
rect 13916 16884 13972 16894
rect 13580 15988 13636 15998
rect 13580 15894 13636 15932
rect 13132 15486 13134 15538
rect 13186 15486 13188 15538
rect 13132 15474 13188 15486
rect 12908 15262 12910 15314
rect 12962 15262 12964 15314
rect 12908 15250 12964 15262
rect 13244 15204 13300 15214
rect 13020 15202 13300 15204
rect 13020 15150 13246 15202
rect 13298 15150 13300 15202
rect 13020 15148 13300 15150
rect 13020 15092 13076 15148
rect 13244 15138 13300 15148
rect 12796 15036 13076 15092
rect 13916 14530 13972 16828
rect 14364 16324 14420 16334
rect 14364 16230 14420 16268
rect 14700 15876 14756 15886
rect 14140 15874 14756 15876
rect 14140 15822 14702 15874
rect 14754 15822 14756 15874
rect 14140 15820 14756 15822
rect 14028 15316 14084 15326
rect 14140 15316 14196 15820
rect 14700 15810 14756 15820
rect 14252 15428 14308 15438
rect 14252 15426 14756 15428
rect 14252 15374 14254 15426
rect 14306 15374 14756 15426
rect 14252 15372 14756 15374
rect 14252 15362 14308 15372
rect 14028 15314 14196 15316
rect 14028 15262 14030 15314
rect 14082 15262 14196 15314
rect 14028 15260 14196 15262
rect 14028 15250 14084 15260
rect 13916 14478 13918 14530
rect 13970 14478 13972 14530
rect 13916 14466 13972 14478
rect 14588 15204 14644 15214
rect 14140 13860 14196 13870
rect 13804 13858 14196 13860
rect 13804 13806 14142 13858
rect 14194 13806 14196 13858
rect 13804 13804 14196 13806
rect 13244 13748 13300 13758
rect 13244 13634 13300 13692
rect 13244 13582 13246 13634
rect 13298 13582 13300 13634
rect 13244 13570 13300 13582
rect 13020 13300 13076 13310
rect 12908 12852 12964 12862
rect 12908 12758 12964 12796
rect 12684 12350 12686 12402
rect 12738 12350 12740 12402
rect 12684 11394 12740 12350
rect 13020 12290 13076 13244
rect 13692 12964 13748 12974
rect 13692 12870 13748 12908
rect 13020 12238 13022 12290
rect 13074 12238 13076 12290
rect 13020 12226 13076 12238
rect 13468 12292 13524 12302
rect 13468 12178 13524 12236
rect 13468 12126 13470 12178
rect 13522 12126 13524 12178
rect 13468 12114 13524 12126
rect 12684 11342 12686 11394
rect 12738 11342 12740 11394
rect 12684 11330 12740 11342
rect 12908 11732 12964 11742
rect 12908 11282 12964 11676
rect 13804 11396 13860 13804
rect 14140 13794 14196 13804
rect 14476 13746 14532 13758
rect 14476 13694 14478 13746
rect 14530 13694 14532 13746
rect 13916 13300 13972 13310
rect 13916 12850 13972 13244
rect 14252 12964 14308 12974
rect 14252 12870 14308 12908
rect 13916 12798 13918 12850
rect 13970 12798 13972 12850
rect 13916 12786 13972 12798
rect 14028 12852 14084 12862
rect 12908 11230 12910 11282
rect 12962 11230 12964 11282
rect 12908 9826 12964 11230
rect 13580 11340 13804 11396
rect 13468 10836 13524 10846
rect 13468 10610 13524 10780
rect 13468 10558 13470 10610
rect 13522 10558 13524 10610
rect 13468 10546 13524 10558
rect 13132 10388 13188 10398
rect 13132 10294 13188 10332
rect 12908 9774 12910 9826
rect 12962 9774 12964 9826
rect 12908 9762 12964 9774
rect 13468 10052 13524 10062
rect 12572 9622 12628 9660
rect 9884 9266 10052 9268
rect 9884 9214 9886 9266
rect 9938 9214 10052 9266
rect 9884 9212 10052 9214
rect 9884 9202 9940 9212
rect 9996 9044 10052 9054
rect 9772 9042 10052 9044
rect 9772 8990 9998 9042
rect 10050 8990 10052 9042
rect 9772 8988 10052 8990
rect 9996 8978 10052 8988
rect 13468 9042 13524 9996
rect 13580 9156 13636 11340
rect 13804 11330 13860 11340
rect 13916 12066 13972 12078
rect 13916 12014 13918 12066
rect 13970 12014 13972 12066
rect 13916 11060 13972 12014
rect 13916 10994 13972 11004
rect 13916 10612 13972 10622
rect 13916 10050 13972 10556
rect 13916 9998 13918 10050
rect 13970 9998 13972 10050
rect 13916 9986 13972 9998
rect 14028 10052 14084 12796
rect 14476 12068 14532 13694
rect 14588 12962 14644 15148
rect 14700 14642 14756 15372
rect 14700 14590 14702 14642
rect 14754 14590 14756 14642
rect 14700 14578 14756 14590
rect 14924 13972 14980 20132
rect 15036 18338 15092 18350
rect 15036 18286 15038 18338
rect 15090 18286 15092 18338
rect 15036 18116 15092 18286
rect 15036 18050 15092 18060
rect 14924 13906 14980 13916
rect 15148 13858 15204 20972
rect 15260 20132 15316 20142
rect 15260 20038 15316 20076
rect 15372 19012 15428 21534
rect 15372 18946 15428 18956
rect 15484 18676 15540 23492
rect 15708 23426 15764 23436
rect 15596 23156 15652 23166
rect 15820 23156 15876 23884
rect 15932 23380 15988 23390
rect 16380 23380 16436 30492
rect 16492 29652 16548 29662
rect 16492 29558 16548 29596
rect 16716 29540 16772 29550
rect 16716 29426 16772 29484
rect 16716 29374 16718 29426
rect 16770 29374 16772 29426
rect 16716 29362 16772 29374
rect 16828 28532 16884 28542
rect 16828 28438 16884 28476
rect 16492 27860 16548 27870
rect 16492 27188 16548 27804
rect 16940 27748 16996 30828
rect 17052 29876 17108 34188
rect 17500 34132 17556 35646
rect 17724 34914 17780 36540
rect 17836 36530 17892 36540
rect 18508 35700 18564 38892
rect 17724 34862 17726 34914
rect 17778 34862 17780 34914
rect 17724 34850 17780 34862
rect 17836 35644 18564 35700
rect 18620 35700 18676 39676
rect 19068 39508 19124 39518
rect 19180 39508 19236 39676
rect 19404 39620 19460 39630
rect 19404 39526 19460 39564
rect 19068 39506 19236 39508
rect 19068 39454 19070 39506
rect 19122 39454 19236 39506
rect 19068 39452 19236 39454
rect 19068 39442 19124 39452
rect 19068 38834 19124 38846
rect 19068 38782 19070 38834
rect 19122 38782 19124 38834
rect 19068 38276 19124 38782
rect 19628 38834 19684 40684
rect 19852 40404 19908 40414
rect 20188 40404 20244 41918
rect 19852 40402 20244 40404
rect 19852 40350 19854 40402
rect 19906 40350 20244 40402
rect 19852 40348 20244 40350
rect 20300 40404 20356 42700
rect 21868 42700 21980 42756
rect 20748 42642 20804 42654
rect 20748 42590 20750 42642
rect 20802 42590 20804 42642
rect 20412 42532 20468 42542
rect 20412 42438 20468 42476
rect 20748 41076 20804 42590
rect 20636 40404 20692 40414
rect 20300 40348 20636 40404
rect 19852 40338 19908 40348
rect 20524 39394 20580 39406
rect 20524 39342 20526 39394
rect 20578 39342 20580 39394
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19628 38782 19630 38834
rect 19682 38782 19684 38834
rect 19628 38770 19684 38782
rect 20524 38834 20580 39342
rect 20524 38782 20526 38834
rect 20578 38782 20580 38834
rect 20524 38770 20580 38782
rect 19068 38210 19124 38220
rect 19180 38164 19236 38174
rect 18844 38052 18900 38062
rect 18844 37938 18900 37996
rect 19180 38050 19236 38108
rect 20188 38164 20244 38174
rect 20188 38070 20244 38108
rect 19180 37998 19182 38050
rect 19234 37998 19236 38050
rect 19180 37986 19236 37998
rect 20636 38050 20692 40348
rect 20748 40068 20804 41020
rect 21308 40628 21364 40638
rect 20748 40012 21140 40068
rect 20972 38948 21028 38958
rect 20972 38854 21028 38892
rect 21084 38948 21140 40012
rect 21308 39618 21364 40572
rect 21308 39566 21310 39618
rect 21362 39566 21364 39618
rect 21308 39554 21364 39566
rect 21644 40404 21700 40414
rect 21644 39506 21700 40348
rect 21644 39454 21646 39506
rect 21698 39454 21700 39506
rect 21644 39442 21700 39454
rect 21756 39396 21812 39406
rect 21756 39058 21812 39340
rect 21756 39006 21758 39058
rect 21810 39006 21812 39058
rect 21756 38994 21812 39006
rect 21308 38948 21364 38958
rect 21084 38946 21364 38948
rect 21084 38894 21310 38946
rect 21362 38894 21364 38946
rect 21084 38892 21364 38894
rect 20636 37998 20638 38050
rect 20690 37998 20692 38050
rect 20636 37986 20692 37998
rect 18844 37886 18846 37938
rect 18898 37886 18900 37938
rect 18732 37268 18788 37278
rect 18844 37268 18900 37886
rect 19516 37828 19572 37838
rect 19852 37828 19908 37866
rect 19516 37826 19684 37828
rect 19516 37774 19518 37826
rect 19570 37774 19684 37826
rect 19516 37772 19684 37774
rect 19516 37762 19572 37772
rect 18732 37266 18900 37268
rect 18732 37214 18734 37266
rect 18786 37214 18900 37266
rect 18732 37212 18900 37214
rect 18956 37378 19012 37390
rect 18956 37326 18958 37378
rect 19010 37326 19012 37378
rect 18732 37202 18788 37212
rect 18956 37156 19012 37326
rect 19516 37156 19572 37166
rect 18956 37154 19572 37156
rect 18956 37102 19518 37154
rect 19570 37102 19572 37154
rect 18956 37100 19572 37102
rect 19516 36482 19572 37100
rect 19628 37044 19684 37772
rect 19852 37762 19908 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19628 36594 19684 36988
rect 19628 36542 19630 36594
rect 19682 36542 19684 36594
rect 19628 36530 19684 36542
rect 19740 37378 19796 37390
rect 19740 37326 19742 37378
rect 19794 37326 19796 37378
rect 19516 36430 19518 36482
rect 19570 36430 19572 36482
rect 19516 36372 19572 36430
rect 19740 36484 19796 37326
rect 20412 37380 20468 37390
rect 19516 36306 19572 36316
rect 19628 36372 19684 36382
rect 19740 36372 19796 36428
rect 19628 36370 19796 36372
rect 19628 36318 19630 36370
rect 19682 36318 19796 36370
rect 19628 36316 19796 36318
rect 20076 37156 20132 37166
rect 19628 35922 19684 36316
rect 20076 36260 20132 37100
rect 20076 36204 20244 36260
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19628 35870 19630 35922
rect 19682 35870 19684 35922
rect 19628 35858 19684 35870
rect 19964 35924 20020 35934
rect 20188 35924 20244 36204
rect 19964 35922 20244 35924
rect 19964 35870 19966 35922
rect 20018 35870 20244 35922
rect 19964 35868 20244 35870
rect 19964 35858 20020 35868
rect 20412 35700 20468 37324
rect 21084 37156 21140 38892
rect 21308 38882 21364 38892
rect 21868 38668 21924 42700
rect 21980 42662 22036 42700
rect 22092 42084 22148 42094
rect 22092 40402 22148 42028
rect 22092 40350 22094 40402
rect 22146 40350 22148 40402
rect 22092 40338 22148 40350
rect 22092 39732 22148 39742
rect 22316 39732 22372 43374
rect 22428 42754 22484 42766
rect 22428 42702 22430 42754
rect 22482 42702 22484 42754
rect 22428 42084 22484 42702
rect 22876 42756 22932 43484
rect 25340 43540 25396 43550
rect 25340 43446 25396 43484
rect 26124 43538 26180 43550
rect 26124 43486 26126 43538
rect 26178 43486 26180 43538
rect 25788 43426 25844 43438
rect 25788 43374 25790 43426
rect 25842 43374 25844 43426
rect 22876 42754 23268 42756
rect 22876 42702 22878 42754
rect 22930 42702 23268 42754
rect 22876 42700 23268 42702
rect 22876 42690 22932 42700
rect 22428 42018 22484 42028
rect 22988 41972 23044 41982
rect 22652 41970 23044 41972
rect 22652 41918 22990 41970
rect 23042 41918 23044 41970
rect 22652 41916 23044 41918
rect 22428 39732 22484 39742
rect 22316 39730 22484 39732
rect 22316 39678 22430 39730
rect 22482 39678 22484 39730
rect 22316 39676 22484 39678
rect 22092 39638 22148 39676
rect 22428 39666 22484 39676
rect 22204 39396 22260 39406
rect 22204 38836 22260 39340
rect 22428 38948 22484 38958
rect 22652 38948 22708 41916
rect 22988 41906 23044 41916
rect 23212 41188 23268 42700
rect 23324 42754 23380 42766
rect 23324 42702 23326 42754
rect 23378 42702 23380 42754
rect 23324 42644 23380 42702
rect 23324 42578 23380 42588
rect 25564 42642 25620 42654
rect 25564 42590 25566 42642
rect 25618 42590 25620 42642
rect 23436 42084 23492 42094
rect 23436 41970 23492 42028
rect 25564 42084 25620 42590
rect 25564 42018 25620 42028
rect 25676 42532 25732 42542
rect 23436 41918 23438 41970
rect 23490 41918 23492 41970
rect 23436 41906 23492 41918
rect 24108 41972 24164 41982
rect 23436 41188 23492 41198
rect 23212 41186 23492 41188
rect 23212 41134 23438 41186
rect 23490 41134 23492 41186
rect 23212 41132 23492 41134
rect 22876 41076 22932 41086
rect 22876 40982 22932 41020
rect 23212 41074 23268 41132
rect 23436 41122 23492 41132
rect 24108 41186 24164 41916
rect 25676 41970 25732 42476
rect 25676 41918 25678 41970
rect 25730 41918 25732 41970
rect 25676 41906 25732 41918
rect 25788 41972 25844 43374
rect 26124 42756 26180 43486
rect 26124 42690 26180 42700
rect 27244 43314 27300 43326
rect 27244 43262 27246 43314
rect 27298 43262 27300 43314
rect 26684 42642 26740 42654
rect 26684 42590 26686 42642
rect 26738 42590 26740 42642
rect 25788 41906 25844 41916
rect 26460 41972 26516 41982
rect 26460 41878 26516 41916
rect 24220 41748 24276 41758
rect 24220 41746 24500 41748
rect 24220 41694 24222 41746
rect 24274 41694 24500 41746
rect 24220 41692 24500 41694
rect 24220 41682 24276 41692
rect 24108 41134 24110 41186
rect 24162 41134 24164 41186
rect 23212 41022 23214 41074
rect 23266 41022 23268 41074
rect 23212 41010 23268 41022
rect 23996 40964 24052 40974
rect 22764 40516 22820 40526
rect 22764 39620 22820 40460
rect 23884 40404 23940 40414
rect 23100 40180 23156 40190
rect 23100 40178 23268 40180
rect 23100 40126 23102 40178
rect 23154 40126 23268 40178
rect 23100 40124 23268 40126
rect 23100 40114 23156 40124
rect 22764 39618 23156 39620
rect 22764 39566 22766 39618
rect 22818 39566 23156 39618
rect 22764 39564 23156 39566
rect 22764 39554 22820 39564
rect 22428 38946 22708 38948
rect 22428 38894 22430 38946
rect 22482 38894 22708 38946
rect 22428 38892 22708 38894
rect 22428 38882 22484 38892
rect 22204 38742 22260 38780
rect 21644 38612 21924 38668
rect 22540 38668 22596 38892
rect 22540 38612 22820 38668
rect 21308 37940 21364 37950
rect 21308 37846 21364 37884
rect 21644 37828 21700 38612
rect 22428 38276 22484 38286
rect 22092 38164 22148 38174
rect 22092 38162 22372 38164
rect 22092 38110 22094 38162
rect 22146 38110 22372 38162
rect 22092 38108 22372 38110
rect 22092 38098 22148 38108
rect 21644 37492 21700 37772
rect 21644 37426 21700 37436
rect 21084 37090 21140 37100
rect 21308 37378 21364 37390
rect 21308 37326 21310 37378
rect 21362 37326 21364 37378
rect 21308 37044 21364 37326
rect 21308 36978 21364 36988
rect 21980 37154 22036 37166
rect 21980 37102 21982 37154
rect 22034 37102 22036 37154
rect 21644 36484 21700 36494
rect 21644 36390 21700 36428
rect 21868 36482 21924 36494
rect 21868 36430 21870 36482
rect 21922 36430 21924 36482
rect 20748 36372 20804 36382
rect 21868 36372 21924 36430
rect 20748 36370 21252 36372
rect 20748 36318 20750 36370
rect 20802 36318 21252 36370
rect 20748 36316 21252 36318
rect 20748 36306 20804 36316
rect 21196 35810 21252 36316
rect 21196 35758 21198 35810
rect 21250 35758 21252 35810
rect 21196 35746 21252 35758
rect 18620 35644 19124 35700
rect 17836 34242 17892 35644
rect 18284 35476 18340 35486
rect 18284 35382 18340 35420
rect 18620 35476 18676 35486
rect 18620 35474 18900 35476
rect 18620 35422 18622 35474
rect 18674 35422 18900 35474
rect 18620 35420 18900 35422
rect 18620 35410 18676 35420
rect 17836 34190 17838 34242
rect 17890 34190 17892 34242
rect 17836 34178 17892 34190
rect 18172 34242 18228 34254
rect 18172 34190 18174 34242
rect 18226 34190 18228 34242
rect 17500 34066 17556 34076
rect 18172 34132 18228 34190
rect 18172 34066 18228 34076
rect 18396 33908 18452 33918
rect 17164 33906 18452 33908
rect 17164 33854 18398 33906
rect 18450 33854 18452 33906
rect 17164 33852 18452 33854
rect 17164 31666 17220 33852
rect 18396 33842 18452 33852
rect 18732 33906 18788 33918
rect 18732 33854 18734 33906
rect 18786 33854 18788 33906
rect 17612 33684 17668 33694
rect 17276 33348 17332 33358
rect 17276 33254 17332 33292
rect 17164 31614 17166 31666
rect 17218 31614 17220 31666
rect 17164 31602 17220 31614
rect 17276 32562 17332 32574
rect 17276 32510 17278 32562
rect 17330 32510 17332 32562
rect 17276 32228 17332 32510
rect 17164 30100 17220 30110
rect 17276 30100 17332 32172
rect 17612 31780 17668 33628
rect 18060 33122 18116 33134
rect 18060 33070 18062 33122
rect 18114 33070 18116 33122
rect 17612 31686 17668 31724
rect 17948 32562 18004 32574
rect 17948 32510 17950 32562
rect 18002 32510 18004 32562
rect 17948 31668 18004 32510
rect 18060 31780 18116 33070
rect 18732 32004 18788 33854
rect 18732 31938 18788 31948
rect 18172 31780 18228 31790
rect 18060 31778 18228 31780
rect 18060 31726 18174 31778
rect 18226 31726 18228 31778
rect 18060 31724 18228 31726
rect 18172 31714 18228 31724
rect 17948 31602 18004 31612
rect 17612 30884 17668 30894
rect 17668 30828 17780 30884
rect 17612 30790 17668 30828
rect 17164 30098 17332 30100
rect 17164 30046 17166 30098
rect 17218 30046 17332 30098
rect 17164 30044 17332 30046
rect 17388 30212 17444 30222
rect 17164 30034 17220 30044
rect 17052 29820 17220 29876
rect 17052 27748 17108 27758
rect 16940 27692 17052 27748
rect 17052 27682 17108 27692
rect 16604 27636 16660 27646
rect 16604 27542 16660 27580
rect 16492 27094 16548 27132
rect 17052 26964 17108 27002
rect 17052 26898 17108 26908
rect 16940 26852 16996 26862
rect 16940 25618 16996 26796
rect 16940 25566 16942 25618
rect 16994 25566 16996 25618
rect 16940 25554 16996 25566
rect 16716 24722 16772 24734
rect 16716 24670 16718 24722
rect 16770 24670 16772 24722
rect 16716 24164 16772 24670
rect 16828 24498 16884 24510
rect 16828 24446 16830 24498
rect 16882 24446 16884 24498
rect 16828 24164 16884 24446
rect 17164 24388 17220 29820
rect 17388 29650 17444 30156
rect 17388 29598 17390 29650
rect 17442 29598 17444 29650
rect 17388 29586 17444 29598
rect 17724 29652 17780 30828
rect 18508 30882 18564 30894
rect 18508 30830 18510 30882
rect 18562 30830 18564 30882
rect 17836 29988 17892 29998
rect 17836 29894 17892 29932
rect 17724 29538 17780 29596
rect 17724 29486 17726 29538
rect 17778 29486 17780 29538
rect 17724 29474 17780 29486
rect 18508 29540 18564 30830
rect 18508 29474 18564 29484
rect 18396 29204 18452 29214
rect 18732 29204 18788 29214
rect 18284 29202 18452 29204
rect 18284 29150 18398 29202
rect 18450 29150 18452 29202
rect 18284 29148 18452 29150
rect 17388 28532 17444 28542
rect 17388 27074 17444 28476
rect 18284 28084 18340 29148
rect 18396 29138 18452 29148
rect 18508 29202 18788 29204
rect 18508 29150 18734 29202
rect 18786 29150 18788 29202
rect 18508 29148 18788 29150
rect 18396 28756 18452 28766
rect 18508 28756 18564 29148
rect 18732 29138 18788 29148
rect 18396 28754 18564 28756
rect 18396 28702 18398 28754
rect 18450 28702 18564 28754
rect 18396 28700 18564 28702
rect 18396 28690 18452 28700
rect 18284 28018 18340 28028
rect 17612 27970 17668 27982
rect 17612 27918 17614 27970
rect 17666 27918 17668 27970
rect 17500 27860 17556 27870
rect 17500 27766 17556 27804
rect 17388 27022 17390 27074
rect 17442 27022 17444 27074
rect 17388 27010 17444 27022
rect 17500 27188 17556 27198
rect 17164 24322 17220 24332
rect 17500 26290 17556 27132
rect 17612 27186 17668 27918
rect 18284 27636 18340 27646
rect 18284 27542 18340 27580
rect 18620 27636 18676 27646
rect 18620 27542 18676 27580
rect 17612 27134 17614 27186
rect 17666 27134 17668 27186
rect 17612 27122 17668 27134
rect 18732 27300 18788 27310
rect 18732 27074 18788 27244
rect 18732 27022 18734 27074
rect 18786 27022 18788 27074
rect 18732 27010 18788 27022
rect 18620 26964 18676 26974
rect 18844 26962 18900 35420
rect 18956 31780 19012 31790
rect 18956 31218 19012 31724
rect 18956 31166 18958 31218
rect 19010 31166 19012 31218
rect 18956 31154 19012 31166
rect 19068 30996 19124 35644
rect 19180 35586 19236 35598
rect 19180 35534 19182 35586
rect 19234 35534 19236 35586
rect 19180 34132 19236 35534
rect 20412 35586 20468 35644
rect 20412 35534 20414 35586
rect 20466 35534 20468 35586
rect 20412 35522 20468 35534
rect 20860 35698 20916 35710
rect 20860 35646 20862 35698
rect 20914 35646 20916 35698
rect 20860 34692 20916 35646
rect 21532 35700 21588 35710
rect 21532 35606 21588 35644
rect 21868 35476 21924 36316
rect 21980 35698 22036 37102
rect 22316 37044 22372 38108
rect 22428 37492 22484 38220
rect 22540 38050 22596 38612
rect 22540 37998 22542 38050
rect 22594 37998 22596 38050
rect 22540 37986 22596 37998
rect 22540 37492 22596 37502
rect 22428 37490 22596 37492
rect 22428 37438 22542 37490
rect 22594 37438 22596 37490
rect 22428 37436 22596 37438
rect 22092 36932 22148 36942
rect 22092 36482 22148 36876
rect 22092 36430 22094 36482
rect 22146 36430 22148 36482
rect 22092 36372 22148 36430
rect 22092 36306 22148 36316
rect 22316 36706 22372 36988
rect 22316 36654 22318 36706
rect 22370 36654 22372 36706
rect 22204 35812 22260 35822
rect 22204 35718 22260 35756
rect 21980 35646 21982 35698
rect 22034 35646 22036 35698
rect 21980 35634 22036 35646
rect 21868 35420 22148 35476
rect 20860 34626 20916 34636
rect 21756 34692 21812 34702
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19292 34132 19348 34142
rect 19180 34076 19292 34132
rect 19292 34018 19348 34076
rect 19292 33966 19294 34018
rect 19346 33966 19348 34018
rect 19292 33908 19348 33966
rect 19292 33842 19348 33852
rect 21308 33348 21364 33358
rect 21196 33346 21364 33348
rect 21196 33294 21310 33346
rect 21362 33294 21364 33346
rect 21196 33292 21364 33294
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20300 32564 20356 32574
rect 20188 32508 20300 32564
rect 19292 32452 19348 32462
rect 19292 31778 19348 32396
rect 19292 31726 19294 31778
rect 19346 31726 19348 31778
rect 19292 31714 19348 31726
rect 19404 31892 19460 31902
rect 18844 26910 18846 26962
rect 18898 26910 18900 26962
rect 18620 26852 18788 26908
rect 18844 26898 18900 26910
rect 18956 30940 19124 30996
rect 17500 26238 17502 26290
rect 17554 26238 17556 26290
rect 17500 24164 17556 26238
rect 17948 26516 18004 26526
rect 17948 26290 18004 26460
rect 17948 26238 17950 26290
rect 18002 26238 18004 26290
rect 17948 26226 18004 26238
rect 18620 26290 18676 26302
rect 18620 26238 18622 26290
rect 18674 26238 18676 26290
rect 18620 26180 18676 26238
rect 18620 26114 18676 26124
rect 18508 26068 18564 26078
rect 18508 25974 18564 26012
rect 17612 25956 17668 25966
rect 17612 25506 17668 25900
rect 18060 25508 18116 25518
rect 17612 25454 17614 25506
rect 17666 25454 17668 25506
rect 17612 25442 17668 25454
rect 17948 25506 18116 25508
rect 17948 25454 18062 25506
rect 18114 25454 18116 25506
rect 17948 25452 18116 25454
rect 17724 25396 17780 25406
rect 17724 25302 17780 25340
rect 17836 24722 17892 24734
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 17836 24164 17892 24670
rect 16828 24108 17892 24164
rect 16716 24098 16772 24108
rect 15932 23378 16436 23380
rect 15932 23326 15934 23378
rect 15986 23326 16436 23378
rect 15932 23324 16436 23326
rect 15932 23314 15988 23324
rect 15820 23100 16100 23156
rect 15596 23062 15652 23100
rect 15708 22820 15764 22830
rect 16044 22820 16100 23100
rect 16380 23154 16436 23324
rect 16380 23102 16382 23154
rect 16434 23102 16436 23154
rect 16380 23090 16436 23102
rect 16492 23826 16548 23838
rect 16492 23774 16494 23826
rect 16546 23774 16548 23826
rect 15764 22764 15876 22820
rect 16044 22764 16436 22820
rect 15708 22754 15764 22764
rect 15708 22484 15764 22494
rect 15708 22390 15764 22428
rect 15820 22370 15876 22764
rect 15820 22318 15822 22370
rect 15874 22318 15876 22370
rect 15820 22306 15876 22318
rect 16380 22370 16436 22764
rect 16492 22484 16548 23774
rect 16604 23266 16660 23278
rect 16604 23214 16606 23266
rect 16658 23214 16660 23266
rect 16604 23044 16660 23214
rect 16604 22978 16660 22988
rect 17388 23154 17444 23166
rect 17388 23102 17390 23154
rect 17442 23102 17444 23154
rect 16492 22418 16548 22428
rect 16380 22318 16382 22370
rect 16434 22318 16436 22370
rect 16044 22260 16100 22270
rect 16044 22258 16324 22260
rect 16044 22206 16046 22258
rect 16098 22206 16324 22258
rect 16044 22204 16324 22206
rect 16044 22194 16100 22204
rect 15596 22146 15652 22158
rect 15596 22094 15598 22146
rect 15650 22094 15652 22146
rect 15596 19346 15652 22094
rect 15708 22036 15764 22046
rect 15708 21586 15764 21980
rect 16044 22036 16100 22046
rect 16044 21810 16100 21980
rect 16044 21758 16046 21810
rect 16098 21758 16100 21810
rect 16044 21746 16100 21758
rect 15932 21588 15988 21598
rect 15708 21534 15710 21586
rect 15762 21534 15764 21586
rect 15708 21522 15764 21534
rect 15820 21586 15988 21588
rect 15820 21534 15934 21586
rect 15986 21534 15988 21586
rect 15820 21532 15988 21534
rect 15596 19294 15598 19346
rect 15650 19294 15652 19346
rect 15596 18788 15652 19294
rect 15708 19796 15764 19806
rect 15820 19796 15876 21532
rect 15932 21522 15988 21532
rect 16156 21588 16212 21598
rect 16268 21588 16324 22204
rect 16380 21812 16436 22318
rect 17164 22258 17220 22270
rect 17164 22206 17166 22258
rect 17218 22206 17220 22258
rect 17164 21924 17220 22206
rect 17164 21858 17220 21868
rect 16380 21756 16548 21812
rect 16492 21700 16548 21756
rect 16492 21634 16548 21644
rect 16828 21700 16884 21710
rect 16828 21606 16884 21644
rect 16380 21588 16436 21598
rect 16268 21586 16436 21588
rect 16268 21534 16382 21586
rect 16434 21534 16436 21586
rect 16268 21532 16436 21534
rect 16156 21494 16212 21532
rect 16044 20692 16100 20702
rect 16044 20598 16100 20636
rect 15764 19740 15876 19796
rect 15932 20580 15988 20590
rect 15708 19458 15764 19740
rect 15708 19406 15710 19458
rect 15762 19406 15764 19458
rect 15708 19348 15764 19406
rect 15708 19282 15764 19292
rect 15932 19234 15988 20524
rect 15932 19182 15934 19234
rect 15986 19182 15988 19234
rect 15932 19170 15988 19182
rect 16268 19122 16324 19134
rect 16268 19070 16270 19122
rect 16322 19070 16324 19122
rect 15596 18722 15652 18732
rect 15932 18900 15988 18910
rect 15372 18620 15484 18676
rect 15372 17668 15428 18620
rect 15484 18610 15540 18620
rect 15484 18450 15540 18462
rect 15484 18398 15486 18450
rect 15538 18398 15540 18450
rect 15484 18228 15540 18398
rect 15932 18450 15988 18844
rect 15932 18398 15934 18450
rect 15986 18398 15988 18450
rect 15484 18162 15540 18172
rect 15708 18340 15764 18350
rect 15260 17612 15372 17668
rect 15260 16210 15316 17612
rect 15372 17602 15428 17612
rect 15708 16994 15764 18284
rect 15932 17444 15988 18398
rect 15932 17378 15988 17388
rect 16268 17108 16324 19070
rect 16380 19012 16436 21532
rect 17388 21364 17444 23102
rect 17836 22372 17892 24108
rect 17836 22306 17892 22316
rect 17948 23156 18004 25452
rect 18060 25442 18116 25452
rect 18508 25506 18564 25518
rect 18508 25454 18510 25506
rect 18562 25454 18564 25506
rect 18172 24610 18228 24622
rect 18172 24558 18174 24610
rect 18226 24558 18228 24610
rect 18172 23716 18228 24558
rect 18172 23650 18228 23660
rect 18508 23268 18564 25454
rect 18620 24724 18676 24734
rect 18620 24630 18676 24668
rect 18620 24164 18676 24174
rect 18620 24050 18676 24108
rect 18620 23998 18622 24050
rect 18674 23998 18676 24050
rect 18620 23986 18676 23998
rect 18508 23202 18564 23212
rect 17948 22148 18004 23100
rect 17612 22092 18004 22148
rect 18172 23042 18228 23054
rect 18172 22990 18174 23042
rect 18226 22990 18228 23042
rect 17612 21698 17668 22092
rect 18172 22036 18228 22990
rect 18172 21970 18228 21980
rect 18396 22260 18452 22270
rect 17612 21646 17614 21698
rect 17666 21646 17668 21698
rect 17612 21634 17668 21646
rect 17836 21812 17892 21822
rect 17500 21588 17556 21598
rect 17500 21494 17556 21532
rect 17388 21298 17444 21308
rect 16828 20916 16884 20926
rect 16828 20804 16884 20860
rect 17164 20804 17220 20814
rect 16828 20802 16996 20804
rect 16828 20750 16830 20802
rect 16882 20750 16996 20802
rect 16828 20748 16996 20750
rect 16828 20738 16884 20748
rect 16716 20020 16772 20030
rect 16716 19796 16772 19964
rect 16716 19730 16772 19740
rect 16380 18946 16436 18956
rect 16604 19234 16660 19246
rect 16604 19182 16606 19234
rect 16658 19182 16660 19234
rect 16380 18676 16436 18686
rect 16380 18450 16436 18620
rect 16380 18398 16382 18450
rect 16434 18398 16436 18450
rect 16380 18386 16436 18398
rect 16604 17780 16660 19182
rect 16716 19124 16772 19134
rect 16716 19030 16772 19068
rect 16828 19122 16884 19134
rect 16828 19070 16830 19122
rect 16882 19070 16884 19122
rect 16828 19012 16884 19070
rect 16828 18946 16884 18956
rect 16940 18564 16996 20748
rect 17164 20710 17220 20748
rect 17836 20802 17892 21756
rect 18396 21588 18452 22204
rect 18396 21522 18452 21532
rect 18060 21474 18116 21486
rect 18060 21422 18062 21474
rect 18114 21422 18116 21474
rect 18060 21364 18116 21422
rect 18060 21298 18116 21308
rect 18284 21476 18340 21486
rect 17836 20750 17838 20802
rect 17890 20750 17892 20802
rect 17836 20738 17892 20750
rect 17276 20692 17332 20702
rect 17276 20598 17332 20636
rect 17388 20580 17444 20590
rect 17388 20486 17444 20524
rect 17388 20132 17444 20142
rect 17388 20038 17444 20076
rect 17612 20018 17668 20030
rect 17612 19966 17614 20018
rect 17666 19966 17668 20018
rect 17612 19460 17668 19966
rect 18172 20018 18228 20030
rect 18172 19966 18174 20018
rect 18226 19966 18228 20018
rect 17612 19394 17668 19404
rect 18060 19794 18116 19806
rect 18060 19742 18062 19794
rect 18114 19742 18116 19794
rect 17164 19234 17220 19246
rect 17164 19182 17166 19234
rect 17218 19182 17220 19234
rect 17164 18564 17220 19182
rect 17948 19124 18004 19134
rect 17948 19030 18004 19068
rect 18060 18788 18116 19742
rect 18172 19796 18228 19966
rect 18172 19730 18228 19740
rect 18060 18722 18116 18732
rect 16604 17714 16660 17724
rect 16716 18508 17220 18564
rect 17836 18564 17892 18574
rect 16268 17042 16324 17052
rect 15708 16942 15710 16994
rect 15762 16942 15764 16994
rect 15708 16930 15764 16942
rect 16380 16884 16436 16894
rect 16716 16884 16772 18508
rect 17388 18452 17444 18462
rect 16940 18450 17444 18452
rect 16940 18398 17390 18450
rect 17442 18398 17444 18450
rect 16940 18396 17444 18398
rect 16828 18338 16884 18350
rect 16828 18286 16830 18338
rect 16882 18286 16884 18338
rect 16828 18228 16884 18286
rect 16828 18162 16884 18172
rect 16940 17778 16996 18396
rect 17388 18386 17444 18396
rect 17612 18340 17668 18350
rect 16940 17726 16942 17778
rect 16994 17726 16996 17778
rect 16940 17714 16996 17726
rect 17500 18284 17612 18340
rect 16436 16828 16772 16884
rect 17388 17444 17444 17454
rect 16380 16790 16436 16828
rect 15260 16158 15262 16210
rect 15314 16158 15316 16210
rect 15260 15428 15316 16158
rect 15932 16660 15988 16670
rect 15932 15988 15988 16604
rect 16604 16660 16660 16670
rect 16604 16322 16660 16604
rect 16604 16270 16606 16322
rect 16658 16270 16660 16322
rect 16604 16258 16660 16270
rect 16268 16098 16324 16110
rect 16268 16046 16270 16098
rect 16322 16046 16324 16098
rect 16268 15988 16324 16046
rect 17388 16100 17444 17388
rect 17500 16882 17556 18284
rect 17612 18274 17668 18284
rect 17836 18116 17892 18508
rect 18172 18452 18228 18462
rect 18172 18358 18228 18396
rect 17948 18338 18004 18350
rect 17948 18286 17950 18338
rect 18002 18286 18004 18338
rect 17948 18228 18004 18286
rect 17948 18162 18004 18172
rect 17836 17780 17892 18060
rect 17948 17780 18004 17790
rect 17836 17778 18004 17780
rect 17836 17726 17950 17778
rect 18002 17726 18004 17778
rect 17836 17724 18004 17726
rect 17948 17714 18004 17724
rect 18060 17108 18116 17118
rect 18060 17014 18116 17052
rect 17500 16830 17502 16882
rect 17554 16830 17556 16882
rect 17500 16818 17556 16830
rect 17724 16660 17780 16670
rect 17388 16034 17444 16044
rect 17500 16212 17556 16222
rect 15932 15986 16324 15988
rect 15932 15934 15934 15986
rect 15986 15934 16324 15986
rect 15932 15932 16324 15934
rect 15932 15922 15988 15932
rect 16268 15540 16324 15932
rect 16268 15474 16324 15484
rect 16828 15540 16884 15550
rect 16828 15446 16884 15484
rect 17500 15540 17556 16156
rect 15260 15362 15316 15372
rect 17500 15314 17556 15484
rect 17500 15262 17502 15314
rect 17554 15262 17556 15314
rect 17500 15250 17556 15262
rect 17724 15314 17780 16604
rect 17724 15262 17726 15314
rect 17778 15262 17780 15314
rect 17724 15250 17780 15262
rect 18172 15876 18228 15886
rect 16828 14756 16884 14766
rect 16828 14642 16884 14700
rect 16828 14590 16830 14642
rect 16882 14590 16884 14642
rect 16828 14578 16884 14590
rect 18172 14306 18228 15820
rect 18284 14644 18340 21420
rect 18620 20018 18676 20030
rect 18620 19966 18622 20018
rect 18674 19966 18676 20018
rect 18508 19794 18564 19806
rect 18508 19742 18510 19794
rect 18562 19742 18564 19794
rect 18508 19348 18564 19742
rect 18620 19684 18676 19966
rect 18620 19618 18676 19628
rect 18508 19282 18564 19292
rect 18396 18562 18452 18574
rect 18396 18510 18398 18562
rect 18450 18510 18452 18562
rect 18396 17556 18452 18510
rect 18508 18564 18564 18574
rect 18508 18470 18564 18508
rect 18396 17490 18452 17500
rect 18620 17780 18676 17790
rect 18732 17780 18788 26852
rect 18844 26290 18900 26302
rect 18844 26238 18846 26290
rect 18898 26238 18900 26290
rect 18844 25172 18900 26238
rect 18844 25106 18900 25116
rect 18956 18900 19012 30940
rect 19404 29540 19460 31836
rect 19852 31780 19908 31790
rect 19852 31686 19908 31724
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20188 30994 20244 32508
rect 20300 32498 20356 32508
rect 20412 32452 20468 32462
rect 20412 32358 20468 32396
rect 20188 30942 20190 30994
rect 20242 30942 20244 30994
rect 20188 30324 20244 30942
rect 20412 32228 20468 32238
rect 20412 31666 20468 32172
rect 21196 32116 21252 33292
rect 21308 33282 21364 33292
rect 21644 33348 21700 33358
rect 21420 33236 21476 33246
rect 21420 32564 21476 33180
rect 21420 32470 21476 32508
rect 21644 32562 21700 33292
rect 21644 32510 21646 32562
rect 21698 32510 21700 32562
rect 21196 32050 21252 32060
rect 21308 32338 21364 32350
rect 21308 32286 21310 32338
rect 21362 32286 21364 32338
rect 20972 32004 21028 32014
rect 21028 31948 21140 32004
rect 20972 31938 21028 31948
rect 20412 31614 20414 31666
rect 20466 31614 20468 31666
rect 20412 30882 20468 31614
rect 20748 31554 20804 31566
rect 20748 31502 20750 31554
rect 20802 31502 20804 31554
rect 20748 31220 20804 31502
rect 20748 31154 20804 31164
rect 20412 30830 20414 30882
rect 20466 30830 20468 30882
rect 20412 30818 20468 30830
rect 20412 30324 20468 30334
rect 20188 30322 20468 30324
rect 20188 30270 20414 30322
rect 20466 30270 20468 30322
rect 20188 30268 20468 30270
rect 19516 30212 19572 30250
rect 19516 30146 19572 30156
rect 20076 30210 20132 30222
rect 20076 30158 20078 30210
rect 20130 30158 20132 30210
rect 19292 29484 19460 29540
rect 19516 29986 19572 29998
rect 19516 29934 19518 29986
rect 19570 29934 19572 29986
rect 19516 29538 19572 29934
rect 19516 29486 19518 29538
rect 19570 29486 19572 29538
rect 19180 29426 19236 29438
rect 19180 29374 19182 29426
rect 19234 29374 19236 29426
rect 19180 28642 19236 29374
rect 19180 28590 19182 28642
rect 19234 28590 19236 28642
rect 19068 28530 19124 28542
rect 19068 28478 19070 28530
rect 19122 28478 19124 28530
rect 19068 27970 19124 28478
rect 19068 27918 19070 27970
rect 19122 27918 19124 27970
rect 19068 27906 19124 27918
rect 19180 27860 19236 28590
rect 19180 27794 19236 27804
rect 19292 27748 19348 29484
rect 19516 29474 19572 29486
rect 19628 29988 19684 29998
rect 20076 29988 20132 30158
rect 20188 30212 20244 30268
rect 20412 30258 20468 30268
rect 20188 30146 20244 30156
rect 20076 29932 20244 29988
rect 19404 29316 19460 29326
rect 19404 27970 19460 29260
rect 19628 28866 19684 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20188 29764 20244 29932
rect 20300 29764 20356 29774
rect 20188 29708 20300 29764
rect 19628 28814 19630 28866
rect 19682 28814 19684 28866
rect 19628 28802 19684 28814
rect 20076 29314 20132 29326
rect 20076 29262 20078 29314
rect 20130 29262 20132 29314
rect 19964 28420 20020 28458
rect 20076 28420 20132 29262
rect 20188 29316 20244 29708
rect 20300 29698 20356 29708
rect 20188 29250 20244 29260
rect 20524 29426 20580 29438
rect 20524 29374 20526 29426
rect 20578 29374 20580 29426
rect 20076 28364 20244 28420
rect 19964 28354 20020 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19404 27918 19406 27970
rect 19458 27918 19460 27970
rect 19404 27906 19460 27918
rect 20188 27858 20244 28364
rect 20188 27806 20190 27858
rect 20242 27806 20244 27858
rect 19292 27692 19684 27748
rect 19516 27412 19572 27422
rect 19404 27076 19460 27086
rect 19404 26982 19460 27020
rect 19292 26962 19348 26974
rect 19292 26910 19294 26962
rect 19346 26910 19348 26962
rect 19180 26852 19236 26862
rect 19068 26850 19236 26852
rect 19068 26798 19182 26850
rect 19234 26798 19236 26850
rect 19068 26796 19236 26798
rect 19068 25506 19124 26796
rect 19180 26786 19236 26796
rect 19292 26740 19348 26910
rect 19292 26674 19348 26684
rect 19516 26516 19572 27356
rect 19068 25454 19070 25506
rect 19122 25454 19124 25506
rect 19068 25442 19124 25454
rect 19180 26460 19572 26516
rect 19180 24946 19236 26460
rect 19628 26404 19684 27692
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19180 24894 19182 24946
rect 19234 24894 19236 24946
rect 19180 24882 19236 24894
rect 19292 26348 19684 26404
rect 19740 26514 19796 26526
rect 19740 26462 19742 26514
rect 19794 26462 19796 26514
rect 19292 24276 19348 26348
rect 19404 26180 19460 26190
rect 19740 26180 19796 26462
rect 19404 26178 19796 26180
rect 19404 26126 19406 26178
rect 19458 26126 19796 26178
rect 19404 26124 19796 26126
rect 20188 26290 20244 27806
rect 20524 27076 20580 29374
rect 20860 29428 20916 29438
rect 20860 29334 20916 29372
rect 20860 28420 20916 28430
rect 20524 26982 20580 27020
rect 20748 28084 20804 28094
rect 20188 26238 20190 26290
rect 20242 26238 20244 26290
rect 19404 26114 19460 26124
rect 18956 18834 19012 18844
rect 19068 24220 19348 24276
rect 19404 25506 19460 25518
rect 19404 25454 19406 25506
rect 19458 25454 19460 25506
rect 19404 25172 19460 25454
rect 19852 25508 19908 25518
rect 19852 25414 19908 25452
rect 18620 17778 19012 17780
rect 18620 17726 18622 17778
rect 18674 17726 19012 17778
rect 18620 17724 19012 17726
rect 18620 17220 18676 17724
rect 18956 17666 19012 17724
rect 18956 17614 18958 17666
rect 19010 17614 19012 17666
rect 18956 17602 19012 17614
rect 18284 14578 18340 14588
rect 18396 17164 18676 17220
rect 18732 17556 18788 17566
rect 18172 14254 18174 14306
rect 18226 14254 18228 14306
rect 18172 14196 18228 14254
rect 17500 14140 18228 14196
rect 15148 13806 15150 13858
rect 15202 13806 15204 13858
rect 14812 13748 14868 13758
rect 14812 13654 14868 13692
rect 14588 12910 14590 12962
rect 14642 12910 14644 12962
rect 14588 12898 14644 12910
rect 14924 13076 14980 13086
rect 14924 12850 14980 13020
rect 15148 12964 15204 13806
rect 15820 13858 15876 13870
rect 15820 13806 15822 13858
rect 15874 13806 15876 13858
rect 15484 13746 15540 13758
rect 15484 13694 15486 13746
rect 15538 13694 15540 13746
rect 15148 12898 15204 12908
rect 15260 12962 15316 12974
rect 15260 12910 15262 12962
rect 15314 12910 15316 12962
rect 14924 12798 14926 12850
rect 14978 12798 14980 12850
rect 14924 12786 14980 12798
rect 14476 12002 14532 12012
rect 14364 11956 14420 11966
rect 14140 11060 14196 11070
rect 14140 10052 14196 11004
rect 14364 10610 14420 11900
rect 15036 11956 15092 11966
rect 14700 11396 14756 11406
rect 14700 11394 14980 11396
rect 14700 11342 14702 11394
rect 14754 11342 14980 11394
rect 14700 11340 14980 11342
rect 14700 11330 14756 11340
rect 14700 11060 14756 11070
rect 14756 11004 14868 11060
rect 14700 10994 14756 11004
rect 14812 10722 14868 11004
rect 14812 10670 14814 10722
rect 14866 10670 14868 10722
rect 14812 10658 14868 10670
rect 14364 10558 14366 10610
rect 14418 10558 14420 10610
rect 14364 10546 14420 10558
rect 14924 10612 14980 11340
rect 15036 11394 15092 11900
rect 15260 11956 15316 12910
rect 15484 12852 15540 13694
rect 15820 13188 15876 13806
rect 15820 12962 15876 13132
rect 16940 13188 16996 13198
rect 16940 13094 16996 13132
rect 16492 13076 16548 13086
rect 15820 12910 15822 12962
rect 15874 12910 15876 12962
rect 15820 12898 15876 12910
rect 16380 12964 16436 12974
rect 15484 12786 15540 12796
rect 15260 11890 15316 11900
rect 15372 12068 15428 12078
rect 15036 11342 15038 11394
rect 15090 11342 15092 11394
rect 15036 11330 15092 11342
rect 14924 10546 14980 10556
rect 14252 10052 14308 10062
rect 14140 10050 14420 10052
rect 14140 9998 14254 10050
rect 14306 9998 14420 10050
rect 14140 9996 14420 9998
rect 14028 9958 14084 9996
rect 14252 9986 14308 9996
rect 13580 9154 13748 9156
rect 13580 9102 13582 9154
rect 13634 9102 13748 9154
rect 13580 9100 13748 9102
rect 13580 9090 13636 9100
rect 13468 8990 13470 9042
rect 13522 8990 13524 9042
rect 13468 8372 13524 8990
rect 13580 8372 13636 8382
rect 13468 8370 13636 8372
rect 13468 8318 13582 8370
rect 13634 8318 13636 8370
rect 13468 8316 13636 8318
rect 13580 8306 13636 8316
rect 13692 8258 13748 9100
rect 14364 9042 14420 9996
rect 14812 9716 14868 9726
rect 15148 9716 15204 9726
rect 14812 9714 15204 9716
rect 14812 9662 14814 9714
rect 14866 9662 15150 9714
rect 15202 9662 15204 9714
rect 14812 9660 15204 9662
rect 14812 9650 14868 9660
rect 15148 9650 15204 9660
rect 14364 8990 14366 9042
rect 14418 8990 14420 9042
rect 14364 8428 14420 8990
rect 14476 8932 14532 8942
rect 14476 8838 14532 8876
rect 13692 8206 13694 8258
rect 13746 8206 13748 8258
rect 13692 8194 13748 8206
rect 14252 8372 14420 8428
rect 14252 8260 14308 8372
rect 14252 8194 14308 8204
rect 15036 8260 15092 8270
rect 15036 8166 15092 8204
rect 5516 7646 5518 7698
rect 5570 7646 5572 7698
rect 5516 7634 5572 7646
rect 5852 6916 5908 6926
rect 5068 6132 5124 6142
rect 4956 6130 5124 6132
rect 4956 6078 5070 6130
rect 5122 6078 5124 6130
rect 4956 6076 5124 6078
rect 5068 6066 5124 6076
rect 5852 6130 5908 6860
rect 15372 6692 15428 12012
rect 15484 11844 15540 11854
rect 15484 9826 15540 11788
rect 16380 11844 16436 12908
rect 16492 12178 16548 13020
rect 16492 12126 16494 12178
rect 16546 12126 16548 12178
rect 16492 12114 16548 12126
rect 16716 12850 16772 12862
rect 16716 12798 16718 12850
rect 16770 12798 16772 12850
rect 15708 11396 15764 11406
rect 15708 11282 15764 11340
rect 16380 11394 16436 11788
rect 16380 11342 16382 11394
rect 16434 11342 16436 11394
rect 16380 11330 16436 11342
rect 16044 11284 16100 11294
rect 15708 11230 15710 11282
rect 15762 11230 15764 11282
rect 15708 11218 15764 11230
rect 15820 11282 16100 11284
rect 15820 11230 16046 11282
rect 16098 11230 16100 11282
rect 15820 11228 16100 11230
rect 15484 9774 15486 9826
rect 15538 9774 15540 9826
rect 15484 8260 15540 9774
rect 15596 9156 15652 9166
rect 15820 9156 15876 11228
rect 16044 11218 16100 11228
rect 16716 10836 16772 12798
rect 17276 12740 17332 12750
rect 17276 12646 17332 12684
rect 17052 12292 17108 12302
rect 16828 11396 16884 11406
rect 16828 11302 16884 11340
rect 17052 11282 17108 12236
rect 17052 11230 17054 11282
rect 17106 11230 17108 11282
rect 17052 11218 17108 11230
rect 17500 11282 17556 14140
rect 18396 14084 18452 17164
rect 18732 17108 18788 17500
rect 18732 16770 18788 17052
rect 18732 16718 18734 16770
rect 18786 16718 18788 16770
rect 18732 16706 18788 16718
rect 18732 16548 18788 16558
rect 18620 15988 18676 15998
rect 18620 14642 18676 15932
rect 18620 14590 18622 14642
rect 18674 14590 18676 14642
rect 18620 14578 18676 14590
rect 18172 14028 18452 14084
rect 17612 13972 17668 13982
rect 17836 13972 17892 13982
rect 17612 13634 17668 13916
rect 17612 13582 17614 13634
rect 17666 13582 17668 13634
rect 17612 13412 17668 13582
rect 17612 13346 17668 13356
rect 17724 13916 17836 13972
rect 17724 12962 17780 13916
rect 17836 13906 17892 13916
rect 17948 13860 18004 13870
rect 17948 13858 18116 13860
rect 17948 13806 17950 13858
rect 18002 13806 18116 13858
rect 17948 13804 18116 13806
rect 17948 13794 18004 13804
rect 18060 12964 18116 13804
rect 17724 12910 17726 12962
rect 17778 12910 17780 12962
rect 17724 12898 17780 12910
rect 17836 12908 18116 12964
rect 18172 13074 18228 14028
rect 18732 13972 18788 16492
rect 19068 16548 19124 24220
rect 19292 24052 19348 24062
rect 19292 23958 19348 23996
rect 19404 23940 19460 25116
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 25060 20244 26238
rect 20748 26292 20804 28028
rect 20860 27858 20916 28364
rect 21084 28308 21140 31948
rect 21308 31890 21364 32286
rect 21644 32228 21700 32510
rect 21644 32162 21700 32172
rect 21756 33346 21812 34636
rect 21980 34692 22036 34702
rect 21980 34598 22036 34636
rect 22092 34580 22148 35420
rect 22092 34514 22148 34524
rect 22204 35252 22260 35262
rect 22092 34244 22148 34254
rect 21980 34242 22148 34244
rect 21980 34190 22094 34242
rect 22146 34190 22148 34242
rect 21980 34188 22148 34190
rect 21868 33684 21924 33694
rect 21980 33684 22036 34188
rect 22092 34178 22148 34188
rect 21924 33628 22036 33684
rect 21868 33618 21924 33628
rect 22204 33572 22260 35196
rect 22316 33908 22372 36654
rect 22428 36372 22484 36382
rect 22428 34580 22484 36316
rect 22540 36260 22596 37436
rect 22764 36932 22820 38612
rect 22876 38610 22932 38622
rect 22876 38558 22878 38610
rect 22930 38558 22932 38610
rect 22876 37492 22932 38558
rect 22988 38052 23044 38062
rect 22988 37958 23044 37996
rect 22876 37436 23044 37492
rect 22764 36866 22820 36876
rect 22876 37266 22932 37278
rect 22876 37214 22878 37266
rect 22930 37214 22932 37266
rect 22876 36484 22932 37214
rect 22540 36194 22596 36204
rect 22652 36428 22932 36484
rect 22652 35028 22708 36428
rect 22764 36258 22820 36270
rect 22764 36206 22766 36258
rect 22818 36206 22820 36258
rect 22764 35028 22820 36206
rect 22876 36260 22932 36270
rect 22876 35698 22932 36204
rect 22876 35646 22878 35698
rect 22930 35646 22932 35698
rect 22876 35476 22932 35646
rect 22876 35410 22932 35420
rect 22876 35252 22932 35262
rect 22988 35252 23044 37436
rect 22932 35196 23044 35252
rect 22876 35186 22932 35196
rect 22876 35028 22932 35038
rect 22764 35026 22932 35028
rect 22764 34974 22878 35026
rect 22930 34974 22932 35026
rect 22764 34972 22932 34974
rect 22652 34962 22708 34972
rect 22876 34962 22932 34972
rect 23100 34916 23156 39564
rect 23212 39618 23268 40124
rect 23212 39566 23214 39618
rect 23266 39566 23268 39618
rect 23212 39554 23268 39566
rect 23436 39396 23492 39406
rect 23212 39394 23492 39396
rect 23212 39342 23438 39394
rect 23490 39342 23492 39394
rect 23212 39340 23492 39342
rect 23212 38834 23268 39340
rect 23436 39330 23492 39340
rect 23212 38782 23214 38834
rect 23266 38782 23268 38834
rect 23212 38770 23268 38782
rect 23772 38834 23828 38846
rect 23772 38782 23774 38834
rect 23826 38782 23828 38834
rect 23772 38276 23828 38782
rect 23772 38210 23828 38220
rect 23884 38164 23940 40348
rect 23996 38946 24052 40908
rect 24108 40626 24164 41134
rect 24108 40574 24110 40626
rect 24162 40574 24164 40626
rect 24108 40562 24164 40574
rect 23996 38894 23998 38946
rect 24050 38894 24052 38946
rect 23996 38882 24052 38894
rect 24108 39618 24164 39630
rect 24108 39566 24110 39618
rect 24162 39566 24164 39618
rect 24108 38724 24164 39566
rect 24444 39618 24500 41692
rect 25564 41412 25620 41422
rect 24444 39566 24446 39618
rect 24498 39566 24500 39618
rect 24444 39554 24500 39566
rect 25452 40404 25508 40414
rect 24108 38658 24164 38668
rect 24556 38722 24612 38734
rect 24556 38670 24558 38722
rect 24610 38670 24612 38722
rect 24556 38276 24612 38670
rect 25452 38724 25508 40348
rect 25564 39618 25620 41356
rect 25564 39566 25566 39618
rect 25618 39566 25620 39618
rect 25564 39554 25620 39566
rect 26348 41186 26404 41198
rect 26348 41134 26350 41186
rect 26402 41134 26404 41186
rect 25452 38612 25732 38668
rect 24556 38210 24612 38220
rect 23884 38108 24164 38164
rect 23436 38050 23492 38062
rect 23436 37998 23438 38050
rect 23490 37998 23492 38050
rect 23436 37828 23492 37998
rect 23884 37940 23940 37950
rect 23436 37266 23492 37772
rect 23436 37214 23438 37266
rect 23490 37214 23492 37266
rect 23324 35698 23380 35710
rect 23324 35646 23326 35698
rect 23378 35646 23380 35698
rect 23212 34916 23268 34926
rect 22988 34914 23268 34916
rect 22988 34862 23214 34914
rect 23266 34862 23268 34914
rect 22988 34860 23268 34862
rect 22540 34804 22596 34814
rect 22988 34804 23044 34860
rect 23212 34850 23268 34860
rect 22540 34802 23044 34804
rect 22540 34750 22542 34802
rect 22594 34750 23044 34802
rect 22540 34748 23044 34750
rect 22540 34738 22596 34748
rect 23212 34580 23268 34590
rect 22428 34524 23044 34580
rect 22428 34244 22484 34254
rect 22428 34150 22484 34188
rect 22876 33908 22932 33918
rect 22316 33906 22932 33908
rect 22316 33854 22878 33906
rect 22930 33854 22932 33906
rect 22316 33852 22932 33854
rect 22876 33842 22932 33852
rect 22988 33906 23044 34524
rect 23212 34130 23268 34524
rect 23324 34354 23380 35646
rect 23324 34302 23326 34354
rect 23378 34302 23380 34354
rect 23324 34290 23380 34302
rect 23212 34078 23214 34130
rect 23266 34078 23268 34130
rect 23212 34066 23268 34078
rect 23436 34130 23492 37214
rect 23772 37938 23940 37940
rect 23772 37886 23886 37938
rect 23938 37886 23940 37938
rect 23772 37884 23940 37886
rect 23548 37044 23604 37054
rect 23548 36370 23604 36988
rect 23548 36318 23550 36370
rect 23602 36318 23604 36370
rect 23548 36306 23604 36318
rect 23436 34078 23438 34130
rect 23490 34078 23492 34130
rect 23436 34066 23492 34078
rect 23548 35812 23604 35822
rect 22988 33854 22990 33906
rect 23042 33854 23044 33906
rect 22988 33842 23044 33854
rect 23212 33908 23268 33918
rect 21756 33294 21758 33346
rect 21810 33294 21812 33346
rect 21756 32004 21812 33294
rect 21308 31838 21310 31890
rect 21362 31838 21364 31890
rect 21308 31826 21364 31838
rect 21420 31948 21812 32004
rect 21980 33516 22260 33572
rect 22652 33684 22708 33694
rect 21420 30098 21476 31948
rect 21756 31780 21812 31790
rect 21756 31686 21812 31724
rect 21644 31668 21700 31678
rect 21644 31106 21700 31612
rect 21644 31054 21646 31106
rect 21698 31054 21700 31106
rect 21644 31042 21700 31054
rect 21980 30884 22036 33516
rect 22428 33348 22484 33358
rect 22428 33254 22484 33292
rect 22204 33236 22260 33246
rect 22204 33142 22260 33180
rect 22204 32676 22260 32686
rect 22204 32582 22260 32620
rect 22540 32674 22596 32686
rect 22540 32622 22542 32674
rect 22594 32622 22596 32674
rect 22204 32340 22260 32350
rect 22092 31892 22148 31902
rect 22092 31790 22148 31836
rect 22092 31738 22094 31790
rect 22146 31738 22148 31790
rect 22092 31726 22148 31738
rect 22204 31668 22260 32284
rect 22092 31612 22260 31668
rect 22092 30996 22148 31612
rect 22316 31554 22372 31566
rect 22316 31502 22318 31554
rect 22370 31502 22372 31554
rect 22204 30996 22260 31006
rect 22092 30994 22260 30996
rect 22092 30942 22206 30994
rect 22258 30942 22260 30994
rect 22092 30940 22260 30942
rect 22204 30930 22260 30940
rect 21420 30046 21422 30098
rect 21474 30046 21476 30098
rect 21420 30034 21476 30046
rect 21868 30828 22036 30884
rect 21756 29988 21812 29998
rect 21196 29764 21252 29774
rect 21196 29650 21252 29708
rect 21196 29598 21198 29650
rect 21250 29598 21252 29650
rect 21196 29586 21252 29598
rect 21308 28532 21364 28542
rect 21308 28438 21364 28476
rect 21420 28420 21476 28430
rect 21644 28420 21700 28430
rect 21420 28326 21476 28364
rect 21532 28418 21700 28420
rect 21532 28366 21646 28418
rect 21698 28366 21700 28418
rect 21532 28364 21700 28366
rect 21084 28252 21364 28308
rect 21084 28082 21140 28094
rect 21084 28030 21086 28082
rect 21138 28030 21140 28082
rect 20860 27806 20862 27858
rect 20914 27806 20916 27858
rect 20860 27794 20916 27806
rect 20972 27970 21028 27982
rect 20972 27918 20974 27970
rect 21026 27918 21028 27970
rect 20972 26516 21028 27918
rect 20860 26292 20916 26302
rect 20748 26290 20916 26292
rect 20748 26238 20862 26290
rect 20914 26238 20916 26290
rect 20748 26236 20916 26238
rect 20860 26226 20916 26236
rect 20972 26068 21028 26460
rect 20972 26002 21028 26012
rect 20524 25508 20580 25518
rect 20524 25506 20692 25508
rect 20524 25454 20526 25506
rect 20578 25454 20692 25506
rect 20524 25452 20692 25454
rect 20524 25442 20580 25452
rect 20188 24994 20244 25004
rect 20412 25394 20468 25406
rect 20412 25342 20414 25394
rect 20466 25342 20468 25394
rect 19740 24948 19796 24958
rect 19740 24834 19796 24892
rect 20412 24948 20468 25342
rect 20412 24882 20468 24892
rect 19740 24782 19742 24834
rect 19794 24782 19796 24834
rect 19292 23826 19348 23838
rect 19292 23774 19294 23826
rect 19346 23774 19348 23826
rect 19292 23716 19348 23774
rect 19292 23650 19348 23660
rect 19292 22482 19348 22494
rect 19292 22430 19294 22482
rect 19346 22430 19348 22482
rect 19292 22148 19348 22430
rect 19292 22082 19348 22092
rect 19404 21586 19460 23884
rect 19516 24722 19572 24734
rect 19516 24670 19518 24722
rect 19570 24670 19572 24722
rect 19516 21812 19572 24670
rect 19516 21746 19572 21756
rect 19628 23938 19684 23950
rect 19628 23886 19630 23938
rect 19682 23886 19684 23938
rect 19404 21534 19406 21586
rect 19458 21534 19460 21586
rect 19404 21522 19460 21534
rect 19628 20916 19684 23886
rect 19740 23716 19796 24782
rect 20188 24836 20244 24846
rect 20188 24742 20244 24780
rect 20524 24722 20580 24734
rect 20524 24670 20526 24722
rect 20578 24670 20580 24722
rect 20188 23940 20244 23950
rect 20524 23940 20580 24670
rect 20244 23884 20580 23940
rect 20188 23846 20244 23884
rect 19740 23650 19796 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20300 23268 20356 23278
rect 20300 23044 20356 23212
rect 20188 23042 20356 23044
rect 20188 22990 20302 23042
rect 20354 22990 20356 23042
rect 20188 22988 20356 22990
rect 19964 22372 20020 22382
rect 19964 22278 20020 22316
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19964 21812 20020 21822
rect 20188 21812 20244 22988
rect 20300 22978 20356 22988
rect 20524 22484 20580 22494
rect 20524 22390 20580 22428
rect 20636 22372 20692 25452
rect 21084 25396 21140 28030
rect 21308 28084 21364 28252
rect 21308 28028 21476 28084
rect 21308 27860 21364 27870
rect 21308 26628 21364 27804
rect 21420 26962 21476 28028
rect 21532 27636 21588 28364
rect 21644 28354 21700 28364
rect 21756 28196 21812 29932
rect 21644 28140 21812 28196
rect 21644 27860 21700 28140
rect 21868 27970 21924 30828
rect 21980 30660 22036 30670
rect 21980 29314 22036 30604
rect 22092 30212 22148 30222
rect 22092 30118 22148 30156
rect 21980 29262 21982 29314
rect 22034 29262 22036 29314
rect 21980 29092 22036 29262
rect 22316 29316 22372 31502
rect 22428 31218 22484 31230
rect 22428 31166 22430 31218
rect 22482 31166 22484 31218
rect 22428 30660 22484 31166
rect 22540 31220 22596 32622
rect 22652 31780 22708 33628
rect 22764 33124 22820 33134
rect 22764 33030 22820 33068
rect 22764 31780 22820 31790
rect 22652 31778 22820 31780
rect 22652 31726 22766 31778
rect 22818 31726 22820 31778
rect 22652 31724 22820 31726
rect 22764 31714 22820 31724
rect 22540 31154 22596 31164
rect 22540 30996 22596 31006
rect 22540 30994 23156 30996
rect 22540 30942 22542 30994
rect 22594 30942 23156 30994
rect 22540 30940 23156 30942
rect 22540 30930 22596 30940
rect 22428 30594 22484 30604
rect 22540 30210 22596 30222
rect 22540 30158 22542 30210
rect 22594 30158 22596 30210
rect 22540 29988 22596 30158
rect 22540 29922 22596 29932
rect 23100 30098 23156 30940
rect 23100 30046 23102 30098
rect 23154 30046 23156 30098
rect 23100 29876 23156 30046
rect 23100 29810 23156 29820
rect 23212 29540 23268 33852
rect 23324 33124 23380 33134
rect 23324 31778 23380 33068
rect 23324 31726 23326 31778
rect 23378 31726 23380 31778
rect 23324 31714 23380 31726
rect 23436 31780 23492 31790
rect 22876 29484 23268 29540
rect 23436 30994 23492 31724
rect 23436 30942 23438 30994
rect 23490 30942 23492 30994
rect 23436 30210 23492 30942
rect 23436 30158 23438 30210
rect 23490 30158 23492 30210
rect 22316 29250 22372 29260
rect 22652 29428 22708 29438
rect 21980 29026 22036 29036
rect 22652 28754 22708 29372
rect 22652 28702 22654 28754
rect 22706 28702 22708 28754
rect 22204 28644 22260 28654
rect 21868 27918 21870 27970
rect 21922 27918 21924 27970
rect 21868 27906 21924 27918
rect 21980 28642 22260 28644
rect 21980 28590 22206 28642
rect 22258 28590 22260 28642
rect 21980 28588 22260 28590
rect 21644 27794 21700 27804
rect 21756 27858 21812 27870
rect 21756 27806 21758 27858
rect 21810 27806 21812 27858
rect 21532 27580 21700 27636
rect 21532 27412 21588 27422
rect 21532 27074 21588 27356
rect 21532 27022 21534 27074
rect 21586 27022 21588 27074
rect 21532 27010 21588 27022
rect 21420 26910 21422 26962
rect 21474 26910 21476 26962
rect 21420 26898 21476 26910
rect 21308 26572 21476 26628
rect 21308 26402 21364 26414
rect 21308 26350 21310 26402
rect 21362 26350 21364 26402
rect 21308 26068 21364 26350
rect 21308 26002 21364 26012
rect 20860 25340 21140 25396
rect 21308 25506 21364 25518
rect 21308 25454 21310 25506
rect 21362 25454 21364 25506
rect 21308 25396 21364 25454
rect 20748 23940 20804 23950
rect 20860 23940 20916 25340
rect 21308 25330 21364 25340
rect 21196 25284 21252 25294
rect 20972 25282 21252 25284
rect 20972 25230 21198 25282
rect 21250 25230 21252 25282
rect 20972 25228 21252 25230
rect 20972 24722 21028 25228
rect 21196 25218 21252 25228
rect 20972 24670 20974 24722
rect 21026 24670 21028 24722
rect 20972 24658 21028 24670
rect 21308 24276 21364 24286
rect 20748 23938 20916 23940
rect 20748 23886 20750 23938
rect 20802 23886 20916 23938
rect 20748 23884 20916 23886
rect 21196 24220 21308 24276
rect 20748 23874 20804 23884
rect 20748 23380 20804 23390
rect 20748 23286 20804 23324
rect 21196 23154 21252 24220
rect 21308 24210 21364 24220
rect 21420 23940 21476 26572
rect 21644 25956 21700 27580
rect 21756 27300 21812 27806
rect 21756 26292 21812 27244
rect 21980 27860 22036 28588
rect 22204 28578 22260 28588
rect 22316 28644 22372 28654
rect 22092 28420 22148 28430
rect 22316 28420 22372 28588
rect 22148 28364 22372 28420
rect 22092 28326 22148 28364
rect 21980 26852 22036 27804
rect 22204 27636 22260 27646
rect 22092 27188 22148 27198
rect 22092 26962 22148 27132
rect 22204 27074 22260 27580
rect 22204 27022 22206 27074
rect 22258 27022 22260 27074
rect 22204 27010 22260 27022
rect 22428 27076 22484 27086
rect 22092 26910 22094 26962
rect 22146 26910 22148 26962
rect 22092 26898 22148 26910
rect 21980 26786 22036 26796
rect 22204 26850 22260 26862
rect 22204 26798 22206 26850
rect 22258 26798 22260 26850
rect 21980 26404 22036 26414
rect 21980 26310 22036 26348
rect 21756 26198 21812 26236
rect 21644 25890 21700 25900
rect 21196 23102 21198 23154
rect 21250 23102 21252 23154
rect 21196 23090 21252 23102
rect 21308 23884 21476 23940
rect 21644 25508 21700 25518
rect 21308 22596 21364 23884
rect 21420 23716 21476 23726
rect 21420 23714 21588 23716
rect 21420 23662 21422 23714
rect 21474 23662 21588 23714
rect 21420 23660 21588 23662
rect 21420 23650 21476 23660
rect 21420 23156 21476 23166
rect 21420 22708 21476 23100
rect 21532 23042 21588 23660
rect 21532 22990 21534 23042
rect 21586 22990 21588 23042
rect 21532 22978 21588 22990
rect 21420 22642 21476 22652
rect 20636 22306 20692 22316
rect 21084 22540 21364 22596
rect 19964 21810 20244 21812
rect 19964 21758 19966 21810
rect 20018 21758 20244 21810
rect 19964 21756 20244 21758
rect 20412 21812 20468 21822
rect 20636 21812 20692 21822
rect 19964 21746 20020 21756
rect 20412 21718 20468 21756
rect 20524 21756 20636 21812
rect 20524 21698 20580 21756
rect 20636 21746 20692 21756
rect 20524 21646 20526 21698
rect 20578 21646 20580 21698
rect 20300 21586 20356 21598
rect 20300 21534 20302 21586
rect 20354 21534 20356 21586
rect 20300 21140 20356 21534
rect 20300 21074 20356 21084
rect 19628 20850 19684 20860
rect 20300 20916 20356 20926
rect 20300 20822 20356 20860
rect 20412 20804 20468 20814
rect 20524 20804 20580 21646
rect 20972 21700 21028 21710
rect 20972 21586 21028 21644
rect 20972 21534 20974 21586
rect 21026 21534 21028 21586
rect 20972 21522 21028 21534
rect 20412 20802 20580 20804
rect 20412 20750 20414 20802
rect 20466 20750 20580 20802
rect 20412 20748 20580 20750
rect 20860 21252 20916 21262
rect 20860 20802 20916 21196
rect 20860 20750 20862 20802
rect 20914 20750 20916 20802
rect 20412 20738 20468 20748
rect 20860 20738 20916 20750
rect 20188 20578 20244 20590
rect 20188 20526 20190 20578
rect 20242 20526 20244 20578
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20076 20132 20132 20142
rect 19852 20018 19908 20030
rect 19852 19966 19854 20018
rect 19906 19966 19908 20018
rect 19628 19908 19684 19918
rect 19852 19908 19908 19966
rect 19628 19906 19908 19908
rect 19628 19854 19630 19906
rect 19682 19854 19908 19906
rect 19628 19852 19908 19854
rect 19628 19572 19684 19852
rect 19628 19506 19684 19516
rect 20076 19346 20132 20076
rect 20076 19294 20078 19346
rect 20130 19294 20132 19346
rect 20076 19282 20132 19294
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19740 18564 19796 18574
rect 19180 18450 19236 18462
rect 19740 18452 19796 18508
rect 19180 18398 19182 18450
rect 19234 18398 19236 18450
rect 19180 16772 19236 18398
rect 19628 18450 19796 18452
rect 19628 18398 19742 18450
rect 19794 18398 19796 18450
rect 19628 18396 19796 18398
rect 19180 16706 19236 16716
rect 19292 18340 19348 18350
rect 19068 16482 19124 16492
rect 19292 14530 19348 18284
rect 19516 17666 19572 17678
rect 19516 17614 19518 17666
rect 19570 17614 19572 17666
rect 19404 17556 19460 17566
rect 19404 16324 19460 17500
rect 19516 16884 19572 17614
rect 19628 16994 19684 18396
rect 19740 18386 19796 18396
rect 20188 17892 20244 20526
rect 21084 20132 21140 22540
rect 21420 22372 21476 22382
rect 21420 22278 21476 22316
rect 21308 22148 21364 22158
rect 21084 20066 21140 20076
rect 21196 22146 21364 22148
rect 21196 22094 21310 22146
rect 21362 22094 21364 22146
rect 21196 22092 21364 22094
rect 20300 19796 20356 19806
rect 20300 19794 20468 19796
rect 20300 19742 20302 19794
rect 20354 19742 20468 19794
rect 20300 19740 20468 19742
rect 20300 19730 20356 19740
rect 20412 17892 20468 19740
rect 21196 18676 21252 22092
rect 21308 22082 21364 22092
rect 21532 22146 21588 22158
rect 21532 22094 21534 22146
rect 21586 22094 21588 22146
rect 21532 21812 21588 22094
rect 21532 21746 21588 21756
rect 21644 21588 21700 25452
rect 21868 24722 21924 24734
rect 21868 24670 21870 24722
rect 21922 24670 21924 24722
rect 21756 23268 21812 23278
rect 21868 23268 21924 24670
rect 22204 24610 22260 26798
rect 22428 26402 22484 27020
rect 22428 26350 22430 26402
rect 22482 26350 22484 26402
rect 22428 26338 22484 26350
rect 22540 26290 22596 26302
rect 22540 26238 22542 26290
rect 22594 26238 22596 26290
rect 22428 26068 22484 26078
rect 22316 25508 22372 25518
rect 22316 25414 22372 25452
rect 22428 25394 22484 26012
rect 22540 25956 22596 26238
rect 22652 26292 22708 28702
rect 22876 27746 22932 29484
rect 23324 29426 23380 29438
rect 23324 29374 23326 29426
rect 23378 29374 23380 29426
rect 22876 27694 22878 27746
rect 22930 27694 22932 27746
rect 22876 27682 22932 27694
rect 22988 29314 23044 29326
rect 22988 29262 22990 29314
rect 23042 29262 23044 29314
rect 22988 29204 23044 29262
rect 22988 26908 23044 29148
rect 23100 29316 23156 29326
rect 23100 28530 23156 29260
rect 23324 29204 23380 29374
rect 23436 29428 23492 30158
rect 23436 29362 23492 29372
rect 23436 29204 23492 29214
rect 23324 29148 23436 29204
rect 23436 29138 23492 29148
rect 23100 28478 23102 28530
rect 23154 28478 23156 28530
rect 23100 28466 23156 28478
rect 23324 28644 23380 28654
rect 23212 28418 23268 28430
rect 23212 28366 23214 28418
rect 23266 28366 23268 28418
rect 23212 28084 23268 28366
rect 23212 28018 23268 28028
rect 23324 28082 23380 28588
rect 23436 28420 23492 28430
rect 23436 28326 23492 28364
rect 23324 28030 23326 28082
rect 23378 28030 23380 28082
rect 23324 28018 23380 28030
rect 23100 27076 23156 27086
rect 23100 26982 23156 27020
rect 23548 26964 23604 35756
rect 23772 34914 23828 37884
rect 23884 37874 23940 37884
rect 23996 37940 24052 37950
rect 23996 37268 24052 37884
rect 23996 37174 24052 37212
rect 24108 36708 24164 38108
rect 24220 37828 24276 37838
rect 24220 37734 24276 37772
rect 24556 37828 24612 37838
rect 24556 37734 24612 37772
rect 24892 37826 24948 37838
rect 24892 37774 24894 37826
rect 24946 37774 24948 37826
rect 24444 37378 24500 37390
rect 24444 37326 24446 37378
rect 24498 37326 24500 37378
rect 24444 37156 24500 37326
rect 24444 37090 24500 37100
rect 24556 37266 24612 37278
rect 24556 37214 24558 37266
rect 24610 37214 24612 37266
rect 24108 36642 24164 36652
rect 24332 37042 24388 37054
rect 24332 36990 24334 37042
rect 24386 36990 24388 37042
rect 24332 35698 24388 36990
rect 24556 37044 24612 37214
rect 24556 36978 24612 36988
rect 24892 36484 24948 37774
rect 25228 37828 25284 37838
rect 25228 37734 25284 37772
rect 25452 37268 25508 37278
rect 25340 37156 25396 37166
rect 24892 36418 24948 36428
rect 25116 37100 25340 37156
rect 25116 36482 25172 37100
rect 25340 37062 25396 37100
rect 25116 36430 25118 36482
rect 25170 36430 25172 36482
rect 25116 36418 25172 36430
rect 25452 36482 25508 37212
rect 25452 36430 25454 36482
rect 25506 36430 25508 36482
rect 25452 36418 25508 36430
rect 25676 36596 25732 38612
rect 26236 38276 26292 38286
rect 25900 37940 25956 37950
rect 25788 37492 25844 37502
rect 25788 37398 25844 37436
rect 24332 35646 24334 35698
rect 24386 35646 24388 35698
rect 24332 35634 24388 35646
rect 24892 36258 24948 36270
rect 24892 36206 24894 36258
rect 24946 36206 24948 36258
rect 23772 34862 23774 34914
rect 23826 34862 23828 34914
rect 23772 34850 23828 34862
rect 24332 35476 24388 35486
rect 24332 34914 24388 35420
rect 24332 34862 24334 34914
rect 24386 34862 24388 34914
rect 24332 34850 24388 34862
rect 24892 34914 24948 36206
rect 25564 35476 25620 35486
rect 25564 35382 25620 35420
rect 24892 34862 24894 34914
rect 24946 34862 24948 34914
rect 24892 34850 24948 34862
rect 23772 34692 23828 34702
rect 23772 34356 23828 34636
rect 23884 34692 23940 34702
rect 23884 34690 24052 34692
rect 23884 34638 23886 34690
rect 23938 34638 24052 34690
rect 23884 34636 24052 34638
rect 23884 34626 23940 34636
rect 23884 34356 23940 34366
rect 23772 34354 23940 34356
rect 23772 34302 23886 34354
rect 23938 34302 23940 34354
rect 23772 34300 23940 34302
rect 23884 34290 23940 34300
rect 23660 34244 23716 34254
rect 23660 29650 23716 34188
rect 23996 33460 24052 34636
rect 25564 34356 25620 34366
rect 25676 34356 25732 36540
rect 25900 35698 25956 37884
rect 26124 37716 26180 37726
rect 26124 37266 26180 37660
rect 26124 37214 26126 37266
rect 26178 37214 26180 37266
rect 26124 37202 26180 37214
rect 25900 35646 25902 35698
rect 25954 35646 25956 35698
rect 25900 35634 25956 35646
rect 26124 37042 26180 37054
rect 26124 36990 26126 37042
rect 26178 36990 26180 37042
rect 26012 34916 26068 34926
rect 26124 34916 26180 36990
rect 26236 35700 26292 38220
rect 26348 36932 26404 41134
rect 26684 40516 26740 42590
rect 26908 42084 26964 42094
rect 26908 41186 26964 42028
rect 27244 41412 27300 43262
rect 27916 42644 27972 42654
rect 27916 42642 28084 42644
rect 27916 42590 27918 42642
rect 27970 42590 28084 42642
rect 27916 42588 28084 42590
rect 27916 42578 27972 42588
rect 28028 42532 28084 42588
rect 28028 42466 28084 42476
rect 28140 42530 28196 42542
rect 28140 42478 28142 42530
rect 28194 42478 28196 42530
rect 27244 41346 27300 41356
rect 26908 41134 26910 41186
rect 26962 41134 26964 41186
rect 26908 41122 26964 41134
rect 27132 41188 27188 41198
rect 26796 40516 26852 40526
rect 26684 40514 26852 40516
rect 26684 40462 26798 40514
rect 26850 40462 26852 40514
rect 26684 40460 26852 40462
rect 26796 40450 26852 40460
rect 27132 40516 27188 41132
rect 27132 40402 27188 40460
rect 27132 40350 27134 40402
rect 27186 40350 27188 40402
rect 27132 40338 27188 40350
rect 27580 41074 27636 41086
rect 27580 41022 27582 41074
rect 27634 41022 27636 41074
rect 27580 40402 27636 41022
rect 27916 40964 27972 40974
rect 27580 40350 27582 40402
rect 27634 40350 27636 40402
rect 27580 40338 27636 40350
rect 27692 40962 27972 40964
rect 27692 40910 27918 40962
rect 27970 40910 27972 40962
rect 27692 40908 27972 40910
rect 27692 40180 27748 40908
rect 27916 40898 27972 40908
rect 27580 40124 27748 40180
rect 27804 40514 27860 40526
rect 27804 40462 27806 40514
rect 27858 40462 27860 40514
rect 27356 39732 27412 39742
rect 26572 37828 26628 37838
rect 26460 37268 26516 37278
rect 26460 37174 26516 37212
rect 26348 36866 26404 36876
rect 26572 36372 26628 37772
rect 26460 36370 26628 36372
rect 26460 36318 26574 36370
rect 26626 36318 26628 36370
rect 26460 36316 26628 36318
rect 26348 35700 26404 35710
rect 26236 35698 26404 35700
rect 26236 35646 26350 35698
rect 26402 35646 26404 35698
rect 26236 35644 26404 35646
rect 26012 34914 26180 34916
rect 26012 34862 26014 34914
rect 26066 34862 26180 34914
rect 26012 34860 26180 34862
rect 26348 35028 26404 35644
rect 26012 34850 26068 34860
rect 25564 34354 25732 34356
rect 25564 34302 25566 34354
rect 25618 34302 25732 34354
rect 25564 34300 25732 34302
rect 25564 34290 25620 34300
rect 25228 34244 25284 34254
rect 25228 34150 25284 34188
rect 24444 34018 24500 34030
rect 24444 33966 24446 34018
rect 24498 33966 24500 34018
rect 24444 33684 24500 33966
rect 26348 33908 26404 34972
rect 26460 34242 26516 36316
rect 26572 36306 26628 36316
rect 27132 37156 27188 37166
rect 26684 36260 26740 36270
rect 26684 35810 26740 36204
rect 26684 35758 26686 35810
rect 26738 35758 26740 35810
rect 26684 35746 26740 35758
rect 27132 35698 27188 37100
rect 27356 35924 27412 39676
rect 27580 39620 27636 40124
rect 27580 38946 27636 39564
rect 27692 39508 27748 39518
rect 27692 39414 27748 39452
rect 27580 38894 27582 38946
rect 27634 38894 27636 38946
rect 27580 38882 27636 38894
rect 27804 37940 27860 40462
rect 28028 39620 28084 39630
rect 28140 39620 28196 42478
rect 28028 39618 28196 39620
rect 28028 39566 28030 39618
rect 28082 39566 28196 39618
rect 28028 39564 28196 39566
rect 28252 40962 28308 43598
rect 28364 42756 28420 43710
rect 30492 43650 30548 43662
rect 30492 43598 30494 43650
rect 30546 43598 30548 43650
rect 29484 43540 29540 43550
rect 29484 43446 29540 43484
rect 30492 43540 30548 43598
rect 28364 42690 28420 42700
rect 28700 43426 28756 43438
rect 28700 43374 28702 43426
rect 28754 43374 28756 43426
rect 28476 42642 28532 42654
rect 28476 42590 28478 42642
rect 28530 42590 28532 42642
rect 28252 40910 28254 40962
rect 28306 40910 28308 40962
rect 28252 40628 28308 40910
rect 28028 39284 28084 39564
rect 28252 39506 28308 40572
rect 28252 39454 28254 39506
rect 28306 39454 28308 39506
rect 28252 39442 28308 39454
rect 28364 42532 28420 42542
rect 28476 42532 28532 42590
rect 28420 42476 28532 42532
rect 28028 39218 28084 39228
rect 27804 37874 27860 37884
rect 28364 37378 28420 42476
rect 28700 41972 28756 43374
rect 30268 43314 30324 43326
rect 30268 43262 30270 43314
rect 30322 43262 30324 43314
rect 29260 42756 29316 42766
rect 29260 42754 29428 42756
rect 29260 42702 29262 42754
rect 29314 42702 29428 42754
rect 29260 42700 29428 42702
rect 29260 42690 29316 42700
rect 28700 41906 28756 41916
rect 28924 41858 28980 41870
rect 28924 41806 28926 41858
rect 28978 41806 28980 41858
rect 28476 41076 28532 41086
rect 28476 40404 28532 41020
rect 28476 40310 28532 40348
rect 28924 40402 28980 41806
rect 29148 41076 29204 41086
rect 29148 41074 29316 41076
rect 29148 41022 29150 41074
rect 29202 41022 29316 41074
rect 29148 41020 29316 41022
rect 29148 41010 29204 41020
rect 28924 40350 28926 40402
rect 28978 40350 28980 40402
rect 28924 40338 28980 40350
rect 29148 39396 29204 39406
rect 29148 39302 29204 39340
rect 29260 39060 29316 41020
rect 29372 40404 29428 42700
rect 30268 42084 30324 43262
rect 30492 43092 30548 43484
rect 30828 43540 30884 43550
rect 30828 43538 31220 43540
rect 30828 43486 30830 43538
rect 30882 43486 31220 43538
rect 30828 43484 31220 43486
rect 30828 43474 30884 43484
rect 30492 43036 30772 43092
rect 30156 42028 30324 42084
rect 30492 42756 30548 42766
rect 30044 41972 30100 41982
rect 30044 41878 30100 41916
rect 29484 41188 29540 41198
rect 29484 41094 29540 41132
rect 29932 41188 29988 41198
rect 30156 41188 30212 42028
rect 29932 41094 29988 41132
rect 30044 41132 30212 41188
rect 29708 40404 29764 40414
rect 29372 40348 29708 40404
rect 29708 39620 29764 40348
rect 29932 40404 29988 40414
rect 30044 40404 30100 41132
rect 30156 40964 30212 40974
rect 30156 40870 30212 40908
rect 30380 40516 30436 40526
rect 30492 40516 30548 42700
rect 30604 41970 30660 41982
rect 30604 41918 30606 41970
rect 30658 41918 30660 41970
rect 30604 41300 30660 41918
rect 30716 41972 30772 43036
rect 30828 41972 30884 41982
rect 30716 41970 30884 41972
rect 30716 41918 30830 41970
rect 30882 41918 30884 41970
rect 30716 41916 30884 41918
rect 30828 41906 30884 41916
rect 30604 41244 30772 41300
rect 30604 41076 30660 41086
rect 30604 40982 30660 41020
rect 29932 40402 30100 40404
rect 29932 40350 29934 40402
rect 29986 40350 30100 40402
rect 29932 40348 30100 40350
rect 30156 40514 30492 40516
rect 30156 40462 30382 40514
rect 30434 40462 30492 40514
rect 30156 40460 30492 40462
rect 29932 40338 29988 40348
rect 30156 39956 30212 40460
rect 30380 40450 30436 40460
rect 30492 40422 30548 40460
rect 29708 39554 29764 39564
rect 29820 39900 30212 39956
rect 29820 39618 29876 39900
rect 29820 39566 29822 39618
rect 29874 39566 29876 39618
rect 29820 39554 29876 39566
rect 30044 39620 30100 39630
rect 30044 39526 30100 39564
rect 29372 39508 29428 39518
rect 29372 39414 29428 39452
rect 29372 39060 29428 39070
rect 29260 39058 29428 39060
rect 29260 39006 29374 39058
rect 29426 39006 29428 39058
rect 29260 39004 29428 39006
rect 29372 38994 29428 39004
rect 30716 38948 30772 41244
rect 30716 38882 30772 38892
rect 30828 40402 30884 40414
rect 30828 40350 30830 40402
rect 30882 40350 30884 40402
rect 30044 38724 30100 38734
rect 28364 37326 28366 37378
rect 28418 37326 28420 37378
rect 27132 35646 27134 35698
rect 27186 35646 27188 35698
rect 27020 35476 27076 35486
rect 26572 35028 26628 35038
rect 26572 34934 26628 34972
rect 26460 34190 26462 34242
rect 26514 34190 26516 34242
rect 26460 34178 26516 34190
rect 26348 33842 26404 33852
rect 24444 33618 24500 33628
rect 25564 33572 25620 33582
rect 24668 33460 24724 33470
rect 23996 33394 24052 33404
rect 24444 33458 24724 33460
rect 24444 33406 24670 33458
rect 24722 33406 24724 33458
rect 24444 33404 24724 33406
rect 24220 33124 24276 33134
rect 23884 33122 24276 33124
rect 23884 33070 24222 33122
rect 24274 33070 24276 33122
rect 23884 33068 24276 33070
rect 23884 29764 23940 33068
rect 24220 33058 24276 33068
rect 24332 32564 24388 32574
rect 24444 32564 24500 33404
rect 24668 33394 24724 33404
rect 25228 33348 25284 33358
rect 25228 33254 25284 33292
rect 24556 33124 24612 33134
rect 24556 32674 24612 33068
rect 25452 33124 25508 33134
rect 25452 33030 25508 33068
rect 24556 32622 24558 32674
rect 24610 32622 24612 32674
rect 24556 32610 24612 32622
rect 24332 32562 24444 32564
rect 24332 32510 24334 32562
rect 24386 32510 24444 32562
rect 24332 32508 24444 32510
rect 24332 32498 24388 32508
rect 24108 32338 24164 32350
rect 24108 32286 24110 32338
rect 24162 32286 24164 32338
rect 24108 31780 24164 32286
rect 24332 31780 24388 31790
rect 24108 31778 24388 31780
rect 24108 31726 24334 31778
rect 24386 31726 24388 31778
rect 24108 31724 24388 31726
rect 24332 31714 24388 31724
rect 23884 29698 23940 29708
rect 24108 31220 24164 31230
rect 23660 29598 23662 29650
rect 23714 29598 23716 29650
rect 23660 29540 23716 29598
rect 24108 29650 24164 31164
rect 24332 30884 24388 30894
rect 24332 30210 24388 30828
rect 24332 30158 24334 30210
rect 24386 30158 24388 30210
rect 24332 30146 24388 30158
rect 24108 29598 24110 29650
rect 24162 29598 24164 29650
rect 24108 29586 24164 29598
rect 24332 29876 24388 29886
rect 23660 29474 23716 29484
rect 23884 28644 23940 28654
rect 23660 28420 23716 28430
rect 23660 28418 23828 28420
rect 23660 28366 23662 28418
rect 23714 28366 23828 28418
rect 23660 28364 23828 28366
rect 23660 28354 23716 28364
rect 23660 27860 23716 27870
rect 23660 27766 23716 27804
rect 23772 26908 23828 28364
rect 22988 26852 23268 26908
rect 23548 26898 23604 26908
rect 22988 26292 23044 26302
rect 22652 26290 23044 26292
rect 22652 26238 22990 26290
rect 23042 26238 23044 26290
rect 22652 26236 23044 26238
rect 22540 25890 22596 25900
rect 22428 25342 22430 25394
rect 22482 25342 22484 25394
rect 22428 25330 22484 25342
rect 22652 25396 22708 25406
rect 22540 24724 22596 24734
rect 22428 24722 22596 24724
rect 22428 24670 22542 24722
rect 22594 24670 22596 24722
rect 22428 24668 22596 24670
rect 22204 24558 22206 24610
rect 22258 24558 22260 24610
rect 22204 24546 22260 24558
rect 22316 24612 22372 24622
rect 22316 24518 22372 24556
rect 21980 23940 22036 23950
rect 21980 23938 22260 23940
rect 21980 23886 21982 23938
rect 22034 23886 22260 23938
rect 21980 23884 22260 23886
rect 21980 23874 22036 23884
rect 21812 23212 21924 23268
rect 21756 23202 21812 23212
rect 22204 23156 22260 23884
rect 22204 23090 22260 23100
rect 22428 22484 22484 24668
rect 22540 24658 22596 24668
rect 22652 23938 22708 25340
rect 22652 23886 22654 23938
rect 22706 23886 22708 23938
rect 22652 23874 22708 23886
rect 22764 25060 22820 25070
rect 22764 23716 22820 25004
rect 22652 23660 22764 23716
rect 21980 22428 22484 22484
rect 22540 23154 22596 23166
rect 22540 23102 22542 23154
rect 22594 23102 22596 23154
rect 21868 22372 21924 22382
rect 21868 22278 21924 22316
rect 21980 21810 22036 22428
rect 21980 21758 21982 21810
rect 22034 21758 22036 21810
rect 21980 21746 22036 21758
rect 22092 21812 22148 21822
rect 21196 18610 21252 18620
rect 21420 21532 21700 21588
rect 21868 21586 21924 21598
rect 21868 21534 21870 21586
rect 21922 21534 21924 21586
rect 20524 18450 20580 18462
rect 21420 18452 21476 21532
rect 21756 19348 21812 19358
rect 21756 19254 21812 19292
rect 21644 19012 21700 19022
rect 20524 18398 20526 18450
rect 20578 18398 20580 18450
rect 20524 18340 20580 18398
rect 20524 18274 20580 18284
rect 21084 18396 21476 18452
rect 21532 19010 21700 19012
rect 21532 18958 21646 19010
rect 21698 18958 21700 19010
rect 21532 18956 21700 18958
rect 20188 17836 20356 17892
rect 19852 17780 19908 17790
rect 19852 17778 20244 17780
rect 19852 17726 19854 17778
rect 19906 17726 20244 17778
rect 19852 17724 20244 17726
rect 19852 17714 19908 17724
rect 20076 17556 20132 17566
rect 20076 17462 20132 17500
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 16942 19630 16994
rect 19682 16942 19684 16994
rect 19628 16930 19684 16942
rect 19516 16818 19572 16828
rect 19404 16258 19460 16268
rect 19516 16548 19572 16558
rect 19516 15988 19572 16492
rect 20188 16322 20244 17724
rect 20300 17444 20356 17836
rect 20412 17826 20468 17836
rect 20412 17668 20468 17678
rect 20412 17666 20580 17668
rect 20412 17614 20414 17666
rect 20466 17614 20580 17666
rect 20412 17612 20580 17614
rect 20412 17602 20468 17612
rect 20300 17388 20468 17444
rect 20188 16270 20190 16322
rect 20242 16270 20244 16322
rect 20188 16258 20244 16270
rect 20300 17220 20356 17230
rect 19740 16100 19796 16110
rect 19964 16100 20020 16110
rect 19740 16098 20020 16100
rect 19740 16046 19742 16098
rect 19794 16046 19966 16098
rect 20018 16046 20020 16098
rect 19740 16044 20020 16046
rect 19740 16034 19796 16044
rect 19964 16034 20020 16044
rect 20300 16098 20356 17164
rect 20300 16046 20302 16098
rect 20354 16046 20356 16098
rect 20300 16034 20356 16046
rect 19516 15426 19572 15932
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20300 15540 20356 15550
rect 20300 15446 20356 15484
rect 19516 15374 19518 15426
rect 19570 15374 19572 15426
rect 19516 15362 19572 15374
rect 19292 14478 19294 14530
rect 19346 14478 19348 14530
rect 19292 14466 19348 14478
rect 19628 15204 19684 15214
rect 18732 13878 18788 13916
rect 18284 13746 18340 13758
rect 18284 13694 18286 13746
rect 18338 13694 18340 13746
rect 18284 13412 18340 13694
rect 18284 13346 18340 13356
rect 19628 13746 19684 15148
rect 19964 14980 20020 14990
rect 19740 14530 19796 14542
rect 19740 14478 19742 14530
rect 19794 14478 19796 14530
rect 19740 14308 19796 14478
rect 19740 14242 19796 14252
rect 19964 14306 20020 14924
rect 19964 14254 19966 14306
rect 20018 14254 20020 14306
rect 19964 14242 20020 14254
rect 20188 14308 20244 14318
rect 20300 14308 20356 14318
rect 20244 14306 20356 14308
rect 20244 14254 20302 14306
rect 20354 14254 20356 14306
rect 20244 14252 20356 14254
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13694 19630 13746
rect 19682 13694 19684 13746
rect 19628 13076 19684 13694
rect 18172 13022 18174 13074
rect 18226 13022 18228 13074
rect 18172 12964 18228 13022
rect 17836 12178 17892 12908
rect 18172 12898 18228 12908
rect 19068 13020 19684 13076
rect 19068 12962 19124 13020
rect 19068 12910 19070 12962
rect 19122 12910 19124 12962
rect 19068 12898 19124 12910
rect 18508 12850 18564 12862
rect 19404 12852 19460 12862
rect 18508 12798 18510 12850
rect 18562 12798 18564 12850
rect 17948 12740 18004 12750
rect 18004 12684 18116 12740
rect 17948 12674 18004 12684
rect 17836 12126 17838 12178
rect 17890 12126 17892 12178
rect 17500 11230 17502 11282
rect 17554 11230 17556 11282
rect 16716 10770 16772 10780
rect 16044 10612 16100 10622
rect 16044 10518 16100 10556
rect 17388 10612 17444 10622
rect 17388 10518 17444 10556
rect 16604 10498 16660 10510
rect 16604 10446 16606 10498
rect 16658 10446 16660 10498
rect 16604 10052 16660 10446
rect 16604 9986 16660 9996
rect 17276 10052 17332 10062
rect 15596 9154 15876 9156
rect 15596 9102 15598 9154
rect 15650 9102 15876 9154
rect 15596 9100 15876 9102
rect 15932 9826 15988 9838
rect 15932 9774 15934 9826
rect 15986 9774 15988 9826
rect 15596 9090 15652 9100
rect 15820 8372 15876 8382
rect 15932 8372 15988 9774
rect 16828 9826 16884 9838
rect 16828 9774 16830 9826
rect 16882 9774 16884 9826
rect 15820 8370 15988 8372
rect 15820 8318 15822 8370
rect 15874 8318 15988 8370
rect 15820 8316 15988 8318
rect 16044 9716 16100 9726
rect 15820 8306 15876 8316
rect 15484 8194 15540 8204
rect 15484 6692 15540 6702
rect 15372 6690 15652 6692
rect 15372 6638 15486 6690
rect 15538 6638 15652 6690
rect 15372 6636 15652 6638
rect 15484 6626 15540 6636
rect 5852 6078 5854 6130
rect 5906 6078 5908 6130
rect 5852 6066 5908 6078
rect 2716 5908 2772 5918
rect 15596 5908 15652 6636
rect 15932 6020 15988 6030
rect 16044 6020 16100 9660
rect 16156 9602 16212 9614
rect 16156 9550 16158 9602
rect 16210 9550 16212 9602
rect 16156 9156 16212 9550
rect 16828 9604 16884 9774
rect 17276 9826 17332 9996
rect 17276 9774 17278 9826
rect 17330 9774 17332 9826
rect 17276 9762 17332 9774
rect 16828 9538 16884 9548
rect 17500 9604 17556 11230
rect 17724 11844 17780 11854
rect 17612 10610 17668 10622
rect 17612 10558 17614 10610
rect 17666 10558 17668 10610
rect 17612 9716 17668 10558
rect 17612 9650 17668 9660
rect 17724 10610 17780 11788
rect 17836 10724 17892 12126
rect 17948 12404 18004 12414
rect 17948 12178 18004 12348
rect 17948 12126 17950 12178
rect 18002 12126 18004 12178
rect 17948 11844 18004 12126
rect 17948 11778 18004 11788
rect 18060 11394 18116 12684
rect 18172 12404 18228 12414
rect 18172 11956 18228 12348
rect 18396 12180 18452 12190
rect 18508 12180 18564 12798
rect 18396 12178 18564 12180
rect 18396 12126 18398 12178
rect 18450 12126 18564 12178
rect 18396 12124 18564 12126
rect 19180 12850 19460 12852
rect 19180 12798 19406 12850
rect 19458 12798 19460 12850
rect 19180 12796 19460 12798
rect 18172 11890 18228 11900
rect 18284 11954 18340 11966
rect 18284 11902 18286 11954
rect 18338 11902 18340 11954
rect 18060 11342 18062 11394
rect 18114 11342 18116 11394
rect 18060 11330 18116 11342
rect 17836 10668 18004 10724
rect 17724 10558 17726 10610
rect 17778 10558 17780 10610
rect 17500 9538 17556 9548
rect 16156 9090 16212 9100
rect 16380 8484 16436 8494
rect 15932 6018 16100 6020
rect 15932 5966 15934 6018
rect 15986 5966 16100 6018
rect 15932 5964 16100 5966
rect 16156 8372 16212 8382
rect 16156 6018 16212 8316
rect 16156 5966 16158 6018
rect 16210 5966 16212 6018
rect 15932 5954 15988 5964
rect 16156 5954 16212 5966
rect 2268 5906 2772 5908
rect 2268 5854 2718 5906
rect 2770 5854 2772 5906
rect 2268 5852 2772 5854
rect 2156 5842 2212 5852
rect 2716 5842 2772 5852
rect 15260 5906 15652 5908
rect 15260 5854 15598 5906
rect 15650 5854 15652 5906
rect 15260 5852 15652 5854
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 15260 5122 15316 5852
rect 15596 5842 15652 5852
rect 16380 5906 16436 8428
rect 17724 8372 17780 10558
rect 17836 8484 17892 8494
rect 17948 8484 18004 10668
rect 18172 10500 18228 10510
rect 18172 10406 18228 10444
rect 18284 9826 18340 11902
rect 18396 11844 18452 12124
rect 18396 11778 18452 11788
rect 19180 11732 19236 12796
rect 19404 12786 19460 12796
rect 19292 12292 19348 12302
rect 19516 12292 19572 12302
rect 19292 12198 19348 12236
rect 19404 12236 19516 12292
rect 18956 11676 19236 11732
rect 18956 10610 19012 11676
rect 19404 11620 19460 12236
rect 19516 12226 19572 12236
rect 18956 10558 18958 10610
rect 19010 10558 19012 10610
rect 18508 10500 18564 10510
rect 18508 10406 18564 10444
rect 18284 9774 18286 9826
rect 18338 9774 18340 9826
rect 18284 9762 18340 9774
rect 18172 9604 18228 9614
rect 18172 9266 18228 9548
rect 18172 9214 18174 9266
rect 18226 9214 18228 9266
rect 18172 9202 18228 9214
rect 18620 9156 18676 9166
rect 18620 9062 18676 9100
rect 17892 8428 18004 8484
rect 18956 8484 19012 10558
rect 19068 11564 19460 11620
rect 19628 11620 19684 13020
rect 19852 13972 19908 13982
rect 19852 12964 19908 13916
rect 19852 12870 19908 12908
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19852 12404 19908 12414
rect 19740 12292 19796 12302
rect 19740 12198 19796 12236
rect 19068 9154 19124 11564
rect 19628 11554 19684 11564
rect 19852 11506 19908 12348
rect 20188 12180 20244 14252
rect 20300 14242 20356 14252
rect 20412 13524 20468 17388
rect 20524 16324 20580 17612
rect 20636 17666 20692 17678
rect 20636 17614 20638 17666
rect 20690 17614 20692 17666
rect 20636 16436 20692 17614
rect 20748 17444 20804 17454
rect 21084 17444 21140 18396
rect 20748 17442 21140 17444
rect 20748 17390 20750 17442
rect 20802 17390 21140 17442
rect 20748 17388 21140 17390
rect 21420 17666 21476 17678
rect 21420 17614 21422 17666
rect 21474 17614 21476 17666
rect 20748 17378 20804 17388
rect 21420 16436 21476 17614
rect 21532 17332 21588 18956
rect 21644 18946 21700 18956
rect 21756 18338 21812 18350
rect 21756 18286 21758 18338
rect 21810 18286 21812 18338
rect 21532 17266 21588 17276
rect 21644 17666 21700 17678
rect 21644 17614 21646 17666
rect 21698 17614 21700 17666
rect 21644 16772 21700 17614
rect 21644 16706 21700 16716
rect 20636 16380 21252 16436
rect 20524 16258 20580 16268
rect 20524 15876 20580 15886
rect 20524 15782 20580 15820
rect 20748 15204 20804 15242
rect 20748 15138 20804 15148
rect 20300 13468 20468 13524
rect 20524 14530 20580 14542
rect 20524 14478 20526 14530
rect 20578 14478 20580 14530
rect 20300 12402 20356 13468
rect 20524 13076 20580 14478
rect 21196 14532 21252 16380
rect 21420 16370 21476 16380
rect 21532 16658 21588 16670
rect 21532 16606 21534 16658
rect 21586 16606 21588 16658
rect 21308 15314 21364 15326
rect 21308 15262 21310 15314
rect 21362 15262 21364 15314
rect 21308 14980 21364 15262
rect 21532 15148 21588 16606
rect 21644 16548 21700 16558
rect 21644 16098 21700 16492
rect 21644 16046 21646 16098
rect 21698 16046 21700 16098
rect 21644 16034 21700 16046
rect 21644 15428 21700 15438
rect 21756 15428 21812 18286
rect 21868 17332 21924 21534
rect 22092 21476 22148 21756
rect 22316 21812 22372 21822
rect 22316 21718 22372 21756
rect 22092 21410 22148 21420
rect 22540 21364 22596 23102
rect 22652 22370 22708 23660
rect 22764 23622 22820 23660
rect 22876 24834 22932 24846
rect 22876 24782 22878 24834
rect 22930 24782 22932 24834
rect 22876 23826 22932 24782
rect 22876 23774 22878 23826
rect 22930 23774 22932 23826
rect 22876 22932 22932 23774
rect 22988 23492 23044 26236
rect 23100 26292 23156 26302
rect 23100 25506 23156 26236
rect 23100 25454 23102 25506
rect 23154 25454 23156 25506
rect 23100 25442 23156 25454
rect 22988 23426 23044 23436
rect 22876 22866 22932 22876
rect 23212 22820 23268 26852
rect 23660 26852 23828 26908
rect 23548 26292 23604 26302
rect 23548 26198 23604 26236
rect 23436 25396 23492 25406
rect 23436 25302 23492 25340
rect 23660 25172 23716 26852
rect 23772 25508 23828 25518
rect 23772 25414 23828 25452
rect 23660 25106 23716 25116
rect 23884 24948 23940 28588
rect 24220 28532 24276 28542
rect 23996 28084 24052 28094
rect 23996 27990 24052 28028
rect 24220 27636 24276 28476
rect 24332 28530 24388 29820
rect 24444 28644 24500 32508
rect 25340 32450 25396 32462
rect 25340 32398 25342 32450
rect 25394 32398 25396 32450
rect 25340 32116 25396 32398
rect 25340 32050 25396 32060
rect 25564 32452 25620 33516
rect 25676 33460 25732 33470
rect 25732 33404 25844 33460
rect 25676 33394 25732 33404
rect 25564 31892 25620 32396
rect 25340 31836 25620 31892
rect 25676 32674 25732 32686
rect 25676 32622 25678 32674
rect 25730 32622 25732 32674
rect 25228 31780 25284 31790
rect 25228 31686 25284 31724
rect 24556 30882 24612 30894
rect 24556 30830 24558 30882
rect 24610 30830 24612 30882
rect 24556 30212 24612 30830
rect 25228 30884 25284 30894
rect 25228 30790 25284 30828
rect 25340 30884 25396 31836
rect 25676 31780 25732 32622
rect 25452 31724 25732 31780
rect 25452 31666 25508 31724
rect 25788 31668 25844 33404
rect 26572 33236 26628 33246
rect 26348 33124 26404 33134
rect 25900 32564 25956 32574
rect 25956 32508 26180 32564
rect 25900 32470 25956 32508
rect 26124 31778 26180 32508
rect 26124 31726 26126 31778
rect 26178 31726 26180 31778
rect 26124 31714 26180 31726
rect 26348 31778 26404 33068
rect 26460 32452 26516 32462
rect 26572 32452 26628 33180
rect 26460 32450 26628 32452
rect 26460 32398 26462 32450
rect 26514 32398 26628 32450
rect 26460 32396 26628 32398
rect 26460 32386 26516 32396
rect 26348 31726 26350 31778
rect 26402 31726 26404 31778
rect 26348 31714 26404 31726
rect 25452 31614 25454 31666
rect 25506 31614 25508 31666
rect 25452 31220 25508 31614
rect 25676 31612 25844 31668
rect 26572 31666 26628 32396
rect 27020 32452 27076 35420
rect 27132 35252 27188 35646
rect 27132 35186 27188 35196
rect 27244 35922 27412 35924
rect 27244 35870 27358 35922
rect 27410 35870 27412 35922
rect 27244 35868 27412 35870
rect 27132 35028 27188 35038
rect 27244 35028 27300 35868
rect 27356 35858 27412 35868
rect 27692 36708 27748 36718
rect 27692 35698 27748 36652
rect 28140 36596 28196 36606
rect 28364 36596 28420 37326
rect 29260 38612 29316 38622
rect 28700 37268 28756 37278
rect 28700 37266 28980 37268
rect 28700 37214 28702 37266
rect 28754 37214 28980 37266
rect 28700 37212 28980 37214
rect 28700 37202 28756 37212
rect 28140 36594 28308 36596
rect 28140 36542 28142 36594
rect 28194 36542 28308 36594
rect 28140 36540 28308 36542
rect 28364 36540 28644 36596
rect 28140 36530 28196 36540
rect 27804 36258 27860 36270
rect 27804 36206 27806 36258
rect 27858 36206 27860 36258
rect 27804 36036 27860 36206
rect 27804 35970 27860 35980
rect 27692 35646 27694 35698
rect 27746 35646 27748 35698
rect 27692 35634 27748 35646
rect 28252 35698 28308 36540
rect 28252 35646 28254 35698
rect 28306 35646 28308 35698
rect 27132 35026 27300 35028
rect 27132 34974 27134 35026
rect 27186 34974 27300 35026
rect 27132 34972 27300 34974
rect 27580 35364 27636 35374
rect 27132 34962 27188 34972
rect 27580 34802 27636 35308
rect 28252 35364 28308 35646
rect 28252 35298 28308 35308
rect 28476 36372 28532 36382
rect 28476 35138 28532 36316
rect 28588 36258 28644 36540
rect 28588 36206 28590 36258
rect 28642 36206 28644 36258
rect 28588 36036 28644 36206
rect 28588 35970 28644 35980
rect 28476 35086 28478 35138
rect 28530 35086 28532 35138
rect 28476 35074 28532 35086
rect 27580 34750 27582 34802
rect 27634 34750 27636 34802
rect 27580 34738 27636 34750
rect 28028 33796 28084 33806
rect 28028 32564 28084 33740
rect 28588 33460 28644 33470
rect 28252 33236 28308 33246
rect 28252 33142 28308 33180
rect 28028 32470 28084 32508
rect 28588 32562 28644 33404
rect 28700 33124 28756 33134
rect 28700 33030 28756 33068
rect 28588 32510 28590 32562
rect 28642 32510 28644 32562
rect 28588 32498 28644 32510
rect 28700 32674 28756 32686
rect 28700 32622 28702 32674
rect 28754 32622 28756 32674
rect 27692 32452 27748 32462
rect 27020 32386 27076 32396
rect 27580 32450 27748 32452
rect 27580 32398 27694 32450
rect 27746 32398 27748 32450
rect 27580 32396 27748 32398
rect 27580 32228 27636 32396
rect 27692 32386 27748 32396
rect 26908 32172 27636 32228
rect 26908 32002 26964 32172
rect 26908 31950 26910 32002
rect 26962 31950 26964 32002
rect 26908 31938 26964 31950
rect 27020 32004 27076 32014
rect 26572 31614 26574 31666
rect 26626 31614 26628 31666
rect 25564 31556 25620 31566
rect 25564 31462 25620 31500
rect 25564 31220 25620 31230
rect 25452 31164 25564 31220
rect 25564 31154 25620 31164
rect 25564 30994 25620 31006
rect 25564 30942 25566 30994
rect 25618 30942 25620 30994
rect 25564 30884 25620 30942
rect 25340 30828 25620 30884
rect 25340 30660 25396 30828
rect 24556 30146 24612 30156
rect 25228 30604 25396 30660
rect 25228 30210 25284 30604
rect 25228 30158 25230 30210
rect 25282 30158 25284 30210
rect 25228 30146 25284 30158
rect 25340 30324 25396 30334
rect 24892 30100 24948 30110
rect 24892 30098 25172 30100
rect 24892 30046 24894 30098
rect 24946 30046 25172 30098
rect 24892 30044 25172 30046
rect 24892 30034 24948 30044
rect 25116 29652 25172 30044
rect 25228 29652 25284 29662
rect 25116 29650 25284 29652
rect 25116 29598 25230 29650
rect 25282 29598 25284 29650
rect 25116 29596 25284 29598
rect 25228 29586 25284 29596
rect 24892 29540 24948 29550
rect 24948 29484 25060 29540
rect 24892 29474 24948 29484
rect 24556 29428 24612 29438
rect 24556 29314 24612 29372
rect 24556 29262 24558 29314
rect 24610 29262 24612 29314
rect 24556 29250 24612 29262
rect 24556 28644 24612 28654
rect 24444 28642 24612 28644
rect 24444 28590 24558 28642
rect 24610 28590 24612 28642
rect 24444 28588 24612 28590
rect 24556 28578 24612 28588
rect 25004 28642 25060 29484
rect 25004 28590 25006 28642
rect 25058 28590 25060 28642
rect 25004 28578 25060 28590
rect 24332 28478 24334 28530
rect 24386 28478 24388 28530
rect 24332 28466 24388 28478
rect 25116 28532 25172 28542
rect 24892 28420 24948 28430
rect 24556 28084 24612 28094
rect 24332 27972 24388 27982
rect 24332 27970 24500 27972
rect 24332 27918 24334 27970
rect 24386 27918 24500 27970
rect 24332 27916 24500 27918
rect 24332 27906 24388 27916
rect 24220 27570 24276 27580
rect 24332 27412 24388 27422
rect 24332 27188 24388 27356
rect 24108 27186 24388 27188
rect 24108 27134 24334 27186
rect 24386 27134 24388 27186
rect 24108 27132 24388 27134
rect 23996 27076 24052 27086
rect 23996 26404 24052 27020
rect 24108 26514 24164 27132
rect 24332 27122 24388 27132
rect 24220 26908 24276 26918
rect 24276 26852 24388 26908
rect 24220 26842 24276 26852
rect 24108 26462 24110 26514
rect 24162 26462 24164 26514
rect 24108 26450 24164 26462
rect 24332 26404 24388 26852
rect 24444 26628 24500 27916
rect 24444 26562 24500 26572
rect 24444 26404 24500 26414
rect 24332 26402 24500 26404
rect 24332 26350 24446 26402
rect 24498 26350 24500 26402
rect 24332 26348 24500 26350
rect 23996 26338 24052 26348
rect 24444 26338 24500 26348
rect 24556 26402 24612 28028
rect 24668 27860 24724 27870
rect 24668 27858 24836 27860
rect 24668 27806 24670 27858
rect 24722 27806 24836 27858
rect 24668 27804 24836 27806
rect 24668 27794 24724 27804
rect 24668 27636 24724 27646
rect 24668 27186 24724 27580
rect 24668 27134 24670 27186
rect 24722 27134 24724 27186
rect 24668 27122 24724 27134
rect 24780 26964 24836 27804
rect 24892 27074 24948 28364
rect 24892 27022 24894 27074
rect 24946 27022 24948 27074
rect 24892 27010 24948 27022
rect 25004 27636 25060 27646
rect 24556 26350 24558 26402
rect 24610 26350 24612 26402
rect 24108 26068 24164 26078
rect 24108 25506 24164 26012
rect 24556 25732 24612 26350
rect 24108 25454 24110 25506
rect 24162 25454 24164 25506
rect 24108 25442 24164 25454
rect 24444 25676 24612 25732
rect 24668 26852 24836 26908
rect 23996 25282 24052 25294
rect 23996 25230 23998 25282
rect 24050 25230 24052 25282
rect 23996 25172 24052 25230
rect 23996 25106 24052 25116
rect 23884 24892 24164 24948
rect 23324 24724 23380 24734
rect 23324 23940 23380 24668
rect 23884 24722 23940 24734
rect 23884 24670 23886 24722
rect 23938 24670 23940 24722
rect 23324 23846 23380 23884
rect 23548 24498 23604 24510
rect 23548 24446 23550 24498
rect 23602 24446 23604 24498
rect 23548 23828 23604 24446
rect 23548 23762 23604 23772
rect 23660 23826 23716 23838
rect 23660 23774 23662 23826
rect 23714 23774 23716 23826
rect 23436 23716 23492 23726
rect 23436 23154 23492 23660
rect 23436 23102 23438 23154
rect 23490 23102 23492 23154
rect 23436 23090 23492 23102
rect 23548 23266 23604 23278
rect 23548 23214 23550 23266
rect 23602 23214 23604 23266
rect 23212 22754 23268 22764
rect 23436 22932 23492 22942
rect 23548 22932 23604 23214
rect 23492 22876 23604 22932
rect 23324 22484 23380 22494
rect 23436 22484 23492 22876
rect 23380 22428 23492 22484
rect 23324 22418 23380 22428
rect 23212 22372 23268 22382
rect 22652 22318 22654 22370
rect 22706 22318 22708 22370
rect 22652 22306 22708 22318
rect 22764 22370 23268 22372
rect 22764 22318 23214 22370
rect 23266 22318 23268 22370
rect 22764 22316 23268 22318
rect 22652 21810 22708 21822
rect 22652 21758 22654 21810
rect 22706 21758 22708 21810
rect 22652 21588 22708 21758
rect 22652 21522 22708 21532
rect 22540 21298 22596 21308
rect 22652 21028 22708 21038
rect 22764 21028 22820 22316
rect 23212 22306 23268 22316
rect 23436 22258 23492 22428
rect 23436 22206 23438 22258
rect 23490 22206 23492 22258
rect 23436 22194 23492 22206
rect 23548 22708 23604 22718
rect 23100 22148 23156 22158
rect 23324 22148 23380 22158
rect 23100 21586 23156 22092
rect 23100 21534 23102 21586
rect 23154 21534 23156 21586
rect 23100 21522 23156 21534
rect 23212 22146 23380 22148
rect 23212 22094 23326 22146
rect 23378 22094 23380 22146
rect 23212 22092 23380 22094
rect 23212 21474 23268 22092
rect 23324 22082 23380 22092
rect 23548 22036 23604 22652
rect 23436 21980 23604 22036
rect 23436 21586 23492 21980
rect 23436 21534 23438 21586
rect 23490 21534 23492 21586
rect 23436 21522 23492 21534
rect 23212 21422 23214 21474
rect 23266 21422 23268 21474
rect 23212 21410 23268 21422
rect 23324 21364 23380 21374
rect 23380 21308 23492 21364
rect 23324 21298 23380 21308
rect 22652 21026 22820 21028
rect 22652 20974 22654 21026
rect 22706 20974 22820 21026
rect 22652 20972 22820 20974
rect 22652 20962 22708 20972
rect 22876 20916 22932 20926
rect 22764 20860 22876 20916
rect 22092 20580 22148 20590
rect 21980 20524 22092 20580
rect 21980 17778 22036 20524
rect 22092 20514 22148 20524
rect 22540 20130 22596 20142
rect 22540 20078 22542 20130
rect 22594 20078 22596 20130
rect 22540 19908 22596 20078
rect 22540 18564 22596 19852
rect 22540 18498 22596 18508
rect 22764 19348 22820 20860
rect 22876 20850 22932 20860
rect 22988 20802 23044 20814
rect 22988 20750 22990 20802
rect 23042 20750 23044 20802
rect 22988 20244 23044 20750
rect 23212 20690 23268 20702
rect 23212 20638 23214 20690
rect 23266 20638 23268 20690
rect 23100 20244 23156 20254
rect 22988 20242 23156 20244
rect 22988 20190 23102 20242
rect 23154 20190 23156 20242
rect 22988 20188 23156 20190
rect 23100 20178 23156 20188
rect 23212 19460 23268 20638
rect 22652 18452 22708 18462
rect 22764 18452 22820 19292
rect 22652 18450 22820 18452
rect 22652 18398 22654 18450
rect 22706 18398 22820 18450
rect 22652 18396 22820 18398
rect 23100 19404 23268 19460
rect 23100 18452 23156 19404
rect 22652 18386 22708 18396
rect 23100 18386 23156 18396
rect 23212 19234 23268 19246
rect 23212 19182 23214 19234
rect 23266 19182 23268 19234
rect 21980 17726 21982 17778
rect 22034 17726 22036 17778
rect 21980 17714 22036 17726
rect 22876 17780 22932 17790
rect 21980 17556 22036 17566
rect 21980 17462 22036 17500
rect 22204 17554 22260 17566
rect 22204 17502 22206 17554
rect 22258 17502 22260 17554
rect 21868 17276 22148 17332
rect 21868 16882 21924 16894
rect 21868 16830 21870 16882
rect 21922 16830 21924 16882
rect 21868 16660 21924 16830
rect 21868 16594 21924 16604
rect 21868 16436 21924 16446
rect 21924 16380 22036 16436
rect 21868 16370 21924 16380
rect 21644 15426 21812 15428
rect 21644 15374 21646 15426
rect 21698 15374 21812 15426
rect 21644 15372 21812 15374
rect 21868 16100 21924 16110
rect 21868 15538 21924 16044
rect 21868 15486 21870 15538
rect 21922 15486 21924 15538
rect 21644 15362 21700 15372
rect 21868 15148 21924 15486
rect 21308 14914 21364 14924
rect 21420 15092 21588 15148
rect 21644 15092 21924 15148
rect 21980 15202 22036 16380
rect 21980 15150 21982 15202
rect 22034 15150 22036 15202
rect 21980 15138 22036 15150
rect 21308 14756 21364 14766
rect 21420 14756 21476 15092
rect 21308 14754 21476 14756
rect 21308 14702 21310 14754
rect 21362 14702 21476 14754
rect 21308 14700 21476 14702
rect 21308 14690 21364 14700
rect 21420 14532 21476 14542
rect 21196 14530 21476 14532
rect 21196 14478 21422 14530
rect 21474 14478 21476 14530
rect 21196 14476 21476 14478
rect 21420 14466 21476 14476
rect 21644 14530 21700 15092
rect 21644 14478 21646 14530
rect 21698 14478 21700 14530
rect 21644 14466 21700 14478
rect 20524 13010 20580 13020
rect 20412 12964 20468 12974
rect 20412 12870 20468 12908
rect 20300 12350 20302 12402
rect 20354 12350 20356 12402
rect 20300 12338 20356 12350
rect 21532 12852 21588 12862
rect 21532 12402 21588 12796
rect 21532 12350 21534 12402
rect 21586 12350 21588 12402
rect 21532 12338 21588 12350
rect 21084 12290 21140 12302
rect 21084 12238 21086 12290
rect 21138 12238 21140 12290
rect 20188 12124 20356 12180
rect 19852 11454 19854 11506
rect 19906 11454 19908 11506
rect 19852 11442 19908 11454
rect 19964 11954 20020 11966
rect 19964 11902 19966 11954
rect 20018 11902 20020 11954
rect 19180 11396 19236 11406
rect 19628 11396 19684 11406
rect 19180 11394 19684 11396
rect 19180 11342 19182 11394
rect 19234 11342 19630 11394
rect 19682 11342 19684 11394
rect 19180 11340 19684 11342
rect 19180 11330 19236 11340
rect 19628 11330 19684 11340
rect 19964 11172 20020 11902
rect 19516 11116 20020 11172
rect 20076 11844 20132 11854
rect 20076 11394 20132 11788
rect 20076 11342 20078 11394
rect 20130 11342 20132 11394
rect 20076 11172 20132 11342
rect 20076 11116 20244 11172
rect 19516 10834 19572 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20188 10836 20244 11116
rect 19516 10782 19518 10834
rect 19570 10782 19572 10834
rect 19516 10770 19572 10782
rect 20076 10780 20244 10836
rect 19292 10610 19348 10622
rect 19292 10558 19294 10610
rect 19346 10558 19348 10610
rect 19292 9938 19348 10558
rect 19964 10612 20020 10622
rect 19964 10518 20020 10556
rect 19292 9886 19294 9938
rect 19346 9886 19348 9938
rect 19292 9874 19348 9886
rect 19628 10164 19684 10174
rect 19068 9102 19070 9154
rect 19122 9102 19124 9154
rect 19068 9090 19124 9102
rect 19628 9044 19684 10108
rect 20076 9828 20132 10780
rect 20188 9828 20244 9838
rect 20076 9772 20188 9828
rect 20188 9734 20244 9772
rect 19964 9714 20020 9726
rect 19964 9662 19966 9714
rect 20018 9662 20020 9714
rect 19964 9604 20020 9662
rect 19964 9548 20244 9604
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19964 9044 20020 9054
rect 19628 8988 19796 9044
rect 19292 8820 19348 8830
rect 19628 8820 19684 8830
rect 19292 8818 19572 8820
rect 19292 8766 19294 8818
rect 19346 8766 19572 8818
rect 19292 8764 19572 8766
rect 19292 8754 19348 8764
rect 18956 8428 19348 8484
rect 17836 8418 17892 8428
rect 17724 8306 17780 8316
rect 18732 8260 18788 8270
rect 19180 8260 19236 8270
rect 18732 8166 18788 8204
rect 19068 8258 19236 8260
rect 19068 8206 19182 8258
rect 19234 8206 19236 8258
rect 19068 8204 19236 8206
rect 18844 8036 18900 8046
rect 18844 7474 18900 7980
rect 18844 7422 18846 7474
rect 18898 7422 18900 7474
rect 18844 7410 18900 7422
rect 18956 8034 19012 8046
rect 18956 7982 18958 8034
rect 19010 7982 19012 8034
rect 18284 6468 18340 6478
rect 18284 6374 18340 6412
rect 18508 6132 18564 6142
rect 16380 5854 16382 5906
rect 16434 5854 16436 5906
rect 16380 5842 16436 5854
rect 17500 6018 17556 6030
rect 17500 5966 17502 6018
rect 17554 5966 17556 6018
rect 15260 5070 15262 5122
rect 15314 5070 15316 5122
rect 15260 5058 15316 5070
rect 16716 5682 16772 5694
rect 16716 5630 16718 5682
rect 16770 5630 16772 5682
rect 1708 4900 1764 4910
rect 1708 4806 1764 4844
rect 16716 4564 16772 5630
rect 16716 4498 16772 4508
rect 17500 4338 17556 5966
rect 18508 6018 18564 6076
rect 18956 6132 19012 7982
rect 18956 6066 19012 6076
rect 19068 7586 19124 8204
rect 19180 8194 19236 8204
rect 19068 7534 19070 7586
rect 19122 7534 19124 7586
rect 18508 5966 18510 6018
rect 18562 5966 18564 6018
rect 18508 5954 18564 5966
rect 18620 5908 18676 5918
rect 17500 4286 17502 4338
rect 17554 4286 17556 4338
rect 17500 4274 17556 4286
rect 18508 4898 18564 4910
rect 18508 4846 18510 4898
rect 18562 4846 18564 4898
rect 18508 4338 18564 4846
rect 18508 4286 18510 4338
rect 18562 4286 18564 4338
rect 18508 4274 18564 4286
rect 18620 4116 18676 5852
rect 19068 5124 19124 7534
rect 19292 7028 19348 8428
rect 19516 7588 19572 8764
rect 19628 8726 19684 8764
rect 19740 8258 19796 8988
rect 19740 8206 19742 8258
rect 19794 8206 19796 8258
rect 19740 8194 19796 8206
rect 19964 8146 20020 8988
rect 19964 8094 19966 8146
rect 20018 8094 20020 8146
rect 19964 8082 20020 8094
rect 20188 8930 20244 9548
rect 20188 8878 20190 8930
rect 20242 8878 20244 8930
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19516 7532 19684 7588
rect 19180 6972 19348 7028
rect 19516 7362 19572 7374
rect 19516 7310 19518 7362
rect 19570 7310 19572 7362
rect 19180 6692 19236 6972
rect 19180 6626 19236 6636
rect 19292 6804 19348 6814
rect 19516 6804 19572 7310
rect 19292 6802 19572 6804
rect 19292 6750 19294 6802
rect 19346 6750 19572 6802
rect 19292 6748 19572 6750
rect 19292 5908 19348 6748
rect 19292 5842 19348 5852
rect 19068 5058 19124 5068
rect 19180 5684 19236 5694
rect 19180 4450 19236 5628
rect 19628 4562 19684 7532
rect 19852 7586 19908 7598
rect 19852 7534 19854 7586
rect 19906 7534 19908 7586
rect 19852 6578 19908 7534
rect 19852 6526 19854 6578
rect 19906 6526 19908 6578
rect 19852 6468 19908 6526
rect 20188 6580 20244 8878
rect 20300 8258 20356 12124
rect 20748 12178 20804 12190
rect 20748 12126 20750 12178
rect 20802 12126 20804 12178
rect 20748 11732 20804 12126
rect 20748 11666 20804 11676
rect 21084 11284 21140 12238
rect 21308 11620 21364 11630
rect 21308 11394 21364 11564
rect 21308 11342 21310 11394
rect 21362 11342 21364 11394
rect 21308 11330 21364 11342
rect 20636 11228 21140 11284
rect 20636 10164 20692 11228
rect 21420 11172 21476 11182
rect 20748 11170 21476 11172
rect 20748 11118 21422 11170
rect 21474 11118 21476 11170
rect 20748 11116 21476 11118
rect 20748 10610 20804 11116
rect 21420 11106 21476 11116
rect 20748 10558 20750 10610
rect 20802 10558 20804 10610
rect 20748 10546 20804 10558
rect 21644 10612 21700 10622
rect 21644 10610 21812 10612
rect 21644 10558 21646 10610
rect 21698 10558 21812 10610
rect 21644 10556 21812 10558
rect 21644 10546 21700 10556
rect 20636 10098 20692 10108
rect 21756 10052 21812 10556
rect 21868 10052 21924 10062
rect 21756 10050 21924 10052
rect 21756 9998 21870 10050
rect 21922 9998 21924 10050
rect 21756 9996 21924 9998
rect 21868 9986 21924 9996
rect 21644 9940 21700 9950
rect 21308 9828 21364 9838
rect 21308 9734 21364 9772
rect 20636 9604 20692 9614
rect 20636 9510 20692 9548
rect 20636 9044 20692 9054
rect 20636 8950 20692 8988
rect 20300 8206 20302 8258
rect 20354 8206 20356 8258
rect 20300 8194 20356 8206
rect 21644 8258 21700 9884
rect 22092 8932 22148 17276
rect 22204 17108 22260 17502
rect 22876 17556 22932 17724
rect 23212 17668 23268 19182
rect 23436 18450 23492 21308
rect 23660 21252 23716 23774
rect 23772 22708 23828 22718
rect 23884 22708 23940 24670
rect 23996 24610 24052 24622
rect 23996 24558 23998 24610
rect 24050 24558 24052 24610
rect 23996 23378 24052 24558
rect 23996 23326 23998 23378
rect 24050 23326 24052 23378
rect 23996 23314 24052 23326
rect 24108 23156 24164 24892
rect 24220 24724 24276 24734
rect 24220 24630 24276 24668
rect 24444 24052 24500 25676
rect 24444 23986 24500 23996
rect 24556 25508 24612 25518
rect 24668 25508 24724 26852
rect 24780 26516 24836 26526
rect 24780 26422 24836 26460
rect 25004 25844 25060 27580
rect 25116 27188 25172 28476
rect 25340 28530 25396 30268
rect 25564 29316 25620 29326
rect 25564 29222 25620 29260
rect 25340 28478 25342 28530
rect 25394 28478 25396 28530
rect 25340 28466 25396 28478
rect 25676 28308 25732 31612
rect 26124 31556 26180 31566
rect 26124 30994 26180 31500
rect 26124 30942 26126 30994
rect 26178 30942 26180 30994
rect 26124 30930 26180 30942
rect 26236 31106 26292 31118
rect 26236 31054 26238 31106
rect 26290 31054 26292 31106
rect 25788 30212 25844 30222
rect 25788 30118 25844 30156
rect 25900 29988 25956 29998
rect 25900 29986 26068 29988
rect 25900 29934 25902 29986
rect 25954 29934 26068 29986
rect 25900 29932 26068 29934
rect 25900 29922 25956 29932
rect 25788 29876 25844 29886
rect 25788 29540 25844 29820
rect 25788 29426 25844 29484
rect 25788 29374 25790 29426
rect 25842 29374 25844 29426
rect 25788 29362 25844 29374
rect 25228 28252 25732 28308
rect 25228 27970 25284 28252
rect 25340 28084 25396 28094
rect 25340 27990 25396 28028
rect 25228 27918 25230 27970
rect 25282 27918 25284 27970
rect 25228 27906 25284 27918
rect 26012 27970 26068 29932
rect 26012 27918 26014 27970
rect 26066 27918 26068 27970
rect 26012 27906 26068 27918
rect 26124 27972 26180 27982
rect 26124 27878 26180 27916
rect 25116 27122 25172 27132
rect 25564 27858 25620 27870
rect 25564 27806 25566 27858
rect 25618 27806 25620 27858
rect 25340 27076 25396 27114
rect 25340 27010 25396 27020
rect 25452 27074 25508 27086
rect 25452 27022 25454 27074
rect 25506 27022 25508 27074
rect 25452 26964 25508 27022
rect 25452 26898 25508 26908
rect 25228 26850 25284 26862
rect 25228 26798 25230 26850
rect 25282 26798 25284 26850
rect 24556 25506 24724 25508
rect 24556 25454 24558 25506
rect 24610 25454 24724 25506
rect 24556 25452 24724 25454
rect 24780 25788 25060 25844
rect 25116 26628 25172 26638
rect 23828 22652 23940 22708
rect 23996 23100 24164 23156
rect 24220 23940 24276 23950
rect 24220 23156 24276 23884
rect 24332 23938 24388 23950
rect 24332 23886 24334 23938
rect 24386 23886 24388 23938
rect 24332 23828 24388 23886
rect 24332 23772 24500 23828
rect 24444 23604 24500 23772
rect 24556 23826 24612 25452
rect 24556 23774 24558 23826
rect 24610 23774 24612 23826
rect 24556 23762 24612 23774
rect 24780 23604 24836 25788
rect 25004 25620 25060 25630
rect 25004 25526 25060 25564
rect 25116 24276 25172 26572
rect 25228 26290 25284 26798
rect 25228 26238 25230 26290
rect 25282 26238 25284 26290
rect 25228 26226 25284 26238
rect 25564 26068 25620 27806
rect 26124 27634 26180 27646
rect 26124 27582 26126 27634
rect 26178 27582 26180 27634
rect 25788 27074 25844 27086
rect 25788 27022 25790 27074
rect 25842 27022 25844 27074
rect 25788 26516 25844 27022
rect 26124 27074 26180 27582
rect 26124 27022 26126 27074
rect 26178 27022 26180 27074
rect 26124 27010 26180 27022
rect 25788 26450 25844 26460
rect 26012 26962 26068 26974
rect 26012 26910 26014 26962
rect 26066 26910 26068 26962
rect 25340 26012 25620 26068
rect 25676 26290 25732 26302
rect 25676 26238 25678 26290
rect 25730 26238 25732 26290
rect 25340 25506 25396 26012
rect 25340 25454 25342 25506
rect 25394 25454 25396 25506
rect 25340 25442 25396 25454
rect 25564 25508 25620 25518
rect 25564 25414 25620 25452
rect 25452 25284 25508 25294
rect 24444 23548 24836 23604
rect 24892 24220 25172 24276
rect 25340 25282 25508 25284
rect 25340 25230 25454 25282
rect 25506 25230 25508 25282
rect 25340 25228 25508 25230
rect 24220 23154 24388 23156
rect 24220 23102 24222 23154
rect 24274 23102 24388 23154
rect 24220 23100 24388 23102
rect 23772 22642 23828 22652
rect 23996 21812 24052 23100
rect 24220 23090 24276 23100
rect 24332 22932 24388 23100
rect 24220 22876 24388 22932
rect 24220 22370 24276 22876
rect 24220 22318 24222 22370
rect 24274 22318 24276 22370
rect 24220 22306 24276 22318
rect 24332 22260 24388 22270
rect 24332 22166 24388 22204
rect 24444 22036 24500 23548
rect 24556 23380 24612 23390
rect 24556 23266 24612 23324
rect 24556 23214 24558 23266
rect 24610 23214 24612 23266
rect 24556 23202 24612 23214
rect 24444 21970 24500 21980
rect 24668 22708 24724 22718
rect 24332 21812 24388 21822
rect 23996 21810 24388 21812
rect 23996 21758 24334 21810
rect 24386 21758 24388 21810
rect 23996 21756 24388 21758
rect 24332 21746 24388 21756
rect 24668 21698 24724 22652
rect 24668 21646 24670 21698
rect 24722 21646 24724 21698
rect 23660 21196 23940 21252
rect 23772 20690 23828 20702
rect 23772 20638 23774 20690
rect 23826 20638 23828 20690
rect 23772 20356 23828 20638
rect 23884 20580 23940 21196
rect 24332 20580 24388 20590
rect 23884 20578 24388 20580
rect 23884 20526 24334 20578
rect 24386 20526 24388 20578
rect 23884 20524 24388 20526
rect 24668 20580 24724 21646
rect 24892 21476 24948 24220
rect 25340 24164 25396 25228
rect 25452 25218 25508 25228
rect 25676 25284 25732 26238
rect 25004 24108 25396 24164
rect 25676 24722 25732 25228
rect 25676 24670 25678 24722
rect 25730 24670 25732 24722
rect 25004 23938 25060 24108
rect 25004 23886 25006 23938
rect 25058 23886 25060 23938
rect 25004 23874 25060 23886
rect 25340 23940 25396 23950
rect 25676 23940 25732 24670
rect 25340 23938 25508 23940
rect 25340 23886 25342 23938
rect 25394 23886 25508 23938
rect 25340 23884 25508 23886
rect 25340 23874 25396 23884
rect 25228 23828 25284 23838
rect 25452 23828 25508 23884
rect 25564 23884 25732 23940
rect 25900 25394 25956 25406
rect 25900 25342 25902 25394
rect 25954 25342 25956 25394
rect 25564 23828 25620 23884
rect 25452 23772 25620 23828
rect 25788 23826 25844 23838
rect 25788 23774 25790 23826
rect 25842 23774 25844 23826
rect 25228 23154 25284 23772
rect 25676 23716 25732 23726
rect 25676 23266 25732 23660
rect 25676 23214 25678 23266
rect 25730 23214 25732 23266
rect 25676 23202 25732 23214
rect 25788 23268 25844 23774
rect 25900 23380 25956 25342
rect 26012 24610 26068 26910
rect 26124 26180 26180 26190
rect 26124 26086 26180 26124
rect 26236 26068 26292 31054
rect 26572 30660 26628 31614
rect 26796 31444 26852 31454
rect 26572 30594 26628 30604
rect 26684 31220 26740 31230
rect 26348 30324 26404 30334
rect 26348 30210 26404 30268
rect 26348 30158 26350 30210
rect 26402 30158 26404 30210
rect 26348 30146 26404 30158
rect 26684 29428 26740 31164
rect 26796 30994 26852 31388
rect 26796 30942 26798 30994
rect 26850 30942 26852 30994
rect 26796 30324 26852 30942
rect 26796 30258 26852 30268
rect 26796 29428 26852 29438
rect 26684 29426 26852 29428
rect 26684 29374 26798 29426
rect 26850 29374 26852 29426
rect 26684 29372 26852 29374
rect 26796 29362 26852 29372
rect 26908 27858 26964 27870
rect 26908 27806 26910 27858
rect 26962 27806 26964 27858
rect 26348 27074 26404 27086
rect 26348 27022 26350 27074
rect 26402 27022 26404 27074
rect 26348 26964 26404 27022
rect 26908 27076 26964 27806
rect 26908 27010 26964 27020
rect 26348 26898 26404 26908
rect 26572 26964 26628 26974
rect 26236 26002 26292 26012
rect 26348 26402 26404 26414
rect 26348 26350 26350 26402
rect 26402 26350 26404 26402
rect 26348 25620 26404 26350
rect 26572 25730 26628 26908
rect 26796 26852 26852 26862
rect 26796 26290 26852 26796
rect 26796 26238 26798 26290
rect 26850 26238 26852 26290
rect 26796 26226 26852 26238
rect 26572 25678 26574 25730
rect 26626 25678 26628 25730
rect 26572 25666 26628 25678
rect 26236 25506 26292 25518
rect 26236 25454 26238 25506
rect 26290 25454 26292 25506
rect 26236 25284 26292 25454
rect 26236 25218 26292 25228
rect 26348 24834 26404 25564
rect 27020 25396 27076 31948
rect 27244 32004 27300 32014
rect 27132 30212 27188 30222
rect 27132 30118 27188 30156
rect 27132 27972 27188 27982
rect 27132 26908 27188 27916
rect 27244 27970 27300 31948
rect 28700 32004 28756 32622
rect 28700 31938 28756 31948
rect 27804 31892 27860 31902
rect 27804 31798 27860 31836
rect 28364 31780 28420 31790
rect 28364 31686 28420 31724
rect 27580 31556 27636 31566
rect 27356 30994 27412 31006
rect 27356 30942 27358 30994
rect 27410 30942 27412 30994
rect 27356 29650 27412 30942
rect 27356 29598 27358 29650
rect 27410 29598 27412 29650
rect 27356 29586 27412 29598
rect 27244 27918 27246 27970
rect 27298 27918 27300 27970
rect 27244 27906 27300 27918
rect 27580 26964 27636 31500
rect 28028 31108 28084 31118
rect 27692 30212 27748 30222
rect 27692 29650 27748 30156
rect 28028 30210 28084 31052
rect 28812 31108 28868 31118
rect 28812 31014 28868 31052
rect 28028 30158 28030 30210
rect 28082 30158 28084 30210
rect 28028 30146 28084 30158
rect 28364 30994 28420 31006
rect 28364 30942 28366 30994
rect 28418 30942 28420 30994
rect 28364 30212 28420 30942
rect 28924 30660 28980 37212
rect 29260 37156 29316 38556
rect 29708 37492 29764 37502
rect 30044 37492 30100 38668
rect 30828 38612 30884 40350
rect 31164 38668 31220 43484
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 33516 42642 33572 42654
rect 33516 42590 33518 42642
rect 33570 42590 33572 42642
rect 31724 42084 31780 42094
rect 31724 41972 31780 42028
rect 33516 42084 33572 42590
rect 46172 42530 46228 42542
rect 46172 42478 46174 42530
rect 46226 42478 46228 42530
rect 46172 42420 46228 42478
rect 46172 42354 46228 42364
rect 33516 41990 33572 42028
rect 31388 41970 31780 41972
rect 31388 41918 31726 41970
rect 31778 41918 31780 41970
rect 31388 41916 31780 41918
rect 31388 41186 31444 41916
rect 31724 41906 31780 41916
rect 32508 41972 32564 41982
rect 32508 41878 32564 41916
rect 33628 41972 33684 41982
rect 31388 41134 31390 41186
rect 31442 41134 31444 41186
rect 31388 41122 31444 41134
rect 31724 41188 31780 41198
rect 31780 41132 31892 41188
rect 31724 41122 31780 41132
rect 31724 40628 31780 40638
rect 31276 40404 31332 40414
rect 31276 40310 31332 40348
rect 31164 38612 31332 38668
rect 30828 38546 30884 38556
rect 29708 37490 30100 37492
rect 29708 37438 29710 37490
rect 29762 37438 30046 37490
rect 30098 37438 30100 37490
rect 29708 37436 30100 37438
rect 29708 37426 29764 37436
rect 30044 37426 30100 37436
rect 31276 37380 31332 38612
rect 31724 38050 31780 40572
rect 31836 40402 31892 41132
rect 31836 40350 31838 40402
rect 31890 40350 31892 40402
rect 31836 40338 31892 40350
rect 32284 41186 32340 41198
rect 32284 41134 32286 41186
rect 32338 41134 32340 41186
rect 32284 39844 32340 41134
rect 32284 39778 32340 39788
rect 33628 39618 33684 41916
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35084 40628 35140 40638
rect 35084 40402 35140 40572
rect 37884 40514 37940 40526
rect 37884 40462 37886 40514
rect 37938 40462 37940 40514
rect 35084 40350 35086 40402
rect 35138 40350 35140 40402
rect 35084 40338 35140 40350
rect 35532 40404 35588 40414
rect 35532 40310 35588 40348
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 34188 39844 34244 39854
rect 34188 39750 34244 39788
rect 33628 39566 33630 39618
rect 33682 39566 33684 39618
rect 33180 39506 33236 39518
rect 33180 39454 33182 39506
rect 33234 39454 33236 39506
rect 33180 39396 33236 39454
rect 33180 39330 33236 39340
rect 33068 39284 33124 39294
rect 32508 38946 32564 38958
rect 32508 38894 32510 38946
rect 32562 38894 32564 38946
rect 31724 37998 31726 38050
rect 31778 37998 31780 38050
rect 31724 37986 31780 37998
rect 32284 38834 32340 38846
rect 32284 38782 32286 38834
rect 32338 38782 32340 38834
rect 32284 38612 32340 38782
rect 30380 37266 30436 37278
rect 30380 37214 30382 37266
rect 30434 37214 30436 37266
rect 29260 37154 29764 37156
rect 29260 37102 29262 37154
rect 29314 37102 29764 37154
rect 29260 37100 29764 37102
rect 29260 37090 29316 37100
rect 29372 36932 29428 36942
rect 29148 36372 29204 36382
rect 29148 36278 29204 36316
rect 29148 35252 29204 35262
rect 29148 34914 29204 35196
rect 29148 34862 29150 34914
rect 29202 34862 29204 34914
rect 29148 34850 29204 34862
rect 29372 34914 29428 36876
rect 29372 34862 29374 34914
rect 29426 34862 29428 34914
rect 29372 34850 29428 34862
rect 29484 36482 29540 36494
rect 29484 36430 29486 36482
rect 29538 36430 29540 36482
rect 29484 33796 29540 36430
rect 29708 34914 29764 37100
rect 29708 34862 29710 34914
rect 29762 34862 29764 34914
rect 29708 34850 29764 34862
rect 29932 36482 29988 36494
rect 29932 36430 29934 36482
rect 29986 36430 29988 36482
rect 29932 34354 29988 36430
rect 30156 36260 30212 36270
rect 30156 36166 30212 36204
rect 30156 35252 30212 35262
rect 30156 34914 30212 35196
rect 30156 34862 30158 34914
rect 30210 34862 30212 34914
rect 30156 34850 30212 34862
rect 29932 34302 29934 34354
rect 29986 34302 29988 34354
rect 29932 34290 29988 34302
rect 29484 33730 29540 33740
rect 29260 33460 29316 33470
rect 29260 33366 29316 33404
rect 29036 33346 29092 33358
rect 29708 33348 29764 33358
rect 29036 33294 29038 33346
rect 29090 33294 29092 33346
rect 29036 33236 29092 33294
rect 29036 33170 29092 33180
rect 29596 33292 29708 33348
rect 29596 33234 29652 33292
rect 29708 33282 29764 33292
rect 29596 33182 29598 33234
rect 29650 33182 29652 33234
rect 29372 33124 29428 33134
rect 29428 33068 29540 33124
rect 29372 33030 29428 33068
rect 29372 32562 29428 32574
rect 29372 32510 29374 32562
rect 29426 32510 29428 32562
rect 29260 31892 29316 31902
rect 29260 31778 29316 31836
rect 29260 31726 29262 31778
rect 29314 31726 29316 31778
rect 29148 31220 29204 31230
rect 29260 31220 29316 31726
rect 29372 31444 29428 32510
rect 29484 31556 29540 33068
rect 29596 31780 29652 33182
rect 29820 32562 29876 32574
rect 29820 32510 29822 32562
rect 29874 32510 29876 32562
rect 29820 32002 29876 32510
rect 29820 31950 29822 32002
rect 29874 31950 29876 32002
rect 29820 31938 29876 31950
rect 29596 31714 29652 31724
rect 30268 31780 30324 31790
rect 29484 31490 29540 31500
rect 29372 31378 29428 31388
rect 29148 31218 29540 31220
rect 29148 31166 29150 31218
rect 29202 31166 29540 31218
rect 29148 31164 29540 31166
rect 29148 31154 29204 31164
rect 29484 30996 29540 31164
rect 29484 30994 29876 30996
rect 29484 30942 29486 30994
rect 29538 30942 29876 30994
rect 29484 30940 29876 30942
rect 29484 30930 29540 30940
rect 28924 30604 29428 30660
rect 28364 30146 28420 30156
rect 29148 30212 29204 30222
rect 29148 30118 29204 30156
rect 27692 29598 27694 29650
rect 27746 29598 27748 29650
rect 27692 29586 27748 29598
rect 28252 29988 28308 29998
rect 27804 29540 27860 29550
rect 27804 29446 27860 29484
rect 28140 28980 28196 28990
rect 28140 28866 28196 28924
rect 28140 28814 28142 28866
rect 28194 28814 28196 28866
rect 28140 28802 28196 28814
rect 27692 28644 27748 28654
rect 27692 28550 27748 28588
rect 28252 27076 28308 29932
rect 28476 29540 28532 29550
rect 28364 28756 28420 28766
rect 28364 28662 28420 28700
rect 28476 27972 28532 29484
rect 28588 29426 28644 29438
rect 28588 29374 28590 29426
rect 28642 29374 28644 29426
rect 28588 28756 28644 29374
rect 29260 29428 29316 29438
rect 29260 29334 29316 29372
rect 28924 28980 28980 28990
rect 28588 28754 28868 28756
rect 28588 28702 28590 28754
rect 28642 28702 28868 28754
rect 28588 28700 28868 28702
rect 28588 28690 28644 28700
rect 28812 28082 28868 28700
rect 28812 28030 28814 28082
rect 28866 28030 28868 28082
rect 28812 28018 28868 28030
rect 27468 26962 27636 26964
rect 27468 26910 27582 26962
rect 27634 26910 27636 26962
rect 27468 26908 27636 26910
rect 27132 26852 27412 26908
rect 27356 25508 27412 26852
rect 27468 26514 27524 26908
rect 27580 26898 27636 26908
rect 27804 27020 28308 27076
rect 27468 26462 27470 26514
rect 27522 26462 27524 26514
rect 27468 26292 27524 26462
rect 27468 26226 27524 26236
rect 27804 26290 27860 27020
rect 28252 26962 28308 27020
rect 28252 26910 28254 26962
rect 28306 26910 28308 26962
rect 28252 26898 28308 26910
rect 28364 27916 28532 27972
rect 28588 27972 28644 27982
rect 27916 26850 27972 26862
rect 27916 26798 27918 26850
rect 27970 26798 27972 26850
rect 27916 26740 27972 26798
rect 28364 26740 28420 27916
rect 28588 27860 28644 27916
rect 27916 26684 28364 26740
rect 28364 26646 28420 26684
rect 28476 27858 28644 27860
rect 28476 27806 28590 27858
rect 28642 27806 28644 27858
rect 28476 27804 28644 27806
rect 28028 26516 28084 26526
rect 28028 26422 28084 26460
rect 28476 26516 28532 27804
rect 28588 27794 28644 27804
rect 28700 27748 28756 27758
rect 28588 27076 28644 27086
rect 28588 26982 28644 27020
rect 28476 26450 28532 26460
rect 28700 26404 28756 27692
rect 28700 26338 28756 26348
rect 27804 26238 27806 26290
rect 27858 26238 27860 26290
rect 27804 26226 27860 26238
rect 28252 26292 28308 26302
rect 27916 25620 27972 25630
rect 27356 25452 27748 25508
rect 27020 25330 27076 25340
rect 26348 24782 26350 24834
rect 26402 24782 26404 24834
rect 26124 24724 26180 24734
rect 26124 24630 26180 24668
rect 26012 24558 26014 24610
rect 26066 24558 26068 24610
rect 26012 24546 26068 24558
rect 26348 23828 26404 24782
rect 26460 25282 26516 25294
rect 26460 25230 26462 25282
rect 26514 25230 26516 25282
rect 26460 24276 26516 25230
rect 26908 25284 26964 25294
rect 26908 25190 26964 25228
rect 27244 25284 27300 25294
rect 27580 25284 27636 25294
rect 27244 25282 27412 25284
rect 27244 25230 27246 25282
rect 27298 25230 27412 25282
rect 27244 25228 27412 25230
rect 27244 25218 27300 25228
rect 27132 25172 27188 25182
rect 26796 24722 26852 24734
rect 26796 24670 26798 24722
rect 26850 24670 26852 24722
rect 26796 24612 26852 24670
rect 27132 24724 27188 25116
rect 27132 24722 27300 24724
rect 27132 24670 27134 24722
rect 27186 24670 27300 24722
rect 27132 24668 27300 24670
rect 27132 24658 27188 24668
rect 26796 24546 26852 24556
rect 27132 24500 27188 24510
rect 26460 24210 26516 24220
rect 26908 24498 27188 24500
rect 26908 24446 27134 24498
rect 27186 24446 27188 24498
rect 26908 24444 27188 24446
rect 26684 24052 26740 24062
rect 26460 23940 26516 23950
rect 26684 23940 26740 23996
rect 26796 23940 26852 23950
rect 26684 23938 26852 23940
rect 26684 23886 26798 23938
rect 26850 23886 26852 23938
rect 26684 23884 26852 23886
rect 26460 23846 26516 23884
rect 26796 23874 26852 23884
rect 26348 23734 26404 23772
rect 26908 23548 26964 24444
rect 27132 24434 27188 24444
rect 27244 23940 27300 24668
rect 27356 24164 27412 25228
rect 27580 25190 27636 25228
rect 27468 25172 27524 25182
rect 27468 24834 27524 25116
rect 27468 24782 27470 24834
rect 27522 24782 27524 24834
rect 27468 24770 27524 24782
rect 27356 24098 27412 24108
rect 27468 23940 27524 23950
rect 27692 23940 27748 25452
rect 27916 25394 27972 25564
rect 28252 25506 28308 26236
rect 28364 26290 28420 26302
rect 28364 26238 28366 26290
rect 28418 26238 28420 26290
rect 28364 26180 28420 26238
rect 28364 25620 28420 26124
rect 28924 26180 28980 28924
rect 29260 28644 29316 28654
rect 29260 28550 29316 28588
rect 29372 27860 29428 30604
rect 29820 30210 29876 30940
rect 29820 30158 29822 30210
rect 29874 30158 29876 30210
rect 29820 30146 29876 30158
rect 30268 30098 30324 31724
rect 30268 30046 30270 30098
rect 30322 30046 30324 30098
rect 30268 30034 30324 30046
rect 30380 29540 30436 37214
rect 31276 37266 31332 37324
rect 31276 37214 31278 37266
rect 31330 37214 31332 37266
rect 31276 37202 31332 37214
rect 32172 37266 32228 37278
rect 32172 37214 32174 37266
rect 32226 37214 32228 37266
rect 30940 37156 30996 37166
rect 30604 36484 30660 36494
rect 30604 36390 30660 36428
rect 30940 35810 30996 37100
rect 31612 37156 31668 37166
rect 31612 37062 31668 37100
rect 31388 36482 31444 36494
rect 31388 36430 31390 36482
rect 31442 36430 31444 36482
rect 31388 35924 31444 36430
rect 31836 35924 31892 35934
rect 31388 35922 31892 35924
rect 31388 35870 31838 35922
rect 31890 35870 31892 35922
rect 31388 35868 31892 35870
rect 31836 35858 31892 35868
rect 30940 35758 30942 35810
rect 30994 35758 30996 35810
rect 30940 35746 30996 35758
rect 32060 33348 32116 33358
rect 32060 33254 32116 33292
rect 30716 32562 30772 32574
rect 30716 32510 30718 32562
rect 30770 32510 30772 32562
rect 30716 30882 30772 32510
rect 32060 31778 32116 31790
rect 32060 31726 32062 31778
rect 32114 31726 32116 31778
rect 30716 30830 30718 30882
rect 30770 30830 30772 30882
rect 30716 30818 30772 30830
rect 30828 31444 30884 31454
rect 30604 29988 30660 29998
rect 30604 29894 30660 29932
rect 30380 29474 30436 29484
rect 29932 29428 29988 29438
rect 29148 27636 29204 27646
rect 29148 27076 29204 27580
rect 29148 26962 29204 27020
rect 29372 27074 29428 27804
rect 29372 27022 29374 27074
rect 29426 27022 29428 27074
rect 29372 27010 29428 27022
rect 29708 28642 29764 28654
rect 29708 28590 29710 28642
rect 29762 28590 29764 28642
rect 29148 26910 29150 26962
rect 29202 26910 29204 26962
rect 29148 26898 29204 26910
rect 29708 26290 29764 28590
rect 29820 27972 29876 27982
rect 29820 27858 29876 27916
rect 29820 27806 29822 27858
rect 29874 27806 29876 27858
rect 29820 27794 29876 27806
rect 29708 26238 29710 26290
rect 29762 26238 29764 26290
rect 28924 26178 29092 26180
rect 28924 26126 28926 26178
rect 28978 26126 29092 26178
rect 28924 26124 29092 26126
rect 28924 26114 28980 26124
rect 28364 25554 28420 25564
rect 28252 25454 28254 25506
rect 28306 25454 28308 25506
rect 28252 25442 28308 25454
rect 27916 25342 27918 25394
rect 27970 25342 27972 25394
rect 27916 25330 27972 25342
rect 28364 25284 28420 25294
rect 27804 24052 27860 24062
rect 27804 23958 27860 23996
rect 28364 24050 28420 25228
rect 28588 25284 28644 25294
rect 28588 25190 28644 25228
rect 28364 23998 28366 24050
rect 28418 23998 28420 24050
rect 28364 23986 28420 23998
rect 27244 23938 27524 23940
rect 27244 23886 27470 23938
rect 27522 23886 27524 23938
rect 27244 23884 27524 23886
rect 27468 23874 27524 23884
rect 27580 23884 27748 23940
rect 29036 23940 29092 26124
rect 29260 26178 29316 26190
rect 29260 26126 29262 26178
rect 29314 26126 29316 26178
rect 29260 24834 29316 26126
rect 29260 24782 29262 24834
rect 29314 24782 29316 24834
rect 29260 24770 29316 24782
rect 29596 24724 29652 24734
rect 29596 24050 29652 24668
rect 29596 23998 29598 24050
rect 29650 23998 29652 24050
rect 29596 23986 29652 23998
rect 27132 23716 27188 23726
rect 26684 23492 26964 23548
rect 27020 23714 27188 23716
rect 27020 23662 27134 23714
rect 27186 23662 27188 23714
rect 27020 23660 27188 23662
rect 26460 23436 26740 23492
rect 25900 23324 26180 23380
rect 25788 23202 25844 23212
rect 25228 23102 25230 23154
rect 25282 23102 25284 23154
rect 25228 23090 25284 23102
rect 25900 23154 25956 23166
rect 25900 23102 25902 23154
rect 25954 23102 25956 23154
rect 25452 23044 25508 23054
rect 25340 22932 25396 22942
rect 25340 22258 25396 22876
rect 25340 22206 25342 22258
rect 25394 22206 25396 22258
rect 25340 22194 25396 22206
rect 25004 22146 25060 22158
rect 25004 22094 25006 22146
rect 25058 22094 25060 22146
rect 25004 22036 25060 22094
rect 25004 21970 25060 21980
rect 24892 21410 24948 21420
rect 24668 20524 24948 20580
rect 24332 20468 24388 20524
rect 24332 20412 24724 20468
rect 23772 20300 24276 20356
rect 24220 20244 24276 20300
rect 24444 20244 24500 20254
rect 24220 20242 24500 20244
rect 24220 20190 24446 20242
rect 24498 20190 24500 20242
rect 24220 20188 24500 20190
rect 24444 20178 24500 20188
rect 23772 20132 23828 20142
rect 23772 20038 23828 20076
rect 24108 20130 24164 20142
rect 24108 20078 24110 20130
rect 24162 20078 24164 20130
rect 23436 18398 23438 18450
rect 23490 18398 23492 18450
rect 23436 18386 23492 18398
rect 23548 18676 23604 18686
rect 23212 17574 23268 17612
rect 23436 17556 23492 17566
rect 22876 17554 23156 17556
rect 22876 17502 22878 17554
rect 22930 17502 23156 17554
rect 22876 17500 23156 17502
rect 22876 17490 22932 17500
rect 22540 17442 22596 17454
rect 22540 17390 22542 17442
rect 22594 17390 22596 17442
rect 22540 17332 22596 17390
rect 22540 17266 22596 17276
rect 22204 17052 23044 17108
rect 22652 16884 22708 16894
rect 22428 16324 22484 16334
rect 22428 15538 22484 16268
rect 22428 15486 22430 15538
rect 22482 15486 22484 15538
rect 22428 15474 22484 15486
rect 22652 15314 22708 16828
rect 22764 16882 22820 16894
rect 22764 16830 22766 16882
rect 22818 16830 22820 16882
rect 22764 15540 22820 16830
rect 22988 16770 23044 17052
rect 22988 16718 22990 16770
rect 23042 16718 23044 16770
rect 22988 16706 23044 16718
rect 23100 17106 23156 17500
rect 23100 17054 23102 17106
rect 23154 17054 23156 17106
rect 23100 16100 23156 17054
rect 23100 16034 23156 16044
rect 23324 16996 23380 17006
rect 23436 16996 23492 17500
rect 23324 16994 23492 16996
rect 23324 16942 23326 16994
rect 23378 16942 23492 16994
rect 23324 16940 23492 16942
rect 22764 15474 22820 15484
rect 23324 15538 23380 16940
rect 23324 15486 23326 15538
rect 23378 15486 23380 15538
rect 23324 15474 23380 15486
rect 22652 15262 22654 15314
rect 22706 15262 22708 15314
rect 22652 15250 22708 15262
rect 22316 15202 22372 15214
rect 22316 15150 22318 15202
rect 22370 15150 22372 15202
rect 22316 13858 22372 15150
rect 22316 13806 22318 13858
rect 22370 13806 22372 13858
rect 22316 13794 22372 13806
rect 22540 14980 22596 14990
rect 22204 13412 22260 13422
rect 22204 12404 22260 13356
rect 22204 12310 22260 12348
rect 22428 12852 22484 12862
rect 22092 8866 22148 8876
rect 22204 11060 22260 11070
rect 22204 10612 22260 11004
rect 21644 8206 21646 8258
rect 21698 8206 21700 8258
rect 21644 8194 21700 8206
rect 21980 8484 22036 8494
rect 20636 8036 20692 8046
rect 20636 7942 20692 7980
rect 21308 8034 21364 8046
rect 21308 7982 21310 8034
rect 21362 7982 21364 8034
rect 20412 7812 20468 7822
rect 20188 6524 20356 6580
rect 19852 6412 20244 6468
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20188 6132 20244 6412
rect 20188 6066 20244 6076
rect 19852 6020 19908 6030
rect 19852 5926 19908 5964
rect 20300 5236 20356 6524
rect 20300 5124 20356 5180
rect 20188 5068 20356 5124
rect 20412 5122 20468 7756
rect 21308 7812 21364 7982
rect 21308 7746 21364 7756
rect 21980 7698 22036 8428
rect 21980 7646 21982 7698
rect 22034 7646 22036 7698
rect 21980 7634 22036 7646
rect 21308 7586 21364 7598
rect 21308 7534 21310 7586
rect 21362 7534 21364 7586
rect 21308 7364 21364 7534
rect 21308 7298 21364 7308
rect 21420 7476 21476 7486
rect 20636 6580 20692 6590
rect 21308 6580 21364 6590
rect 20636 6578 21364 6580
rect 20636 6526 20638 6578
rect 20690 6526 21310 6578
rect 21362 6526 21364 6578
rect 20636 6524 21364 6526
rect 20636 6514 20692 6524
rect 21308 6514 21364 6524
rect 20412 5070 20414 5122
rect 20466 5070 20468 5122
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 4510 19630 4562
rect 19682 4510 19684 4562
rect 19628 4498 19684 4510
rect 19740 4564 19796 4574
rect 20188 4564 20244 5068
rect 20412 5058 20468 5070
rect 20524 6468 20580 6478
rect 19180 4398 19182 4450
rect 19234 4398 19236 4450
rect 19180 4386 19236 4398
rect 19740 4338 19796 4508
rect 19740 4286 19742 4338
rect 19794 4286 19796 4338
rect 19740 4274 19796 4286
rect 19852 4508 20244 4564
rect 18620 4050 18676 4060
rect 19516 4116 19572 4126
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 19516 3442 19572 4060
rect 19852 3554 19908 4508
rect 20524 4452 20580 6412
rect 21420 6356 21476 7420
rect 20748 6300 21476 6356
rect 21532 7364 21588 7374
rect 20748 5010 20804 6300
rect 20972 6132 21028 6142
rect 20748 4958 20750 5010
rect 20802 4958 20804 5010
rect 20748 4946 20804 4958
rect 20860 5796 20916 5806
rect 20636 4452 20692 4462
rect 20524 4450 20692 4452
rect 20524 4398 20638 4450
rect 20690 4398 20692 4450
rect 20524 4396 20692 4398
rect 20636 4386 20692 4396
rect 20300 4338 20356 4350
rect 20300 4286 20302 4338
rect 20354 4286 20356 4338
rect 20300 4228 20356 4286
rect 20860 4228 20916 5740
rect 20972 4450 21028 6076
rect 21308 6020 21364 6030
rect 21532 6020 21588 7308
rect 21644 7364 21700 7374
rect 21644 7362 21812 7364
rect 21644 7310 21646 7362
rect 21698 7310 21812 7362
rect 21644 7308 21812 7310
rect 21644 7298 21700 7308
rect 21364 5964 21588 6020
rect 21644 6692 21700 6702
rect 21756 6692 21812 7308
rect 22092 6692 22148 6702
rect 21756 6690 22148 6692
rect 21756 6638 22094 6690
rect 22146 6638 22148 6690
rect 21756 6636 22148 6638
rect 21196 5908 21252 5918
rect 21196 5814 21252 5852
rect 20972 4398 20974 4450
rect 21026 4398 21028 4450
rect 20972 4386 21028 4398
rect 21308 4340 21364 5964
rect 21644 5908 21700 6636
rect 22092 6626 22148 6636
rect 22204 6468 22260 10556
rect 22316 8146 22372 8158
rect 22316 8094 22318 8146
rect 22370 8094 22372 8146
rect 22316 6578 22372 8094
rect 22316 6526 22318 6578
rect 22370 6526 22372 6578
rect 22316 6514 22372 6526
rect 22428 7362 22484 12796
rect 22540 12290 22596 14924
rect 23324 12850 23380 12862
rect 23324 12798 23326 12850
rect 23378 12798 23380 12850
rect 22540 12238 22542 12290
rect 22594 12238 22596 12290
rect 22540 12226 22596 12238
rect 22876 12290 22932 12302
rect 22876 12238 22878 12290
rect 22930 12238 22932 12290
rect 22652 11396 22708 11406
rect 22876 11396 22932 12238
rect 23212 12290 23268 12302
rect 23212 12238 23214 12290
rect 23266 12238 23268 12290
rect 23100 11396 23156 11406
rect 22652 11394 22932 11396
rect 22652 11342 22654 11394
rect 22706 11342 22932 11394
rect 22652 11340 22932 11342
rect 22988 11340 23100 11396
rect 22652 11172 22708 11340
rect 22652 11106 22708 11116
rect 22428 7310 22430 7362
rect 22482 7310 22484 7362
rect 22092 6412 22260 6468
rect 21756 5908 21812 5918
rect 21644 5906 21812 5908
rect 21644 5854 21758 5906
rect 21810 5854 21812 5906
rect 21644 5852 21812 5854
rect 21420 5796 21476 5806
rect 21756 5796 21812 5852
rect 21420 5794 21700 5796
rect 21420 5742 21422 5794
rect 21474 5742 21700 5794
rect 21420 5740 21700 5742
rect 21420 5730 21476 5740
rect 21420 5236 21476 5246
rect 21420 5142 21476 5180
rect 21532 5124 21588 5134
rect 21532 5030 21588 5068
rect 21644 5012 21700 5740
rect 21756 5730 21812 5740
rect 22092 5684 22148 6412
rect 22428 6356 22484 7310
rect 22316 6300 22484 6356
rect 22540 10722 22596 10734
rect 22540 10670 22542 10722
rect 22594 10670 22596 10722
rect 22204 5908 22260 5918
rect 22204 5814 22260 5852
rect 22092 5618 22148 5628
rect 22316 5012 22372 6300
rect 22540 6244 22596 10670
rect 22988 9826 23044 11340
rect 23100 11302 23156 11340
rect 23212 11060 23268 12238
rect 23212 10994 23268 11004
rect 23324 12292 23380 12798
rect 23324 10836 23380 12236
rect 23436 12740 23492 12750
rect 23436 12178 23492 12684
rect 23548 12628 23604 18620
rect 24108 18564 24164 20078
rect 24556 19908 24612 19918
rect 24556 19814 24612 19852
rect 24668 19348 24724 20412
rect 24780 19348 24836 19358
rect 24668 19292 24780 19348
rect 24780 19282 24836 19292
rect 23884 18452 23940 18462
rect 23772 18226 23828 18238
rect 23772 18174 23774 18226
rect 23826 18174 23828 18226
rect 23772 17890 23828 18174
rect 23772 17838 23774 17890
rect 23826 17838 23828 17890
rect 23772 17826 23828 17838
rect 23884 17106 23940 18396
rect 23884 17054 23886 17106
rect 23938 17054 23940 17106
rect 23884 16884 23940 17054
rect 23884 16818 23940 16828
rect 23772 16772 23828 16782
rect 23772 16678 23828 16716
rect 23660 16658 23716 16670
rect 23660 16606 23662 16658
rect 23714 16606 23716 16658
rect 23660 16210 23716 16606
rect 23660 16158 23662 16210
rect 23714 16158 23716 16210
rect 23660 16146 23716 16158
rect 23660 15652 23716 15662
rect 23660 15314 23716 15596
rect 24108 15538 24164 18508
rect 24556 19122 24612 19134
rect 24556 19070 24558 19122
rect 24610 19070 24612 19122
rect 24556 18562 24612 19070
rect 24556 18510 24558 18562
rect 24610 18510 24612 18562
rect 24556 18498 24612 18510
rect 24220 18452 24276 18462
rect 24220 18358 24276 18396
rect 24668 18116 24724 18126
rect 24668 17108 24724 18060
rect 24668 17014 24724 17052
rect 24108 15486 24110 15538
rect 24162 15486 24164 15538
rect 24108 15474 24164 15486
rect 24332 15876 24388 15886
rect 23660 15262 23662 15314
rect 23714 15262 23716 15314
rect 23660 14642 23716 15262
rect 24332 15428 24388 15820
rect 24332 15148 24388 15372
rect 24668 15202 24724 15214
rect 24668 15150 24670 15202
rect 24722 15150 24724 15202
rect 24668 15148 24724 15150
rect 24332 15092 24612 15148
rect 24668 15092 24836 15148
rect 24220 14868 24276 14878
rect 23660 14590 23662 14642
rect 23714 14590 23716 14642
rect 23660 14578 23716 14590
rect 24108 14644 24164 14654
rect 24108 14550 24164 14588
rect 24108 13972 24164 13982
rect 24220 13972 24276 14812
rect 24556 14644 24612 15092
rect 24668 14644 24724 14654
rect 24556 14642 24724 14644
rect 24556 14590 24670 14642
rect 24722 14590 24724 14642
rect 24556 14588 24724 14590
rect 24668 14578 24724 14588
rect 24780 14532 24836 15092
rect 24892 14868 24948 20524
rect 25452 20020 25508 22988
rect 25788 23042 25844 23054
rect 25788 22990 25790 23042
rect 25842 22990 25844 23042
rect 25788 21700 25844 22990
rect 25900 22482 25956 23102
rect 26124 23044 26180 23324
rect 26460 23378 26516 23436
rect 26460 23326 26462 23378
rect 26514 23326 26516 23378
rect 26460 23314 26516 23326
rect 26124 22978 26180 22988
rect 26236 23154 26292 23166
rect 26796 23156 26852 23166
rect 26236 23102 26238 23154
rect 26290 23102 26292 23154
rect 25900 22430 25902 22482
rect 25954 22430 25956 22482
rect 25900 22418 25956 22430
rect 26012 22932 26068 22942
rect 25900 22146 25956 22158
rect 25900 22094 25902 22146
rect 25954 22094 25956 22146
rect 25900 21812 25956 22094
rect 26012 21812 26068 22876
rect 26236 22372 26292 23102
rect 26684 23154 26852 23156
rect 26684 23102 26798 23154
rect 26850 23102 26852 23154
rect 26684 23100 26852 23102
rect 26348 23044 26404 23054
rect 26684 23044 26740 23100
rect 26796 23090 26852 23100
rect 26348 23042 26628 23044
rect 26348 22990 26350 23042
rect 26402 22990 26628 23042
rect 26348 22988 26628 22990
rect 26348 22978 26404 22988
rect 26236 22316 26404 22372
rect 26124 22258 26180 22270
rect 26124 22206 26126 22258
rect 26178 22206 26180 22258
rect 26124 22036 26180 22206
rect 26124 21970 26180 21980
rect 26124 21812 26180 21822
rect 25900 21810 26180 21812
rect 25900 21758 26126 21810
rect 26178 21758 26180 21810
rect 25900 21756 26180 21758
rect 25788 21634 25844 21644
rect 26124 20804 26180 21756
rect 26236 21812 26292 21822
rect 26348 21812 26404 22316
rect 26236 21810 26404 21812
rect 26236 21758 26238 21810
rect 26290 21758 26404 21810
rect 26236 21756 26404 21758
rect 26236 21746 26292 21756
rect 26348 21364 26404 21374
rect 26348 21362 26516 21364
rect 26348 21310 26350 21362
rect 26402 21310 26516 21362
rect 26348 21308 26516 21310
rect 26348 21298 26404 21308
rect 26124 20738 26180 20748
rect 25452 19954 25508 19964
rect 26124 19908 26180 19918
rect 25340 18340 25396 18350
rect 25340 18246 25396 18284
rect 25004 17668 25060 17678
rect 25004 16098 25060 17612
rect 26124 16882 26180 19852
rect 26124 16830 26126 16882
rect 26178 16830 26180 16882
rect 26124 16818 26180 16830
rect 26236 18340 26292 18350
rect 26236 16884 26292 18284
rect 26348 16884 26404 16894
rect 26236 16882 26404 16884
rect 26236 16830 26350 16882
rect 26402 16830 26404 16882
rect 26236 16828 26404 16830
rect 25676 16660 25732 16670
rect 25900 16660 25956 16670
rect 25676 16566 25732 16604
rect 25788 16658 25956 16660
rect 25788 16606 25902 16658
rect 25954 16606 25956 16658
rect 25788 16604 25956 16606
rect 25788 16324 25844 16604
rect 25900 16594 25956 16604
rect 26012 16660 26068 16670
rect 26236 16660 26292 16670
rect 25452 16268 25844 16324
rect 25452 16210 25508 16268
rect 25452 16158 25454 16210
rect 25506 16158 25508 16210
rect 25452 16146 25508 16158
rect 25004 16046 25006 16098
rect 25058 16046 25060 16098
rect 25004 16034 25060 16046
rect 25340 15986 25396 15998
rect 25340 15934 25342 15986
rect 25394 15934 25396 15986
rect 24892 14802 24948 14812
rect 25116 15652 25172 15662
rect 25004 14644 25060 14654
rect 25004 14550 25060 14588
rect 24780 14466 24836 14476
rect 23884 13970 24276 13972
rect 23884 13918 24110 13970
rect 24162 13918 24276 13970
rect 23884 13916 24276 13918
rect 23884 12962 23940 13916
rect 24108 13906 24164 13916
rect 25116 13412 25172 15596
rect 25228 15316 25284 15326
rect 25228 15222 25284 15260
rect 25340 14642 25396 15934
rect 25564 15538 25620 16268
rect 25564 15486 25566 15538
rect 25618 15486 25620 15538
rect 25564 15474 25620 15486
rect 25900 16098 25956 16110
rect 25900 16046 25902 16098
rect 25954 16046 25956 16098
rect 25900 15314 25956 16046
rect 26012 16098 26068 16604
rect 26012 16046 26014 16098
rect 26066 16046 26068 16098
rect 26012 15428 26068 16046
rect 26012 15334 26068 15372
rect 26124 16658 26292 16660
rect 26124 16606 26238 16658
rect 26290 16606 26292 16658
rect 26124 16604 26292 16606
rect 25900 15262 25902 15314
rect 25954 15262 25956 15314
rect 25340 14590 25342 14642
rect 25394 14590 25396 14642
rect 25340 14578 25396 14590
rect 25452 14756 25508 14766
rect 25452 13972 25508 14700
rect 25900 14644 25956 15262
rect 25900 14578 25956 14588
rect 26012 15204 26068 15214
rect 25788 14532 25844 14542
rect 25452 13970 25732 13972
rect 25452 13918 25454 13970
rect 25506 13918 25732 13970
rect 25452 13916 25732 13918
rect 25452 13906 25508 13916
rect 25676 13858 25732 13916
rect 25676 13806 25678 13858
rect 25730 13806 25732 13858
rect 25676 13794 25732 13806
rect 25116 13356 25620 13412
rect 23884 12910 23886 12962
rect 23938 12910 23940 12962
rect 23884 12898 23940 12910
rect 23996 12964 24052 12974
rect 23548 12572 23716 12628
rect 23436 12126 23438 12178
rect 23490 12126 23492 12178
rect 23436 12114 23492 12126
rect 22988 9774 22990 9826
rect 23042 9774 23044 9826
rect 22988 9762 23044 9774
rect 23100 10780 23380 10836
rect 23660 10834 23716 12572
rect 23660 10782 23662 10834
rect 23714 10782 23716 10834
rect 23100 10722 23156 10780
rect 23660 10770 23716 10782
rect 23884 12068 23940 12078
rect 23996 12068 24052 12908
rect 24444 12964 24500 12974
rect 24444 12962 24948 12964
rect 24444 12910 24446 12962
rect 24498 12910 24948 12962
rect 24444 12908 24948 12910
rect 24444 12898 24500 12908
rect 24556 12738 24612 12750
rect 24556 12686 24558 12738
rect 24610 12686 24612 12738
rect 24556 12404 24612 12686
rect 23884 12066 24052 12068
rect 23884 12014 23886 12066
rect 23938 12014 24052 12066
rect 23884 12012 24052 12014
rect 24220 12348 24612 12404
rect 24780 12738 24836 12750
rect 24780 12686 24782 12738
rect 24834 12686 24836 12738
rect 23884 11394 23940 12012
rect 23884 11342 23886 11394
rect 23938 11342 23940 11394
rect 23100 10670 23102 10722
rect 23154 10670 23156 10722
rect 23100 9604 23156 10670
rect 23884 10612 23940 11342
rect 24220 11396 24276 12348
rect 24332 12180 24388 12190
rect 24332 12086 24388 12124
rect 24556 12068 24612 12078
rect 24276 11340 24388 11396
rect 24220 11302 24276 11340
rect 24332 10836 24388 11340
rect 24444 10836 24500 10846
rect 24332 10834 24500 10836
rect 24332 10782 24446 10834
rect 24498 10782 24500 10834
rect 24332 10780 24500 10782
rect 24444 10770 24500 10780
rect 24556 10834 24612 12012
rect 24556 10782 24558 10834
rect 24610 10782 24612 10834
rect 24556 10770 24612 10782
rect 24668 11508 24724 11518
rect 24668 10834 24724 11452
rect 24668 10782 24670 10834
rect 24722 10782 24724 10834
rect 23996 10612 24052 10622
rect 23884 10610 24052 10612
rect 23884 10558 23998 10610
rect 24050 10558 24052 10610
rect 23884 10556 24052 10558
rect 23324 10386 23380 10398
rect 23324 10334 23326 10386
rect 23378 10334 23380 10386
rect 22764 9548 23156 9604
rect 23212 10052 23268 10062
rect 22764 8146 22820 9548
rect 23212 9492 23268 9996
rect 23324 9716 23380 10334
rect 23996 9940 24052 10556
rect 23996 9874 24052 9884
rect 24108 10164 24164 10174
rect 23324 9650 23380 9660
rect 23548 9716 23604 9726
rect 23996 9716 24052 9726
rect 23548 9714 24052 9716
rect 23548 9662 23550 9714
rect 23602 9662 23998 9714
rect 24050 9662 24052 9714
rect 23548 9660 24052 9662
rect 23548 9650 23604 9660
rect 23996 9650 24052 9660
rect 23212 9436 23716 9492
rect 23324 9156 23380 9166
rect 23324 9154 23492 9156
rect 23324 9102 23326 9154
rect 23378 9102 23492 9154
rect 23324 9100 23492 9102
rect 23324 9090 23380 9100
rect 22988 9042 23044 9054
rect 22988 8990 22990 9042
rect 23042 8990 23044 9042
rect 22988 8708 23044 8990
rect 22764 8094 22766 8146
rect 22818 8094 22820 8146
rect 22764 8082 22820 8094
rect 22876 8652 23044 8708
rect 23324 8932 23380 8942
rect 22876 7476 22932 8652
rect 23324 8370 23380 8876
rect 23324 8318 23326 8370
rect 23378 8318 23380 8370
rect 23324 8306 23380 8318
rect 22988 8258 23044 8270
rect 22988 8206 22990 8258
rect 23042 8206 23044 8258
rect 22988 7700 23044 8206
rect 22988 7634 23044 7644
rect 23436 7588 23492 9100
rect 23660 9042 23716 9436
rect 23660 8990 23662 9042
rect 23714 8990 23716 9042
rect 23660 8978 23716 8990
rect 24108 9042 24164 10108
rect 24668 10052 24724 10782
rect 24668 9986 24724 9996
rect 24108 8990 24110 9042
rect 24162 8990 24164 9042
rect 24108 8978 24164 8990
rect 24444 9826 24500 9838
rect 24444 9774 24446 9826
rect 24498 9774 24500 9826
rect 24444 8596 24500 9774
rect 24780 9826 24836 12686
rect 24780 9774 24782 9826
rect 24834 9774 24836 9826
rect 24780 9762 24836 9774
rect 24892 8932 24948 12908
rect 25564 12850 25620 13356
rect 25564 12798 25566 12850
rect 25618 12798 25620 12850
rect 25564 12786 25620 12798
rect 25228 12740 25284 12750
rect 25228 12646 25284 12684
rect 25564 12180 25620 12190
rect 25788 12180 25844 14476
rect 26012 14084 26068 15148
rect 26124 14530 26180 16604
rect 26236 16594 26292 16604
rect 26348 15316 26404 16828
rect 26348 15250 26404 15260
rect 26124 14478 26126 14530
rect 26178 14478 26180 14530
rect 26124 14466 26180 14478
rect 26348 14420 26404 14430
rect 26460 14420 26516 21308
rect 26572 21252 26628 22988
rect 26684 22372 26740 22988
rect 26796 22932 26852 22942
rect 26796 22596 26852 22876
rect 27020 22596 27076 23660
rect 27132 23650 27188 23660
rect 27244 23380 27300 23390
rect 27244 23154 27300 23324
rect 27468 23380 27524 23390
rect 27580 23380 27636 23884
rect 29036 23874 29092 23884
rect 27692 23716 27748 23726
rect 27692 23622 27748 23660
rect 29372 23716 29428 23726
rect 27916 23380 27972 23390
rect 27468 23378 27860 23380
rect 27468 23326 27470 23378
rect 27522 23326 27860 23378
rect 27468 23324 27860 23326
rect 27468 23314 27524 23324
rect 27244 23102 27246 23154
rect 27298 23102 27300 23154
rect 27244 22820 27300 23102
rect 27244 22754 27300 22764
rect 26796 22540 27076 22596
rect 27804 22484 27860 23324
rect 27916 23286 27972 23324
rect 29372 23380 29428 23660
rect 29372 23314 29428 23324
rect 29036 23266 29092 23278
rect 29036 23214 29038 23266
rect 29090 23214 29092 23266
rect 28700 23154 28756 23166
rect 28700 23102 28702 23154
rect 28754 23102 28756 23154
rect 28364 23044 28420 23054
rect 28700 23044 28756 23102
rect 28364 23042 28756 23044
rect 28364 22990 28366 23042
rect 28418 22990 28756 23042
rect 28364 22988 28756 22990
rect 28364 22596 28420 22988
rect 28364 22530 28420 22540
rect 27804 22428 28308 22484
rect 26908 22372 26964 22382
rect 26684 22370 26852 22372
rect 26684 22318 26686 22370
rect 26738 22318 26852 22370
rect 26684 22316 26852 22318
rect 26684 22306 26740 22316
rect 26572 21186 26628 21196
rect 26684 22036 26740 22046
rect 26572 16658 26628 16670
rect 26572 16606 26574 16658
rect 26626 16606 26628 16658
rect 26572 16212 26628 16606
rect 26572 15876 26628 16156
rect 26572 15810 26628 15820
rect 26684 15148 26740 21980
rect 26796 21810 26852 22316
rect 26796 21758 26798 21810
rect 26850 21758 26852 21810
rect 26796 21746 26852 21758
rect 26908 21252 26964 22316
rect 27020 22372 27076 22382
rect 27580 22372 27636 22382
rect 27020 22370 27524 22372
rect 27020 22318 27022 22370
rect 27074 22318 27524 22370
rect 27020 22316 27524 22318
rect 27020 22306 27076 22316
rect 27132 22146 27188 22158
rect 27132 22094 27134 22146
rect 27186 22094 27188 22146
rect 27132 21812 27188 22094
rect 27244 22148 27300 22158
rect 27244 22146 27412 22148
rect 27244 22094 27246 22146
rect 27298 22094 27412 22146
rect 27244 22092 27412 22094
rect 27244 22082 27300 22092
rect 27132 21746 27188 21756
rect 27356 21700 27412 22092
rect 27468 21924 27524 22316
rect 27580 22278 27636 22316
rect 27468 21868 27748 21924
rect 27356 21644 27524 21700
rect 27020 21586 27076 21598
rect 27020 21534 27022 21586
rect 27074 21534 27076 21586
rect 27020 21476 27076 21534
rect 27244 21588 27300 21598
rect 27244 21494 27300 21532
rect 27020 21410 27076 21420
rect 27132 21474 27188 21486
rect 27132 21422 27134 21474
rect 27186 21422 27188 21474
rect 27132 21252 27188 21422
rect 26908 21196 27188 21252
rect 27244 21140 27300 21150
rect 26796 20804 26852 20814
rect 27132 20804 27188 20814
rect 26852 20748 27132 20804
rect 26796 20738 26852 20748
rect 27132 20710 27188 20748
rect 27244 20356 27300 21084
rect 27356 20916 27412 20926
rect 27468 20916 27524 21644
rect 27692 21474 27748 21868
rect 27804 21810 27860 22428
rect 28252 22372 28308 22428
rect 29036 22372 29092 23214
rect 29484 22930 29540 22942
rect 29484 22878 29486 22930
rect 29538 22878 29540 22930
rect 28252 22316 28532 22372
rect 27916 22260 27972 22270
rect 27916 22166 27972 22204
rect 27804 21758 27806 21810
rect 27858 21758 27860 21810
rect 27804 21746 27860 21758
rect 28252 22146 28308 22158
rect 28252 22094 28254 22146
rect 28306 22094 28308 22146
rect 28028 21700 28084 21710
rect 28028 21606 28084 21644
rect 27692 21422 27694 21474
rect 27746 21422 27748 21474
rect 27692 21410 27748 21422
rect 27804 21588 27860 21598
rect 27804 21026 27860 21532
rect 27804 20974 27806 21026
rect 27858 20974 27860 21026
rect 27804 20962 27860 20974
rect 28252 21252 28308 22094
rect 28476 21810 28532 22316
rect 28588 22146 28644 22158
rect 28588 22094 28590 22146
rect 28642 22094 28644 22146
rect 28588 21924 28644 22094
rect 29036 22036 29092 22316
rect 29260 22372 29316 22382
rect 29260 22278 29316 22316
rect 29036 21970 29092 21980
rect 29148 22260 29204 22270
rect 28588 21858 28644 21868
rect 28476 21758 28478 21810
rect 28530 21758 28532 21810
rect 28476 21746 28532 21758
rect 28588 21588 28644 21598
rect 28364 21476 28420 21486
rect 28364 21382 28420 21420
rect 28364 21252 28420 21262
rect 28252 21196 28364 21252
rect 27356 20914 27524 20916
rect 27356 20862 27358 20914
rect 27410 20862 27524 20914
rect 27356 20860 27524 20862
rect 27356 20850 27412 20860
rect 27804 20804 27860 20814
rect 27804 20710 27860 20748
rect 27132 20300 27300 20356
rect 27468 20690 27524 20702
rect 27468 20638 27470 20690
rect 27522 20638 27524 20690
rect 26796 17108 26852 17118
rect 26796 16770 26852 17052
rect 26796 16718 26798 16770
rect 26850 16718 26852 16770
rect 26796 16706 26852 16718
rect 26908 16436 26964 16446
rect 26908 16098 26964 16380
rect 26908 16046 26910 16098
rect 26962 16046 26964 16098
rect 26908 16034 26964 16046
rect 27132 15148 27188 20300
rect 27468 20244 27524 20638
rect 27468 20178 27524 20188
rect 28140 20690 28196 20702
rect 28140 20638 28142 20690
rect 28194 20638 28196 20690
rect 27244 16770 27300 16782
rect 27244 16718 27246 16770
rect 27298 16718 27300 16770
rect 27244 16436 27300 16718
rect 27244 16370 27300 16380
rect 27468 16772 27524 16782
rect 27356 16098 27412 16110
rect 27356 16046 27358 16098
rect 27410 16046 27412 16098
rect 27356 15428 27412 16046
rect 27356 15362 27412 15372
rect 26348 14418 26516 14420
rect 26348 14366 26350 14418
rect 26402 14366 26516 14418
rect 26348 14364 26516 14366
rect 26572 15092 26740 15148
rect 27020 15092 27188 15148
rect 26348 14354 26404 14364
rect 26012 14028 26180 14084
rect 26012 13858 26068 13870
rect 26012 13806 26014 13858
rect 26066 13806 26068 13858
rect 26012 13748 26068 13806
rect 26012 12740 26068 13692
rect 26124 13188 26180 14028
rect 26348 13860 26404 13870
rect 26348 13766 26404 13804
rect 26572 13412 26628 15092
rect 26796 14418 26852 14430
rect 26796 14366 26798 14418
rect 26850 14366 26852 14418
rect 26796 13860 26852 14366
rect 26684 13748 26740 13758
rect 26684 13654 26740 13692
rect 26124 13122 26180 13132
rect 26236 13356 26628 13412
rect 26012 12674 26068 12684
rect 26236 12402 26292 13356
rect 26236 12350 26238 12402
rect 26290 12350 26292 12402
rect 26236 12338 26292 12350
rect 26348 13188 26404 13198
rect 26348 12404 26404 13132
rect 26460 12964 26516 12974
rect 26460 12870 26516 12908
rect 25564 12178 25844 12180
rect 25564 12126 25566 12178
rect 25618 12126 25844 12178
rect 25564 12124 25844 12126
rect 26124 12178 26180 12190
rect 26124 12126 26126 12178
rect 26178 12126 26180 12178
rect 25228 12068 25284 12078
rect 25228 11974 25284 12012
rect 25004 9716 25060 9726
rect 25004 9622 25060 9660
rect 25452 9714 25508 9726
rect 25452 9662 25454 9714
rect 25506 9662 25508 9714
rect 25228 9044 25284 9054
rect 25228 8950 25284 8988
rect 25004 8932 25060 8942
rect 24892 8876 25004 8932
rect 24556 8596 24612 8606
rect 24444 8540 24556 8596
rect 24556 8530 24612 8540
rect 24220 8372 24276 8382
rect 24108 8316 24220 8372
rect 23884 8036 23940 8046
rect 23884 7942 23940 7980
rect 22876 7382 22932 7420
rect 23324 7532 23492 7588
rect 23324 6916 23380 7532
rect 24108 7474 24164 8316
rect 24220 8306 24276 8316
rect 24892 8372 24948 8382
rect 24892 8258 24948 8316
rect 24892 8206 24894 8258
rect 24946 8206 24948 8258
rect 24892 8194 24948 8206
rect 24668 8146 24724 8158
rect 24668 8094 24670 8146
rect 24722 8094 24724 8146
rect 24220 8036 24276 8046
rect 24220 8034 24612 8036
rect 24220 7982 24222 8034
rect 24274 7982 24612 8034
rect 24220 7980 24612 7982
rect 24220 7970 24276 7980
rect 24108 7422 24110 7474
rect 24162 7422 24164 7474
rect 23436 7364 23492 7374
rect 23492 7308 23604 7364
rect 23436 7270 23492 7308
rect 23324 6860 23492 6916
rect 22428 6188 22596 6244
rect 22876 6690 22932 6702
rect 23324 6692 23380 6702
rect 22876 6638 22878 6690
rect 22930 6638 22932 6690
rect 22428 6130 22484 6188
rect 22428 6078 22430 6130
rect 22482 6078 22484 6130
rect 22428 6066 22484 6078
rect 22876 5906 22932 6638
rect 22876 5854 22878 5906
rect 22930 5854 22932 5906
rect 22876 5684 22932 5854
rect 22876 5618 22932 5628
rect 22988 6690 23380 6692
rect 22988 6638 23326 6690
rect 23378 6638 23380 6690
rect 22988 6636 23380 6638
rect 22988 5234 23044 6636
rect 23324 6626 23380 6636
rect 22988 5182 22990 5234
rect 23042 5182 23044 5234
rect 22988 5170 23044 5182
rect 23436 5796 23492 6860
rect 21644 4956 22148 5012
rect 21644 4788 21700 4798
rect 21420 4340 21476 4350
rect 21308 4338 21476 4340
rect 21308 4286 21422 4338
rect 21474 4286 21476 4338
rect 21308 4284 21476 4286
rect 21420 4274 21476 4284
rect 21644 4338 21700 4732
rect 22092 4562 22148 4956
rect 22316 4946 22372 4956
rect 23100 5012 23156 5022
rect 22092 4510 22094 4562
rect 22146 4510 22148 4562
rect 22092 4498 22148 4510
rect 23100 4450 23156 4956
rect 23100 4398 23102 4450
rect 23154 4398 23156 4450
rect 23100 4386 23156 4398
rect 21644 4286 21646 4338
rect 21698 4286 21700 4338
rect 21644 4274 21700 4286
rect 23436 4340 23492 5740
rect 23548 5122 23604 7308
rect 23548 5070 23550 5122
rect 23602 5070 23604 5122
rect 23548 5058 23604 5070
rect 23660 5906 23716 5918
rect 23660 5854 23662 5906
rect 23714 5854 23716 5906
rect 23660 4562 23716 5854
rect 24108 5684 24164 7422
rect 24556 6804 24612 7980
rect 24668 7812 24724 8094
rect 24668 7746 24724 7756
rect 24668 7474 24724 7486
rect 24668 7422 24670 7474
rect 24722 7422 24724 7474
rect 24668 7364 24724 7422
rect 25004 7364 25060 8876
rect 25452 8260 25508 9662
rect 25564 8596 25620 12124
rect 26012 11508 26068 11518
rect 26012 11394 26068 11452
rect 26124 11506 26180 12126
rect 26124 11454 26126 11506
rect 26178 11454 26180 11506
rect 26124 11442 26180 11454
rect 26012 11342 26014 11394
rect 26066 11342 26068 11394
rect 26012 11330 26068 11342
rect 26348 11394 26404 12348
rect 26348 11342 26350 11394
rect 26402 11342 26404 11394
rect 26348 11330 26404 11342
rect 26796 12178 26852 13804
rect 26908 12964 26964 12974
rect 26908 12870 26964 12908
rect 27020 12404 27076 15092
rect 27468 13858 27524 16716
rect 28028 16324 28084 16334
rect 27580 16212 27636 16222
rect 27580 15314 27636 16156
rect 28028 16098 28084 16268
rect 28028 16046 28030 16098
rect 28082 16046 28084 16098
rect 28028 16034 28084 16046
rect 27580 15262 27582 15314
rect 27634 15262 27636 15314
rect 27580 15250 27636 15262
rect 27692 15426 27748 15438
rect 27692 15374 27694 15426
rect 27746 15374 27748 15426
rect 27580 14532 27636 14542
rect 27692 14532 27748 15374
rect 28140 15148 28196 20638
rect 28252 17556 28308 21196
rect 28364 21186 28420 21196
rect 28588 20914 28644 21532
rect 28700 21364 28756 21374
rect 28700 21270 28756 21308
rect 28588 20862 28590 20914
rect 28642 20862 28644 20914
rect 28588 20804 28644 20862
rect 28588 20738 28644 20748
rect 28700 20356 28756 20366
rect 28700 20130 28756 20300
rect 28700 20078 28702 20130
rect 28754 20078 28756 20130
rect 28700 20066 28756 20078
rect 28252 17462 28308 17500
rect 28364 20018 28420 20030
rect 28364 19966 28366 20018
rect 28418 19966 28420 20018
rect 28364 17108 28420 19966
rect 29148 19796 29204 22204
rect 29484 22036 29540 22878
rect 29260 21980 29540 22036
rect 29260 21698 29316 21980
rect 29260 21646 29262 21698
rect 29314 21646 29316 21698
rect 29260 21634 29316 21646
rect 29596 21924 29652 21934
rect 29260 20804 29316 20814
rect 29260 20710 29316 20748
rect 29260 20356 29316 20366
rect 29260 20018 29316 20300
rect 29596 20130 29652 21868
rect 29708 21586 29764 26238
rect 29820 27076 29876 27086
rect 29820 23938 29876 27020
rect 29932 27074 29988 29372
rect 30156 29202 30212 29214
rect 30156 29150 30158 29202
rect 30210 29150 30212 29202
rect 30156 28642 30212 29150
rect 30156 28590 30158 28642
rect 30210 28590 30212 28642
rect 30156 28578 30212 28590
rect 30492 28644 30548 28654
rect 30268 28418 30324 28430
rect 30268 28366 30270 28418
rect 30322 28366 30324 28418
rect 29932 27022 29934 27074
rect 29986 27022 29988 27074
rect 29932 26628 29988 27022
rect 29932 26562 29988 26572
rect 30044 27748 30100 27758
rect 30044 25506 30100 27692
rect 30268 27188 30324 28366
rect 30268 27122 30324 27132
rect 30380 27188 30436 27198
rect 30492 27188 30548 28588
rect 30828 28642 30884 31388
rect 32060 29540 32116 31726
rect 32060 29474 32116 29484
rect 31500 29426 31556 29438
rect 31500 29374 31502 29426
rect 31554 29374 31556 29426
rect 31164 29314 31220 29326
rect 31164 29262 31166 29314
rect 31218 29262 31220 29314
rect 31164 28980 31220 29262
rect 31164 28914 31220 28924
rect 31276 29202 31332 29214
rect 31276 29150 31278 29202
rect 31330 29150 31332 29202
rect 30828 28590 30830 28642
rect 30882 28590 30884 28642
rect 30828 28578 30884 28590
rect 31276 28642 31332 29150
rect 31276 28590 31278 28642
rect 31330 28590 31332 28642
rect 31276 28578 31332 28590
rect 31500 27748 31556 29374
rect 31836 29426 31892 29438
rect 31836 29374 31838 29426
rect 31890 29374 31892 29426
rect 31836 28644 31892 29374
rect 31836 28578 31892 28588
rect 32172 28196 32228 37214
rect 32284 37156 32340 38556
rect 32508 38836 32564 38894
rect 32508 38050 32564 38780
rect 33068 38834 33124 39228
rect 33068 38782 33070 38834
rect 33122 38782 33124 38834
rect 33068 38770 33124 38782
rect 33516 38836 33572 38846
rect 33516 38742 33572 38780
rect 33628 38668 33684 39566
rect 37660 39732 37716 39742
rect 37884 39732 37940 40462
rect 38668 40180 38724 40190
rect 38668 40178 39060 40180
rect 38668 40126 38670 40178
rect 38722 40126 39060 40178
rect 38668 40124 39060 40126
rect 38668 40114 38724 40124
rect 37660 39730 37940 39732
rect 37660 39678 37662 39730
rect 37714 39678 37940 39730
rect 37660 39676 37940 39678
rect 37324 39508 37380 39518
rect 37100 39506 37380 39508
rect 37100 39454 37326 39506
rect 37378 39454 37380 39506
rect 37100 39452 37380 39454
rect 34748 39396 34804 39406
rect 34804 39340 34916 39396
rect 34748 39302 34804 39340
rect 33628 38612 34692 38668
rect 32508 37998 32510 38050
rect 32562 37998 32564 38050
rect 32508 37986 32564 37998
rect 34636 37938 34692 38612
rect 34636 37886 34638 37938
rect 34690 37886 34692 37938
rect 34636 37874 34692 37886
rect 32396 37380 32452 37390
rect 32396 37286 32452 37324
rect 33516 37380 33572 37390
rect 32284 37100 33012 37156
rect 32284 36482 32340 36494
rect 32284 36430 32286 36482
rect 32338 36430 32340 36482
rect 32284 35140 32340 36430
rect 32956 36482 33012 37100
rect 33516 36932 33572 37324
rect 34636 37380 34692 37390
rect 34636 37378 34804 37380
rect 34636 37326 34638 37378
rect 34690 37326 34804 37378
rect 34636 37324 34804 37326
rect 34636 37314 34692 37324
rect 34412 37266 34468 37278
rect 34412 37214 34414 37266
rect 34466 37214 34468 37266
rect 33964 37154 34020 37166
rect 33964 37102 33966 37154
rect 34018 37102 34020 37154
rect 33964 37044 34020 37102
rect 33964 36978 34020 36988
rect 33516 36876 33684 36932
rect 32956 36430 32958 36482
rect 33010 36430 33012 36482
rect 32956 36418 33012 36430
rect 33180 35140 33236 35150
rect 32284 35138 33236 35140
rect 32284 35086 33182 35138
rect 33234 35086 33236 35138
rect 32284 35084 33236 35086
rect 33180 35074 33236 35084
rect 33628 35140 33684 36876
rect 34188 36484 34244 36494
rect 34188 35698 34244 36428
rect 34188 35646 34190 35698
rect 34242 35646 34244 35698
rect 34188 35634 34244 35646
rect 34300 36482 34356 36494
rect 34300 36430 34302 36482
rect 34354 36430 34356 36482
rect 34300 35364 34356 36430
rect 34300 35298 34356 35308
rect 33628 35074 33684 35084
rect 32396 33346 32452 33358
rect 32396 33294 32398 33346
rect 32450 33294 32452 33346
rect 32396 32564 32452 33294
rect 32396 31778 32452 32508
rect 32956 33348 33012 33358
rect 32956 32562 33012 33292
rect 32956 32510 32958 32562
rect 33010 32510 33012 32562
rect 32956 32498 33012 32510
rect 33516 32564 33572 32574
rect 33516 32470 33572 32508
rect 32508 32452 32564 32462
rect 32620 32452 32676 32462
rect 32508 32450 32620 32452
rect 32508 32398 32510 32450
rect 32562 32398 32620 32450
rect 32508 32396 32620 32398
rect 32508 32386 32564 32396
rect 32396 31726 32398 31778
rect 32450 31726 32452 31778
rect 32284 28756 32340 28766
rect 32284 28642 32340 28700
rect 32284 28590 32286 28642
rect 32338 28590 32340 28642
rect 32284 28578 32340 28590
rect 32396 28420 32452 31726
rect 31500 27654 31556 27692
rect 32060 28140 32228 28196
rect 32284 28364 32452 28420
rect 30380 27186 30548 27188
rect 30380 27134 30382 27186
rect 30434 27134 30548 27186
rect 30380 27132 30548 27134
rect 30716 27188 30772 27198
rect 30380 27076 30436 27132
rect 30716 27094 30772 27132
rect 30380 27010 30436 27020
rect 31164 27076 31220 27114
rect 31164 27010 31220 27020
rect 31500 27074 31556 27086
rect 31500 27022 31502 27074
rect 31554 27022 31556 27074
rect 31500 26908 31556 27022
rect 31836 27076 31892 27086
rect 30492 26852 31556 26908
rect 31724 26964 31780 27002
rect 31724 26898 31780 26908
rect 30268 26516 30324 26526
rect 30492 26516 30548 26852
rect 30268 26514 30548 26516
rect 30268 26462 30270 26514
rect 30322 26462 30548 26514
rect 30268 26460 30548 26462
rect 31724 26628 31780 26638
rect 30268 26450 30324 26460
rect 30044 25454 30046 25506
rect 30098 25454 30100 25506
rect 30044 24724 30100 25454
rect 30044 24630 30100 24668
rect 30156 26290 30212 26302
rect 30156 26238 30158 26290
rect 30210 26238 30212 26290
rect 30156 24164 30212 26238
rect 30940 26292 30996 26302
rect 30604 24164 30660 24174
rect 30156 24162 30660 24164
rect 30156 24110 30606 24162
rect 30658 24110 30660 24162
rect 30156 24108 30660 24110
rect 30604 24098 30660 24108
rect 29820 23886 29822 23938
rect 29874 23886 29876 23938
rect 29820 23874 29876 23886
rect 29932 23940 29988 23950
rect 29932 23846 29988 23884
rect 30380 23940 30436 23950
rect 30380 23846 30436 23884
rect 30604 23492 30660 23502
rect 30604 23266 30660 23436
rect 30604 23214 30606 23266
rect 30658 23214 30660 23266
rect 30268 22932 30324 22942
rect 30268 22930 30436 22932
rect 30268 22878 30270 22930
rect 30322 22878 30436 22930
rect 30268 22876 30436 22878
rect 30268 22866 30324 22876
rect 30156 22484 30212 22494
rect 29820 22372 29876 22382
rect 29876 22316 30100 22372
rect 29820 22306 29876 22316
rect 29708 21534 29710 21586
rect 29762 21534 29764 21586
rect 29708 20916 29764 21534
rect 30044 21586 30100 22316
rect 30044 21534 30046 21586
rect 30098 21534 30100 21586
rect 30044 21522 30100 21534
rect 30156 21364 30212 22428
rect 30268 21700 30324 21710
rect 30268 21606 30324 21644
rect 30380 21700 30436 22876
rect 30604 22484 30660 23214
rect 30604 22390 30660 22428
rect 30716 22036 30772 22046
rect 30604 21700 30660 21710
rect 30380 21644 30604 21700
rect 29708 20822 29764 20860
rect 29932 21308 30212 21364
rect 29596 20078 29598 20130
rect 29650 20078 29652 20130
rect 29596 20066 29652 20078
rect 29260 19966 29262 20018
rect 29314 19966 29316 20018
rect 29260 19954 29316 19966
rect 29148 19740 29428 19796
rect 29372 19234 29428 19740
rect 29372 19182 29374 19234
rect 29426 19182 29428 19234
rect 29372 19012 29428 19182
rect 29708 19124 29764 19134
rect 29932 19124 29988 21308
rect 29708 19122 29988 19124
rect 29708 19070 29710 19122
rect 29762 19070 29988 19122
rect 29708 19068 29988 19070
rect 30156 20690 30212 20702
rect 30156 20638 30158 20690
rect 30210 20638 30212 20690
rect 29708 19058 29764 19068
rect 29372 18946 29428 18956
rect 30156 18676 30212 20638
rect 30380 20356 30436 21644
rect 30604 21634 30660 21644
rect 30492 20916 30548 20926
rect 30492 20802 30548 20860
rect 30492 20750 30494 20802
rect 30546 20750 30548 20802
rect 30492 20738 30548 20750
rect 30380 20290 30436 20300
rect 30156 18620 30324 18676
rect 29708 18562 29764 18574
rect 29708 18510 29710 18562
rect 29762 18510 29764 18562
rect 29484 18450 29540 18462
rect 29484 18398 29486 18450
rect 29538 18398 29540 18450
rect 29372 18004 29428 18014
rect 29372 17778 29428 17948
rect 29372 17726 29374 17778
rect 29426 17726 29428 17778
rect 29372 17714 29428 17726
rect 28588 17554 28644 17566
rect 28588 17502 28590 17554
rect 28642 17502 28644 17554
rect 28588 17332 28644 17502
rect 29484 17444 29540 18398
rect 29596 18004 29652 18014
rect 29596 17780 29652 17948
rect 29708 17892 29764 18510
rect 30156 18450 30212 18462
rect 30156 18398 30158 18450
rect 30210 18398 30212 18450
rect 29708 17836 29988 17892
rect 29596 17724 29876 17780
rect 29820 17666 29876 17724
rect 29820 17614 29822 17666
rect 29874 17614 29876 17666
rect 29820 17602 29876 17614
rect 29708 17556 29764 17566
rect 29596 17444 29652 17454
rect 29484 17442 29652 17444
rect 29484 17390 29598 17442
rect 29650 17390 29652 17442
rect 29484 17388 29652 17390
rect 28588 17266 28644 17276
rect 28364 17042 28420 17052
rect 28476 16994 28532 17006
rect 28476 16942 28478 16994
rect 28530 16942 28532 16994
rect 28364 16882 28420 16894
rect 28364 16830 28366 16882
rect 28418 16830 28420 16882
rect 28364 16324 28420 16830
rect 28364 16258 28420 16268
rect 28476 16212 28532 16942
rect 29596 16772 29652 17388
rect 29596 16706 29652 16716
rect 28476 16146 28532 16156
rect 29260 16324 29316 16334
rect 29260 16210 29316 16268
rect 29260 16158 29262 16210
rect 29314 16158 29316 16210
rect 29260 16146 29316 16158
rect 28588 16098 28644 16110
rect 28588 16046 28590 16098
rect 28642 16046 28644 16098
rect 28588 15540 28644 16046
rect 29708 16098 29764 17500
rect 29932 17332 29988 17836
rect 30044 17332 30100 17342
rect 29932 17276 30044 17332
rect 30044 17266 30100 17276
rect 29708 16046 29710 16098
rect 29762 16046 29764 16098
rect 29708 16034 29764 16046
rect 30044 16212 30100 16222
rect 28588 15474 28644 15484
rect 29932 15540 29988 15550
rect 29260 15428 29316 15438
rect 29932 15428 29988 15484
rect 29260 15148 29316 15372
rect 29596 15426 29988 15428
rect 29596 15374 29934 15426
rect 29986 15374 29988 15426
rect 29596 15372 29988 15374
rect 28140 15092 28308 15148
rect 29260 15092 29428 15148
rect 27580 14530 27748 14532
rect 27580 14478 27582 14530
rect 27634 14478 27748 14530
rect 27580 14476 27748 14478
rect 27580 14466 27636 14476
rect 27804 14196 27860 14206
rect 27804 13970 27860 14140
rect 27804 13918 27806 13970
rect 27858 13918 27860 13970
rect 27804 13906 27860 13918
rect 27468 13806 27470 13858
rect 27522 13806 27524 13858
rect 27468 13794 27524 13806
rect 28140 13748 28196 13758
rect 28140 13654 28196 13692
rect 27580 12962 27636 12974
rect 27580 12910 27582 12962
rect 27634 12910 27636 12962
rect 26796 12126 26798 12178
rect 26850 12126 26852 12178
rect 26236 10724 26292 10734
rect 25676 10498 25732 10510
rect 25676 10446 25678 10498
rect 25730 10446 25732 10498
rect 25676 10164 25732 10446
rect 25676 10098 25732 10108
rect 26124 9826 26180 9838
rect 26124 9774 26126 9826
rect 26178 9774 26180 9826
rect 26124 9154 26180 9774
rect 26124 9102 26126 9154
rect 26178 9102 26180 9154
rect 26124 9090 26180 9102
rect 26236 9042 26292 10668
rect 26236 8990 26238 9042
rect 26290 8990 26292 9042
rect 26236 8978 26292 8990
rect 25676 8932 25732 8942
rect 25676 8838 25732 8876
rect 25564 8530 25620 8540
rect 26124 8596 26180 8606
rect 25452 8194 25508 8204
rect 24668 7308 25060 7364
rect 24556 6748 24948 6804
rect 24444 6692 24500 6702
rect 24444 6598 24500 6636
rect 24892 6690 24948 6748
rect 24892 6638 24894 6690
rect 24946 6638 24948 6690
rect 23884 5012 23940 5022
rect 23884 4918 23940 4956
rect 23660 4510 23662 4562
rect 23714 4510 23716 4562
rect 23660 4498 23716 4510
rect 23548 4340 23604 4350
rect 23436 4338 23604 4340
rect 23436 4286 23550 4338
rect 23602 4286 23604 4338
rect 23436 4284 23604 4286
rect 23548 4274 23604 4284
rect 24108 4338 24164 5628
rect 24556 5906 24612 5918
rect 24780 5908 24836 5918
rect 24556 5854 24558 5906
rect 24610 5854 24612 5906
rect 24556 5234 24612 5854
rect 24556 5182 24558 5234
rect 24610 5182 24612 5234
rect 24556 5170 24612 5182
rect 24668 5852 24780 5908
rect 24668 4450 24724 5852
rect 24780 5842 24836 5852
rect 24892 5010 24948 6638
rect 25004 5122 25060 7308
rect 25116 8148 25172 8158
rect 25116 6916 25172 8092
rect 25900 8036 25956 8046
rect 25788 8034 25956 8036
rect 25788 7982 25902 8034
rect 25954 7982 25956 8034
rect 25788 7980 25956 7982
rect 25788 7586 25844 7980
rect 25900 7970 25956 7980
rect 25788 7534 25790 7586
rect 25842 7534 25844 7586
rect 25788 7522 25844 7534
rect 26124 7474 26180 8540
rect 26796 8260 26852 12126
rect 26908 12348 27076 12404
rect 27468 12738 27524 12750
rect 27468 12686 27470 12738
rect 27522 12686 27524 12738
rect 26908 8820 26964 12348
rect 27020 12180 27076 12190
rect 27020 10610 27076 12124
rect 27468 12178 27524 12686
rect 27468 12126 27470 12178
rect 27522 12126 27524 12178
rect 27468 12114 27524 12126
rect 27580 11508 27636 12910
rect 27580 11442 27636 11452
rect 27804 12850 27860 12862
rect 27804 12798 27806 12850
rect 27858 12798 27860 12850
rect 27804 11508 27860 12798
rect 28252 12404 28308 15092
rect 29148 14644 29204 14654
rect 28476 14532 28532 14542
rect 28476 14438 28532 14476
rect 29148 14530 29204 14588
rect 29148 14478 29150 14530
rect 29202 14478 29204 14530
rect 29036 13972 29092 13982
rect 29148 13972 29204 14478
rect 29372 14530 29428 15092
rect 29372 14478 29374 14530
rect 29426 14478 29428 14530
rect 29372 14466 29428 14478
rect 29484 14532 29540 14542
rect 29484 14438 29540 14476
rect 29596 14530 29652 15372
rect 29932 15362 29988 15372
rect 30044 15316 30100 16156
rect 30044 15148 30100 15260
rect 29596 14478 29598 14530
rect 29650 14478 29652 14530
rect 29596 14466 29652 14478
rect 29820 15092 30100 15148
rect 29820 14530 29876 15092
rect 30156 14532 30212 18398
rect 30268 16882 30324 18620
rect 30380 18562 30436 18574
rect 30380 18510 30382 18562
rect 30434 18510 30436 18562
rect 30380 17780 30436 18510
rect 30380 17714 30436 17724
rect 30268 16830 30270 16882
rect 30322 16830 30324 16882
rect 30268 16818 30324 16830
rect 30604 16996 30660 17006
rect 30604 16098 30660 16940
rect 30604 16046 30606 16098
rect 30658 16046 30660 16098
rect 30604 16034 30660 16046
rect 29820 14478 29822 14530
rect 29874 14478 29876 14530
rect 29820 14466 29876 14478
rect 29932 14530 30212 14532
rect 29932 14478 30158 14530
rect 30210 14478 30212 14530
rect 29932 14476 30212 14478
rect 29932 14308 29988 14476
rect 30156 14466 30212 14476
rect 30268 15988 30324 15998
rect 30268 14532 30324 15932
rect 30492 15316 30548 15326
rect 30492 15222 30548 15260
rect 30716 15148 30772 21980
rect 30940 21588 30996 26236
rect 31276 26290 31332 26302
rect 31276 26238 31278 26290
rect 31330 26238 31332 26290
rect 31276 25618 31332 26238
rect 31276 25566 31278 25618
rect 31330 25566 31332 25618
rect 31276 25554 31332 25566
rect 31724 24722 31780 26572
rect 31724 24670 31726 24722
rect 31778 24670 31780 24722
rect 31724 24658 31780 24670
rect 31500 24388 31556 24398
rect 31052 23940 31108 23950
rect 31052 23846 31108 23884
rect 31388 23716 31444 23726
rect 31388 23622 31444 23660
rect 31500 23380 31556 24332
rect 31836 24164 31892 27020
rect 32060 26908 32116 28140
rect 32172 27970 32228 27982
rect 32172 27918 32174 27970
rect 32226 27918 32228 27970
rect 32172 27860 32228 27918
rect 32172 27794 32228 27804
rect 32172 27412 32228 27422
rect 32172 27074 32228 27356
rect 32172 27022 32174 27074
rect 32226 27022 32228 27074
rect 32172 27010 32228 27022
rect 32060 26852 32228 26908
rect 31836 24050 31892 24108
rect 31836 23998 31838 24050
rect 31890 23998 31892 24050
rect 31836 23986 31892 23998
rect 32172 23940 32228 26852
rect 32284 25284 32340 28364
rect 32396 27858 32452 27870
rect 32396 27806 32398 27858
rect 32450 27806 32452 27858
rect 32396 27524 32452 27806
rect 32396 27458 32452 27468
rect 32396 26290 32452 26302
rect 32396 26238 32398 26290
rect 32450 26238 32452 26290
rect 32396 26068 32452 26238
rect 32396 26002 32452 26012
rect 32284 24946 32340 25228
rect 32284 24894 32286 24946
rect 32338 24894 32340 24946
rect 32284 24882 32340 24894
rect 32284 23940 32340 23950
rect 32060 23938 32340 23940
rect 32060 23886 32286 23938
rect 32338 23886 32340 23938
rect 32060 23884 32340 23886
rect 32060 23548 32116 23884
rect 32284 23874 32340 23884
rect 32620 23940 32676 32396
rect 34300 32340 34356 32350
rect 34300 31220 34356 32284
rect 34076 31218 34356 31220
rect 34076 31166 34302 31218
rect 34354 31166 34356 31218
rect 34076 31164 34356 31166
rect 33964 30882 34020 30894
rect 33964 30830 33966 30882
rect 34018 30830 34020 30882
rect 33740 30098 33796 30110
rect 33740 30046 33742 30098
rect 33794 30046 33796 30098
rect 33180 29988 33236 29998
rect 33516 29988 33572 29998
rect 33740 29988 33796 30046
rect 33068 29652 33124 29662
rect 32956 28756 33012 28766
rect 32956 28662 33012 28700
rect 32844 28644 32900 28654
rect 32844 28550 32900 28588
rect 32956 28532 33012 28542
rect 32956 27074 33012 28476
rect 33068 27970 33124 29596
rect 33180 29650 33236 29932
rect 33180 29598 33182 29650
rect 33234 29598 33236 29650
rect 33180 29586 33236 29598
rect 33404 29986 33796 29988
rect 33404 29934 33518 29986
rect 33570 29934 33796 29986
rect 33404 29932 33796 29934
rect 33404 29204 33460 29932
rect 33516 29922 33572 29932
rect 33404 29138 33460 29148
rect 33516 29540 33572 29550
rect 33516 28644 33572 29484
rect 33964 29092 34020 30830
rect 33964 29026 34020 29036
rect 34076 30098 34132 31164
rect 34300 31154 34356 31164
rect 34412 30324 34468 37214
rect 34748 35698 34804 37324
rect 34860 37044 34916 39340
rect 36316 38948 36372 38958
rect 35868 38834 35924 38846
rect 36316 38836 36372 38892
rect 35868 38782 35870 38834
rect 35922 38782 35924 38834
rect 35868 38668 35924 38782
rect 36204 38834 36372 38836
rect 36204 38782 36318 38834
rect 36370 38782 36372 38834
rect 36204 38780 36372 38782
rect 35868 38612 36036 38668
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35420 37266 35476 37278
rect 35420 37214 35422 37266
rect 35474 37214 35476 37266
rect 35420 37156 35476 37214
rect 35868 37266 35924 37278
rect 35868 37214 35870 37266
rect 35922 37214 35924 37266
rect 35420 37090 35476 37100
rect 35756 37154 35812 37166
rect 35756 37102 35758 37154
rect 35810 37102 35812 37154
rect 34860 36978 34916 36988
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35420 36708 35476 36718
rect 35420 36706 35588 36708
rect 35420 36654 35422 36706
rect 35474 36654 35588 36706
rect 35420 36652 35588 36654
rect 35420 36642 35476 36652
rect 35532 35810 35588 36652
rect 35532 35758 35534 35810
rect 35586 35758 35588 35810
rect 35532 35746 35588 35758
rect 34748 35646 34750 35698
rect 34802 35646 34804 35698
rect 34748 34916 34804 35646
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34748 34850 34804 34860
rect 35756 34468 35812 37102
rect 35868 37044 35924 37214
rect 35868 36978 35924 36988
rect 35980 37156 36036 38612
rect 36092 37940 36148 37950
rect 36092 37846 36148 37884
rect 35980 36594 36036 37100
rect 35980 36542 35982 36594
rect 36034 36542 36036 36594
rect 35980 36530 36036 36542
rect 36092 37380 36148 37390
rect 35980 35700 36036 35710
rect 36092 35700 36148 37324
rect 36204 36484 36260 38780
rect 36316 38770 36372 38780
rect 36988 37940 37044 37950
rect 36988 37846 37044 37884
rect 36652 37266 36708 37278
rect 36652 37214 36654 37266
rect 36706 37214 36708 37266
rect 36204 36390 36260 36428
rect 36540 37042 36596 37054
rect 36540 36990 36542 37042
rect 36594 36990 36596 37042
rect 36540 36372 36596 36990
rect 36652 37044 36708 37214
rect 37100 37268 37156 39452
rect 37324 39442 37380 39452
rect 37660 38836 37716 39676
rect 37884 39506 37940 39518
rect 37884 39454 37886 39506
rect 37938 39454 37940 39506
rect 37660 38770 37716 38780
rect 37772 39060 37828 39070
rect 37884 39060 37940 39454
rect 37828 39004 37940 39060
rect 38668 39506 38724 39518
rect 38668 39454 38670 39506
rect 38722 39454 38724 39506
rect 37772 38834 37828 39004
rect 37772 38782 37774 38834
rect 37826 38782 37828 38834
rect 37772 38770 37828 38782
rect 38556 38836 38612 38874
rect 38556 38770 38612 38780
rect 38220 38722 38276 38734
rect 38220 38670 38222 38722
rect 38274 38670 38276 38722
rect 37212 38610 37268 38622
rect 37212 38558 37214 38610
rect 37266 38558 37268 38610
rect 37212 38388 37268 38558
rect 37212 38332 37492 38388
rect 37324 38050 37380 38062
rect 37324 37998 37326 38050
rect 37378 37998 37380 38050
rect 37324 37940 37380 37998
rect 37436 38052 37492 38332
rect 37772 38052 37828 38062
rect 37436 38050 37828 38052
rect 37436 37998 37774 38050
rect 37826 37998 37828 38050
rect 37436 37996 37828 37998
rect 37772 37986 37828 37996
rect 37324 37884 37604 37940
rect 37436 37716 37492 37726
rect 37100 37202 37156 37212
rect 37212 37660 37436 37716
rect 36652 36978 36708 36988
rect 37100 37044 37156 37054
rect 37100 36594 37156 36988
rect 37100 36542 37102 36594
rect 37154 36542 37156 36594
rect 37100 36530 37156 36542
rect 35980 35698 36148 35700
rect 35980 35646 35982 35698
rect 36034 35646 36148 35698
rect 35980 35644 36148 35646
rect 35980 35634 36036 35644
rect 35756 34402 35812 34412
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34748 33124 34804 33134
rect 34636 33122 34804 33124
rect 34636 33070 34750 33122
rect 34802 33070 34804 33122
rect 34636 33068 34804 33070
rect 34636 31780 34692 33068
rect 34748 33058 34804 33068
rect 35532 33124 35588 33134
rect 35532 33122 35924 33124
rect 35532 33070 35534 33122
rect 35586 33070 35924 33122
rect 35532 33068 35924 33070
rect 35532 33058 35588 33068
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35756 31892 35812 31902
rect 34076 30046 34078 30098
rect 34130 30046 34132 30098
rect 33516 28578 33572 28588
rect 33628 28980 33684 28990
rect 33628 28530 33684 28924
rect 33628 28478 33630 28530
rect 33682 28478 33684 28530
rect 33628 28466 33684 28478
rect 33404 28084 33460 28094
rect 33404 27990 33460 28028
rect 33964 28084 34020 28094
rect 33068 27918 33070 27970
rect 33122 27918 33124 27970
rect 33068 27860 33124 27918
rect 33068 27794 33124 27804
rect 33852 27746 33908 27758
rect 33852 27694 33854 27746
rect 33906 27694 33908 27746
rect 33852 27524 33908 27694
rect 33852 27458 33908 27468
rect 32956 27022 32958 27074
rect 33010 27022 33012 27074
rect 32956 27010 33012 27022
rect 33852 27074 33908 27086
rect 33852 27022 33854 27074
rect 33906 27022 33908 27074
rect 33068 26740 33124 26750
rect 33068 26514 33124 26684
rect 33068 26462 33070 26514
rect 33122 26462 33124 26514
rect 33068 26450 33124 26462
rect 33292 26404 33348 26414
rect 33292 26292 33348 26348
rect 33740 26402 33796 26414
rect 33740 26350 33742 26402
rect 33794 26350 33796 26402
rect 33292 26290 33684 26292
rect 33292 26238 33294 26290
rect 33346 26238 33684 26290
rect 33292 26236 33684 26238
rect 33292 26226 33348 26236
rect 32844 26068 32900 26078
rect 32900 26012 33124 26068
rect 32844 26002 32900 26012
rect 33068 24610 33124 26012
rect 33628 24946 33684 26236
rect 33740 25396 33796 26350
rect 33852 25732 33908 27022
rect 33964 26290 34020 28028
rect 34076 27076 34132 30046
rect 34300 30268 34468 30324
rect 34524 31778 34692 31780
rect 34524 31726 34638 31778
rect 34690 31726 34692 31778
rect 34524 31724 34692 31726
rect 34188 29538 34244 29550
rect 34188 29486 34190 29538
rect 34242 29486 34244 29538
rect 34188 27972 34244 29486
rect 34300 28084 34356 30268
rect 34300 28018 34356 28028
rect 34412 30100 34468 30110
rect 34524 30100 34580 31724
rect 34636 31714 34692 31724
rect 35644 31836 35756 31892
rect 34636 31108 34692 31118
rect 34636 31014 34692 31052
rect 34972 30996 35028 31006
rect 34860 30994 35028 30996
rect 34860 30942 34974 30994
rect 35026 30942 35028 30994
rect 34860 30940 35028 30942
rect 34748 30100 34804 30110
rect 34412 30098 34580 30100
rect 34412 30046 34414 30098
rect 34466 30046 34580 30098
rect 34412 30044 34580 30046
rect 34636 30044 34748 30100
rect 34188 27906 34244 27916
rect 34300 27860 34356 27870
rect 34300 27766 34356 27804
rect 34076 27010 34132 27020
rect 33964 26238 33966 26290
rect 34018 26238 34020 26290
rect 33964 26226 34020 26238
rect 34300 26962 34356 26974
rect 34300 26910 34302 26962
rect 34354 26910 34356 26962
rect 34300 26292 34356 26910
rect 33852 25666 33908 25676
rect 33740 25330 33796 25340
rect 34300 25396 34356 26236
rect 34412 26180 34468 30044
rect 34636 29314 34692 30044
rect 34748 30006 34804 30044
rect 34748 29652 34804 29662
rect 34748 29538 34804 29596
rect 34748 29486 34750 29538
rect 34802 29486 34804 29538
rect 34748 29428 34804 29486
rect 34748 29362 34804 29372
rect 34636 29262 34638 29314
rect 34690 29262 34692 29314
rect 34636 29250 34692 29262
rect 34860 29092 34916 30940
rect 34972 30930 35028 30940
rect 35532 30884 35588 30894
rect 35532 30790 35588 30828
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35532 30210 35588 30222
rect 35532 30158 35534 30210
rect 35586 30158 35588 30210
rect 35196 29988 35252 29998
rect 34524 28644 34580 28654
rect 34524 28550 34580 28588
rect 34748 28084 34804 28094
rect 34748 27858 34804 28028
rect 34748 27806 34750 27858
rect 34802 27806 34804 27858
rect 34748 27794 34804 27806
rect 34524 27076 34580 27086
rect 34524 26516 34580 27020
rect 34524 26450 34580 26460
rect 34412 26114 34468 26124
rect 34860 26290 34916 29036
rect 35084 29986 35252 29988
rect 35084 29934 35198 29986
rect 35250 29934 35252 29986
rect 35084 29932 35252 29934
rect 34972 28532 35028 28542
rect 34972 28082 35028 28476
rect 34972 28030 34974 28082
rect 35026 28030 35028 28082
rect 34972 28018 35028 28030
rect 35084 27972 35140 29932
rect 35196 29922 35252 29932
rect 35532 29652 35588 30158
rect 35532 29586 35588 29596
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35308 27972 35364 27982
rect 35084 27970 35364 27972
rect 35084 27918 35310 27970
rect 35362 27918 35364 27970
rect 35084 27916 35364 27918
rect 35308 27906 35364 27916
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35644 27412 35700 31836
rect 35756 31826 35812 31836
rect 35868 31106 35924 33068
rect 35868 31054 35870 31106
rect 35922 31054 35924 31106
rect 35868 31042 35924 31054
rect 36092 30996 36148 35644
rect 36428 36316 36596 36372
rect 36428 35698 36484 36316
rect 36428 35646 36430 35698
rect 36482 35646 36484 35698
rect 36428 35634 36484 35646
rect 36540 35810 36596 35822
rect 36540 35758 36542 35810
rect 36594 35758 36596 35810
rect 36428 32562 36484 32574
rect 36428 32510 36430 32562
rect 36482 32510 36484 32562
rect 36428 32452 36484 32510
rect 36428 32116 36484 32396
rect 36428 32050 36484 32060
rect 36540 31892 36596 35758
rect 37212 35698 37268 37660
rect 37436 37650 37492 37660
rect 37548 37380 37604 37884
rect 37996 37828 38052 37838
rect 37548 37314 37604 37324
rect 37884 37826 38052 37828
rect 37884 37774 37998 37826
rect 38050 37774 38052 37826
rect 37884 37772 38052 37774
rect 37660 37266 37716 37278
rect 37660 37214 37662 37266
rect 37714 37214 37716 37266
rect 37212 35646 37214 35698
rect 37266 35646 37268 35698
rect 37212 35634 37268 35646
rect 37436 37156 37492 37166
rect 37436 34914 37492 37100
rect 37660 36372 37716 37214
rect 37660 36306 37716 36316
rect 37548 36260 37604 36270
rect 37548 36166 37604 36204
rect 37436 34862 37438 34914
rect 37490 34862 37492 34914
rect 37436 34850 37492 34862
rect 37772 35698 37828 35710
rect 37772 35646 37774 35698
rect 37826 35646 37828 35698
rect 37660 34804 37716 34814
rect 37660 34710 37716 34748
rect 37100 34692 37156 34702
rect 37100 34598 37156 34636
rect 37212 34692 37268 34702
rect 37212 34690 37380 34692
rect 37212 34638 37214 34690
rect 37266 34638 37380 34690
rect 37212 34636 37380 34638
rect 37212 34626 37268 34636
rect 37212 34468 37268 34478
rect 36988 34020 37044 34030
rect 36988 33926 37044 33964
rect 37212 33684 37268 34412
rect 37212 33618 37268 33628
rect 37100 33234 37156 33246
rect 37100 33182 37102 33234
rect 37154 33182 37156 33234
rect 36540 31826 36596 31836
rect 36764 32564 36820 32574
rect 36204 31668 36260 31678
rect 36204 31666 36708 31668
rect 36204 31614 36206 31666
rect 36258 31614 36708 31666
rect 36204 31612 36708 31614
rect 36204 31602 36260 31612
rect 36540 31332 36596 31342
rect 36204 30996 36260 31006
rect 36092 30994 36260 30996
rect 36092 30942 36206 30994
rect 36258 30942 36260 30994
rect 36092 30940 36260 30942
rect 36092 30884 36148 30940
rect 36204 30930 36260 30940
rect 36092 30818 36148 30828
rect 35756 30100 35812 30110
rect 35756 30006 35812 30044
rect 36316 30098 36372 30110
rect 36316 30046 36318 30098
rect 36370 30046 36372 30098
rect 36316 29540 36372 30046
rect 36540 29876 36596 31276
rect 36652 30994 36708 31612
rect 36652 30942 36654 30994
rect 36706 30942 36708 30994
rect 36652 30930 36708 30942
rect 36764 30660 36820 32508
rect 36988 32564 37044 32574
rect 37100 32564 37156 33182
rect 36988 32562 37156 32564
rect 36988 32510 36990 32562
rect 37042 32510 37156 32562
rect 36988 32508 37156 32510
rect 36988 32452 37044 32508
rect 36988 32386 37044 32396
rect 37324 31332 37380 34636
rect 37772 34690 37828 35646
rect 37772 34638 37774 34690
rect 37826 34638 37828 34690
rect 37772 34626 37828 34638
rect 37884 34468 37940 37772
rect 37996 37762 38052 37772
rect 38108 37156 38164 37166
rect 38108 37062 38164 37100
rect 37996 37044 38052 37054
rect 37996 35026 38052 36988
rect 38220 36484 38276 38670
rect 38556 38612 38612 38622
rect 38220 36418 38276 36428
rect 38444 37938 38500 37950
rect 38444 37886 38446 37938
rect 38498 37886 38500 37938
rect 38444 37716 38500 37886
rect 37996 34974 37998 35026
rect 38050 34974 38052 35026
rect 37996 34962 38052 34974
rect 38108 36372 38164 36382
rect 38108 35028 38164 36316
rect 38220 35028 38276 35038
rect 38108 35026 38276 35028
rect 38108 34974 38222 35026
rect 38274 34974 38276 35026
rect 38108 34972 38276 34974
rect 37548 34412 37940 34468
rect 37436 34132 37492 34142
rect 37436 34038 37492 34076
rect 37548 32340 37604 34412
rect 37660 34244 37716 34254
rect 37660 34242 37940 34244
rect 37660 34190 37662 34242
rect 37714 34190 37940 34242
rect 37660 34188 37940 34190
rect 37660 34178 37716 34188
rect 37660 33124 37716 33134
rect 37660 33030 37716 33068
rect 37772 32562 37828 32574
rect 37772 32510 37774 32562
rect 37826 32510 37828 32562
rect 37548 32284 37716 32340
rect 37548 31892 37604 31902
rect 37548 31798 37604 31836
rect 37324 31266 37380 31276
rect 36876 31106 36932 31118
rect 36876 31054 36878 31106
rect 36930 31054 36932 31106
rect 36876 30884 36932 31054
rect 37548 31108 37604 31118
rect 37548 30994 37604 31052
rect 37548 30942 37550 30994
rect 37602 30942 37604 30994
rect 37548 30930 37604 30942
rect 36876 30818 36932 30828
rect 37324 30884 37380 30894
rect 37380 30828 37492 30884
rect 37324 30818 37380 30828
rect 36764 30604 36932 30660
rect 36092 29202 36148 29214
rect 36092 29150 36094 29202
rect 36146 29150 36148 29202
rect 35868 28868 35924 28878
rect 35868 28642 35924 28812
rect 35868 28590 35870 28642
rect 35922 28590 35924 28642
rect 35868 28578 35924 28590
rect 35196 27402 35460 27412
rect 35532 27356 35700 27412
rect 35756 27858 35812 27870
rect 35756 27806 35758 27858
rect 35810 27806 35812 27858
rect 35420 27300 35476 27310
rect 35532 27300 35588 27356
rect 35420 27298 35588 27300
rect 35420 27246 35422 27298
rect 35474 27246 35588 27298
rect 35420 27244 35588 27246
rect 35420 27234 35476 27244
rect 35196 27188 35252 27198
rect 35084 26852 35140 26862
rect 35084 26758 35140 26796
rect 34860 26238 34862 26290
rect 34914 26238 34916 26290
rect 34860 25618 34916 26238
rect 35196 26180 35252 27132
rect 35756 26628 35812 27806
rect 36092 27858 36148 29150
rect 36316 28532 36372 29484
rect 36428 29820 36596 29876
rect 36764 30436 36820 30446
rect 36428 29092 36484 29820
rect 36764 29426 36820 30380
rect 36764 29374 36766 29426
rect 36818 29374 36820 29426
rect 36764 29362 36820 29374
rect 36428 28754 36484 29036
rect 36428 28702 36430 28754
rect 36482 28702 36484 28754
rect 36428 28690 36484 28702
rect 36540 28868 36596 28878
rect 36316 28466 36372 28476
rect 36092 27806 36094 27858
rect 36146 27806 36148 27858
rect 36092 27794 36148 27806
rect 36316 27970 36372 27982
rect 36316 27918 36318 27970
rect 36370 27918 36372 27970
rect 36092 27076 36148 27086
rect 36092 26982 36148 27020
rect 36204 26964 36260 26974
rect 36316 26964 36372 27918
rect 36204 26962 36372 26964
rect 36204 26910 36206 26962
rect 36258 26910 36372 26962
rect 36204 26908 36372 26910
rect 36204 26898 36260 26908
rect 35756 26514 35812 26572
rect 35756 26462 35758 26514
rect 35810 26462 35812 26514
rect 35756 26450 35812 26462
rect 36428 26516 36484 26526
rect 36540 26516 36596 28812
rect 36428 26514 36596 26516
rect 36428 26462 36430 26514
rect 36482 26462 36596 26514
rect 36428 26460 36596 26462
rect 36764 27858 36820 27870
rect 36764 27806 36766 27858
rect 36818 27806 36820 27858
rect 36428 26450 36484 26460
rect 34860 25566 34862 25618
rect 34914 25566 34916 25618
rect 34860 25554 34916 25566
rect 35084 26178 35252 26180
rect 35084 26126 35198 26178
rect 35250 26126 35252 26178
rect 35084 26124 35252 26126
rect 35084 25396 35140 26124
rect 35196 26114 35252 26124
rect 36764 26178 36820 27806
rect 36764 26126 36766 26178
rect 36818 26126 36820 26178
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34300 25330 34356 25340
rect 34524 25340 35140 25396
rect 35196 25732 35252 25742
rect 33628 24894 33630 24946
rect 33682 24894 33684 24946
rect 33628 24882 33684 24894
rect 34524 24722 34580 25340
rect 35196 24946 35252 25676
rect 36428 25508 36484 25518
rect 36428 25414 36484 25452
rect 36764 25508 36820 26126
rect 36764 25442 36820 25452
rect 35196 24894 35198 24946
rect 35250 24894 35252 24946
rect 35196 24882 35252 24894
rect 35644 25396 35700 25406
rect 35644 24834 35700 25340
rect 35644 24782 35646 24834
rect 35698 24782 35700 24834
rect 35644 24770 35700 24782
rect 34972 24724 35028 24734
rect 34524 24670 34526 24722
rect 34578 24670 34580 24722
rect 34524 24658 34580 24670
rect 34636 24722 35028 24724
rect 34636 24670 34974 24722
rect 35026 24670 35028 24722
rect 34636 24668 35028 24670
rect 34188 24612 34244 24622
rect 33068 24558 33070 24610
rect 33122 24558 33124 24610
rect 33068 24546 33124 24558
rect 34076 24610 34244 24612
rect 34076 24558 34190 24610
rect 34242 24558 34244 24610
rect 34076 24556 34244 24558
rect 32620 23826 32676 23884
rect 33628 23940 33684 23950
rect 33628 23938 33796 23940
rect 33628 23886 33630 23938
rect 33682 23886 33796 23938
rect 33628 23884 33796 23886
rect 33628 23874 33684 23884
rect 32620 23774 32622 23826
rect 32674 23774 32676 23826
rect 32620 23762 32676 23774
rect 32732 23828 32788 23838
rect 32788 23772 32900 23828
rect 32732 23762 32788 23772
rect 31052 23266 31108 23278
rect 31052 23214 31054 23266
rect 31106 23214 31108 23266
rect 31052 22260 31108 23214
rect 31500 23266 31556 23324
rect 31836 23492 32116 23548
rect 31836 23378 31892 23492
rect 31836 23326 31838 23378
rect 31890 23326 31892 23378
rect 31836 23314 31892 23326
rect 32284 23380 32340 23390
rect 32284 23286 32340 23324
rect 31500 23214 31502 23266
rect 31554 23214 31556 23266
rect 31500 23202 31556 23214
rect 32620 23156 32676 23166
rect 32396 22594 32452 22606
rect 32396 22542 32398 22594
rect 32450 22542 32452 22594
rect 32284 22370 32340 22382
rect 32284 22318 32286 22370
rect 32338 22318 32340 22370
rect 31164 22260 31220 22270
rect 31052 22258 31220 22260
rect 31052 22206 31166 22258
rect 31218 22206 31220 22258
rect 31052 22204 31220 22206
rect 31164 21924 31220 22204
rect 32284 22260 32340 22318
rect 32284 22194 32340 22204
rect 31164 21858 31220 21868
rect 31276 22146 31332 22158
rect 31276 22094 31278 22146
rect 31330 22094 31332 22146
rect 31276 21700 31332 22094
rect 31276 21634 31332 21644
rect 32284 22036 32340 22046
rect 31500 21588 31556 21598
rect 30940 21586 31108 21588
rect 30940 21534 30942 21586
rect 30994 21534 31108 21586
rect 30940 21532 31108 21534
rect 30940 21522 30996 21532
rect 30940 20804 30996 20814
rect 30828 20802 30996 20804
rect 30828 20750 30942 20802
rect 30994 20750 30996 20802
rect 30828 20748 30996 20750
rect 30828 20242 30884 20748
rect 30940 20738 30996 20748
rect 31052 20468 31108 21532
rect 31500 21494 31556 21532
rect 31164 21364 31220 21374
rect 31164 20690 31220 21308
rect 32060 21028 32116 21038
rect 31164 20638 31166 20690
rect 31218 20638 31220 20690
rect 31164 20626 31220 20638
rect 31612 20690 31668 20702
rect 31612 20638 31614 20690
rect 31666 20638 31668 20690
rect 31612 20468 31668 20638
rect 31052 20412 31668 20468
rect 30828 20190 30830 20242
rect 30882 20190 30884 20242
rect 30828 20178 30884 20190
rect 31724 20020 31780 20030
rect 31724 19926 31780 19964
rect 32060 19906 32116 20972
rect 32060 19854 32062 19906
rect 32114 19854 32116 19906
rect 32060 19842 32116 19854
rect 32172 19684 32228 19694
rect 32172 19010 32228 19628
rect 32172 18958 32174 19010
rect 32226 18958 32228 19010
rect 32172 18900 32228 18958
rect 31836 18844 32228 18900
rect 31724 18340 31780 18350
rect 31724 18246 31780 18284
rect 31388 17780 31444 17790
rect 31276 17668 31332 17678
rect 31052 17666 31332 17668
rect 31052 17614 31278 17666
rect 31330 17614 31332 17666
rect 31052 17612 31332 17614
rect 30940 17442 30996 17454
rect 30940 17390 30942 17442
rect 30994 17390 30996 17442
rect 30828 16996 30884 17006
rect 30828 15988 30884 16940
rect 30940 16772 30996 17390
rect 30940 16706 30996 16716
rect 30940 15988 30996 15998
rect 30828 15986 30996 15988
rect 30828 15934 30942 15986
rect 30994 15934 30996 15986
rect 30828 15932 30996 15934
rect 30940 15922 30996 15932
rect 31052 15540 31108 17612
rect 31276 17602 31332 17612
rect 31276 16100 31332 16110
rect 31388 16100 31444 17724
rect 31724 17668 31780 17678
rect 31724 17574 31780 17612
rect 31500 16660 31556 16670
rect 31500 16658 31780 16660
rect 31500 16606 31502 16658
rect 31554 16606 31780 16658
rect 31500 16604 31780 16606
rect 31500 16594 31556 16604
rect 31724 16210 31780 16604
rect 31724 16158 31726 16210
rect 31778 16158 31780 16210
rect 31724 16146 31780 16158
rect 31276 16098 31444 16100
rect 31276 16046 31278 16098
rect 31330 16046 31444 16098
rect 31276 16044 31444 16046
rect 31276 16034 31332 16044
rect 31052 15446 31108 15484
rect 31836 15148 31892 18844
rect 32284 18788 32340 21980
rect 32396 21586 32452 22542
rect 32620 22370 32676 23100
rect 32620 22318 32622 22370
rect 32674 22318 32676 22370
rect 32620 22306 32676 22318
rect 32396 21534 32398 21586
rect 32450 21534 32452 21586
rect 32396 21522 32452 21534
rect 32396 20802 32452 20814
rect 32396 20750 32398 20802
rect 32450 20750 32452 20802
rect 32396 19124 32452 20750
rect 32508 20018 32564 20030
rect 32508 19966 32510 20018
rect 32562 19966 32564 20018
rect 32508 19796 32564 19966
rect 32508 19730 32564 19740
rect 32396 19058 32452 19068
rect 32732 19234 32788 19246
rect 32732 19182 32734 19234
rect 32786 19182 32788 19234
rect 32060 18732 32340 18788
rect 31948 18564 32004 18574
rect 31948 18470 32004 18508
rect 30716 15092 30884 15148
rect 30268 14466 30324 14476
rect 30828 14530 30884 15092
rect 30828 14478 30830 14530
rect 30882 14478 30884 14530
rect 30828 14466 30884 14478
rect 31612 15092 31892 15148
rect 29596 14252 29988 14308
rect 30492 14306 30548 14318
rect 30492 14254 30494 14306
rect 30546 14254 30548 14306
rect 29036 13970 29204 13972
rect 29036 13918 29038 13970
rect 29090 13918 29204 13970
rect 29036 13916 29204 13918
rect 29484 14196 29540 14206
rect 29036 13906 29092 13916
rect 28252 12338 28308 12348
rect 28476 13858 28532 13870
rect 28476 13806 28478 13858
rect 28530 13806 28532 13858
rect 28476 12292 28532 13806
rect 29260 13746 29316 13758
rect 29260 13694 29262 13746
rect 29314 13694 29316 13746
rect 29260 13300 29316 13694
rect 29260 13234 29316 13244
rect 28476 12226 28532 12236
rect 27804 11394 27860 11452
rect 27804 11342 27806 11394
rect 27858 11342 27860 11394
rect 27356 11284 27412 11294
rect 27020 10558 27022 10610
rect 27074 10558 27076 10610
rect 27020 10546 27076 10558
rect 27132 11282 27412 11284
rect 27132 11230 27358 11282
rect 27410 11230 27412 11282
rect 27132 11228 27412 11230
rect 27132 9826 27188 11228
rect 27356 11218 27412 11228
rect 27804 10724 27860 11342
rect 27804 10658 27860 10668
rect 28252 12178 28308 12190
rect 28252 12126 28254 12178
rect 28306 12126 28308 12178
rect 28252 10722 28308 12126
rect 29260 12066 29316 12078
rect 29260 12014 29262 12066
rect 29314 12014 29316 12066
rect 29148 11172 29204 11182
rect 29148 11078 29204 11116
rect 28252 10670 28254 10722
rect 28306 10670 28308 10722
rect 28252 10658 28308 10670
rect 29260 10500 29316 12014
rect 29260 10434 29316 10444
rect 27132 9774 27134 9826
rect 27186 9774 27188 9826
rect 27132 9762 27188 9774
rect 29484 9492 29540 14140
rect 29596 13970 29652 14252
rect 29596 13918 29598 13970
rect 29650 13918 29652 13970
rect 29596 13906 29652 13918
rect 29708 13972 29764 13982
rect 29596 12178 29652 12190
rect 29596 12126 29598 12178
rect 29650 12126 29652 12178
rect 29596 11956 29652 12126
rect 29596 11890 29652 11900
rect 29596 11508 29652 11518
rect 29596 11414 29652 11452
rect 29596 10500 29652 10510
rect 29596 10406 29652 10444
rect 29596 9828 29652 9838
rect 29708 9828 29764 13916
rect 30492 13972 30548 14254
rect 31164 14308 31220 14318
rect 31164 14214 31220 14252
rect 30492 13906 30548 13916
rect 30492 13746 30548 13758
rect 30492 13694 30494 13746
rect 30546 13694 30548 13746
rect 29932 13634 29988 13646
rect 29932 13582 29934 13634
rect 29986 13582 29988 13634
rect 29820 13412 29876 13422
rect 29820 12962 29876 13356
rect 29820 12910 29822 12962
rect 29874 12910 29876 12962
rect 29820 12898 29876 12910
rect 29932 12852 29988 13582
rect 29932 10610 29988 12796
rect 30044 13186 30100 13198
rect 30044 13134 30046 13186
rect 30098 13134 30100 13186
rect 30044 12178 30100 13134
rect 30268 12962 30324 12974
rect 30268 12910 30270 12962
rect 30322 12910 30324 12962
rect 30268 12628 30324 12910
rect 30380 12962 30436 12974
rect 30380 12910 30382 12962
rect 30434 12910 30436 12962
rect 30380 12852 30436 12910
rect 30380 12786 30436 12796
rect 30268 12562 30324 12572
rect 30268 12404 30324 12414
rect 30268 12310 30324 12348
rect 30044 12126 30046 12178
rect 30098 12126 30100 12178
rect 30044 12114 30100 12126
rect 30156 12068 30212 12078
rect 30156 11396 30212 12012
rect 29932 10558 29934 10610
rect 29986 10558 29988 10610
rect 29932 10546 29988 10558
rect 30044 11394 30212 11396
rect 30044 11342 30158 11394
rect 30210 11342 30212 11394
rect 30044 11340 30212 11342
rect 30044 10164 30100 11340
rect 30156 11330 30212 11340
rect 30268 11844 30324 11854
rect 29596 9826 29764 9828
rect 29596 9774 29598 9826
rect 29650 9774 29764 9826
rect 29596 9772 29764 9774
rect 29820 10108 30100 10164
rect 29596 9762 29652 9772
rect 29820 9714 29876 10108
rect 29820 9662 29822 9714
rect 29874 9662 29876 9714
rect 29820 9650 29876 9662
rect 29484 9436 29876 9492
rect 26908 8754 26964 8764
rect 29596 9154 29652 9166
rect 29596 9102 29598 9154
rect 29650 9102 29652 9154
rect 29596 8484 29652 9102
rect 29820 9042 29876 9436
rect 29820 8990 29822 9042
rect 29874 8990 29876 9042
rect 29820 8978 29876 8990
rect 26796 8194 26852 8204
rect 26908 8258 26964 8270
rect 26908 8206 26910 8258
rect 26962 8206 26964 8258
rect 26124 7422 26126 7474
rect 26178 7422 26180 7474
rect 26124 7410 26180 7422
rect 26684 8146 26740 8158
rect 26684 8094 26686 8146
rect 26738 8094 26740 8146
rect 26684 7474 26740 8094
rect 26908 8036 26964 8206
rect 27244 8260 27300 8270
rect 27020 8148 27076 8158
rect 27020 8054 27076 8092
rect 26908 7970 26964 7980
rect 26796 7700 26852 7710
rect 26796 7606 26852 7644
rect 27244 7586 27300 8204
rect 29484 8260 29540 8270
rect 27580 8148 27636 8158
rect 27580 8054 27636 8092
rect 27244 7534 27246 7586
rect 27298 7534 27300 7586
rect 27244 7522 27300 7534
rect 26684 7422 26686 7474
rect 26738 7422 26740 7474
rect 26684 7410 26740 7422
rect 28028 7474 28084 7486
rect 28028 7422 28030 7474
rect 28082 7422 28084 7474
rect 25116 6860 25508 6916
rect 25340 6692 25396 6702
rect 25340 6130 25396 6636
rect 25452 6692 25508 6860
rect 28028 6914 28084 7422
rect 28028 6862 28030 6914
rect 28082 6862 28084 6914
rect 28028 6850 28084 6862
rect 28364 7476 28420 7486
rect 27580 6804 27636 6814
rect 25452 6690 25732 6692
rect 25452 6638 25454 6690
rect 25506 6638 25732 6690
rect 25452 6636 25732 6638
rect 25452 6626 25508 6636
rect 25340 6078 25342 6130
rect 25394 6078 25396 6130
rect 25340 6066 25396 6078
rect 25228 5906 25284 5918
rect 25228 5854 25230 5906
rect 25282 5854 25284 5906
rect 25228 5796 25284 5854
rect 25676 5908 25732 6636
rect 25676 5814 25732 5852
rect 27580 5906 27636 6748
rect 28364 6804 28420 7420
rect 28364 6690 28420 6748
rect 28812 7474 28868 7486
rect 28812 7422 28814 7474
rect 28866 7422 28868 7474
rect 28364 6638 28366 6690
rect 28418 6638 28420 6690
rect 28364 6626 28420 6638
rect 28588 6692 28644 6702
rect 27580 5854 27582 5906
rect 27634 5854 27636 5906
rect 25228 5730 25284 5740
rect 25452 5684 25508 5694
rect 25452 5590 25508 5628
rect 27580 5346 27636 5854
rect 27580 5294 27582 5346
rect 27634 5294 27636 5346
rect 27580 5282 27636 5294
rect 25004 5070 25006 5122
rect 25058 5070 25060 5122
rect 25004 5058 25060 5070
rect 28588 5122 28644 6636
rect 28812 5794 28868 7422
rect 29484 7476 29540 8204
rect 29484 7382 29540 7420
rect 29148 6692 29204 6702
rect 29148 6578 29204 6636
rect 29484 6692 29540 6702
rect 29596 6692 29652 8428
rect 30044 8148 30100 10108
rect 30268 9938 30324 11788
rect 30492 11396 30548 13694
rect 31612 13746 31668 15092
rect 31724 14868 31780 14878
rect 31724 14644 31780 14812
rect 32060 14756 32116 18732
rect 32732 18452 32788 19182
rect 32732 18386 32788 18396
rect 32508 18338 32564 18350
rect 32508 18286 32510 18338
rect 32562 18286 32564 18338
rect 32508 18116 32564 18286
rect 32508 18050 32564 18060
rect 32284 16884 32340 16894
rect 32284 16770 32340 16828
rect 32284 16718 32286 16770
rect 32338 16718 32340 16770
rect 32172 16100 32228 16110
rect 32172 16006 32228 16044
rect 32284 15652 32340 16718
rect 32844 16660 32900 23772
rect 33180 23826 33236 23838
rect 33180 23774 33182 23826
rect 33234 23774 33236 23826
rect 33180 23492 33236 23774
rect 33236 23436 33348 23492
rect 33180 23426 33236 23436
rect 33180 23156 33236 23166
rect 33180 23042 33236 23100
rect 33180 22990 33182 23042
rect 33234 22990 33236 23042
rect 33180 22978 33236 22990
rect 33292 22148 33348 23436
rect 33516 23154 33572 23166
rect 33516 23102 33518 23154
rect 33570 23102 33572 23154
rect 33516 22932 33572 23102
rect 33516 22866 33572 22876
rect 33628 23044 33684 23054
rect 33628 22596 33684 22988
rect 33740 22820 33796 23884
rect 33964 23938 34020 23950
rect 33964 23886 33966 23938
rect 34018 23886 34020 23938
rect 33852 23156 33908 23166
rect 33964 23156 34020 23886
rect 34076 23380 34132 24556
rect 34188 24546 34244 24556
rect 34636 24164 34692 24668
rect 34972 24658 35028 24668
rect 36316 24722 36372 24734
rect 36316 24670 36318 24722
rect 36370 24670 36372 24722
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 34188 24108 34692 24164
rect 34188 23826 34244 24108
rect 34860 23940 34916 23950
rect 34860 23938 35028 23940
rect 34860 23886 34862 23938
rect 34914 23886 35028 23938
rect 34860 23884 35028 23886
rect 34860 23874 34916 23884
rect 34188 23774 34190 23826
rect 34242 23774 34244 23826
rect 34188 23762 34244 23774
rect 34076 23324 34692 23380
rect 34076 23156 34132 23166
rect 33964 23100 34076 23156
rect 33852 23062 33908 23100
rect 34076 23090 34132 23100
rect 33740 22764 34132 22820
rect 33404 22540 33908 22596
rect 33404 22370 33460 22540
rect 33404 22318 33406 22370
rect 33458 22318 33460 22370
rect 33404 22306 33460 22318
rect 33516 22372 33572 22382
rect 33516 22278 33572 22316
rect 33292 22092 33684 22148
rect 33292 21924 33348 21934
rect 32956 21588 33012 21598
rect 32956 21494 33012 21532
rect 33292 21586 33348 21868
rect 33292 21534 33294 21586
rect 33346 21534 33348 21586
rect 33292 21522 33348 21534
rect 33292 20804 33348 20814
rect 33628 20804 33684 22092
rect 33740 21700 33796 21710
rect 33740 21586 33796 21644
rect 33740 21534 33742 21586
rect 33794 21534 33796 21586
rect 33740 21522 33796 21534
rect 33740 21028 33796 21038
rect 33852 21028 33908 22540
rect 33796 20972 33908 21028
rect 33964 21588 34020 21598
rect 33740 20934 33796 20972
rect 33852 20804 33908 20814
rect 33628 20802 33908 20804
rect 33628 20750 33854 20802
rect 33906 20750 33908 20802
rect 33628 20748 33908 20750
rect 33292 20710 33348 20748
rect 33852 20738 33908 20748
rect 33516 20244 33572 20254
rect 33516 20132 33572 20188
rect 33404 20130 33572 20132
rect 33404 20078 33518 20130
rect 33570 20078 33572 20130
rect 33404 20076 33572 20078
rect 33180 20020 33236 20030
rect 33180 19926 33236 19964
rect 33404 19124 33460 20076
rect 33516 20066 33572 20076
rect 33964 19796 34020 21532
rect 33740 19794 34020 19796
rect 33740 19742 33966 19794
rect 34018 19742 34020 19794
rect 33740 19740 34020 19742
rect 33516 19348 33572 19358
rect 33516 19254 33572 19292
rect 33404 19068 33572 19124
rect 32844 16594 32900 16604
rect 33068 19010 33124 19022
rect 33068 18958 33070 19010
rect 33122 18958 33124 19010
rect 33068 18564 33124 18958
rect 33068 16660 33124 18508
rect 33180 18340 33236 18350
rect 33180 17220 33236 18284
rect 33180 17164 33460 17220
rect 33180 16882 33236 17164
rect 33180 16830 33182 16882
rect 33234 16830 33236 16882
rect 33180 16818 33236 16830
rect 33292 16994 33348 17006
rect 33292 16942 33294 16994
rect 33346 16942 33348 16994
rect 33068 16594 33124 16604
rect 33292 16548 33348 16942
rect 33180 16492 33348 16548
rect 33180 16436 33236 16492
rect 32732 16380 33236 16436
rect 32508 16100 32564 16110
rect 32284 15586 32340 15596
rect 32396 16098 32564 16100
rect 32396 16046 32510 16098
rect 32562 16046 32564 16098
rect 32396 16044 32564 16046
rect 32396 15538 32452 16044
rect 32508 16034 32564 16044
rect 32732 15986 32788 16380
rect 33404 16324 33460 17164
rect 33292 16268 33460 16324
rect 32732 15934 32734 15986
rect 32786 15934 32788 15986
rect 32732 15922 32788 15934
rect 33180 15986 33236 15998
rect 33180 15934 33182 15986
rect 33234 15934 33236 15986
rect 33180 15652 33236 15934
rect 33180 15586 33236 15596
rect 32396 15486 32398 15538
rect 32450 15486 32452 15538
rect 32396 15474 32452 15486
rect 33068 15428 33124 15438
rect 32060 14690 32116 14700
rect 32844 15426 33124 15428
rect 32844 15374 33070 15426
rect 33122 15374 33124 15426
rect 32844 15372 33124 15374
rect 32620 14644 32676 14654
rect 31724 14642 32004 14644
rect 31724 14590 31726 14642
rect 31778 14590 32004 14642
rect 31724 14588 32004 14590
rect 31724 14578 31780 14588
rect 31948 14532 32004 14588
rect 32620 14550 32676 14588
rect 32060 14532 32116 14542
rect 31948 14530 32116 14532
rect 31948 14478 32062 14530
rect 32114 14478 32116 14530
rect 31948 14476 32116 14478
rect 32060 14466 32116 14476
rect 32396 14420 32452 14430
rect 32284 14308 32340 14318
rect 32060 13860 32116 13870
rect 31612 13694 31614 13746
rect 31666 13694 31668 13746
rect 31276 13634 31332 13646
rect 31276 13582 31278 13634
rect 31330 13582 31332 13634
rect 31164 13412 31220 13422
rect 31052 12964 31108 12974
rect 31052 12870 31108 12908
rect 30492 11330 30548 11340
rect 30604 12628 30660 12638
rect 30604 11506 30660 12572
rect 30940 12292 30996 12302
rect 30940 12178 30996 12236
rect 30940 12126 30942 12178
rect 30994 12126 30996 12178
rect 30940 12114 30996 12126
rect 31164 11844 31220 13356
rect 31276 13188 31332 13582
rect 31388 13188 31444 13198
rect 31276 13132 31388 13188
rect 31388 12962 31444 13132
rect 31388 12910 31390 12962
rect 31442 12910 31444 12962
rect 31388 12898 31444 12910
rect 31500 12740 31556 12750
rect 31500 12178 31556 12684
rect 31500 12126 31502 12178
rect 31554 12126 31556 12178
rect 31500 12114 31556 12126
rect 31220 11788 31556 11844
rect 31164 11750 31220 11788
rect 30604 11454 30606 11506
rect 30658 11454 30660 11506
rect 30604 11172 30660 11454
rect 30380 11116 30660 11172
rect 30380 10610 30436 11116
rect 30380 10558 30382 10610
rect 30434 10558 30436 10610
rect 30380 10546 30436 10558
rect 31500 10610 31556 11788
rect 31500 10558 31502 10610
rect 31554 10558 31556 10610
rect 31500 10546 31556 10558
rect 30268 9886 30270 9938
rect 30322 9886 30324 9938
rect 30268 9874 30324 9886
rect 31164 9940 31220 9950
rect 31164 9826 31220 9884
rect 31164 9774 31166 9826
rect 31218 9774 31220 9826
rect 31164 9762 31220 9774
rect 31388 9828 31444 9838
rect 31388 9714 31444 9772
rect 31388 9662 31390 9714
rect 31442 9662 31444 9714
rect 31388 9650 31444 9662
rect 30716 9602 30772 9614
rect 30716 9550 30718 9602
rect 30770 9550 30772 9602
rect 30716 8484 30772 9550
rect 30940 9268 30996 9278
rect 30940 9174 30996 9212
rect 31276 8932 31332 8942
rect 31612 8932 31668 13694
rect 31948 13858 32116 13860
rect 31948 13806 32062 13858
rect 32114 13806 32116 13858
rect 31948 13804 32116 13806
rect 31836 12964 31892 12974
rect 31836 12850 31892 12908
rect 31836 12798 31838 12850
rect 31890 12798 31892 12850
rect 31836 11844 31892 12798
rect 31836 11778 31892 11788
rect 31724 11396 31780 11406
rect 31724 9714 31780 11340
rect 31724 9662 31726 9714
rect 31778 9662 31780 9714
rect 31724 9650 31780 9662
rect 31948 9940 32004 13804
rect 32060 13794 32116 13804
rect 32284 13746 32340 14252
rect 32284 13694 32286 13746
rect 32338 13694 32340 13746
rect 32284 13682 32340 13694
rect 32284 13188 32340 13198
rect 32284 13094 32340 13132
rect 32060 12852 32116 12862
rect 32060 12180 32116 12796
rect 32172 12740 32228 12750
rect 32172 12646 32228 12684
rect 32396 12516 32452 14364
rect 32844 13748 32900 15372
rect 33068 15362 33124 15372
rect 33292 14644 33348 16268
rect 33404 15428 33460 15438
rect 33516 15428 33572 19068
rect 33404 15426 33572 15428
rect 33404 15374 33406 15426
rect 33458 15374 33572 15426
rect 33404 15372 33572 15374
rect 33628 18116 33684 18126
rect 33404 15362 33460 15372
rect 33628 15148 33684 18060
rect 33740 17668 33796 19740
rect 33964 19730 34020 19740
rect 34076 20690 34132 22764
rect 34300 22372 34356 22382
rect 34300 22370 34468 22372
rect 34300 22318 34302 22370
rect 34354 22318 34468 22370
rect 34300 22316 34468 22318
rect 34300 22306 34356 22316
rect 34076 20638 34078 20690
rect 34130 20638 34132 20690
rect 34076 19684 34132 20638
rect 34412 20802 34468 22316
rect 34524 22258 34580 22270
rect 34524 22206 34526 22258
rect 34578 22206 34580 22258
rect 34524 21700 34580 22206
rect 34636 21812 34692 23324
rect 34972 23154 35028 23884
rect 35420 23938 35476 23950
rect 35420 23886 35422 23938
rect 35474 23886 35476 23938
rect 35420 23828 35476 23886
rect 35420 23762 35476 23772
rect 36204 23938 36260 23950
rect 36204 23886 36206 23938
rect 36258 23886 36260 23938
rect 36204 23716 36260 23886
rect 36204 23650 36260 23660
rect 34972 23102 34974 23154
rect 35026 23102 35028 23154
rect 34972 22260 35028 23102
rect 35756 23154 35812 23166
rect 35756 23102 35758 23154
rect 35810 23102 35812 23154
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34860 22146 34916 22158
rect 34860 22094 34862 22146
rect 34914 22094 34916 22146
rect 34748 21812 34804 21822
rect 34636 21810 34804 21812
rect 34636 21758 34750 21810
rect 34802 21758 34804 21810
rect 34636 21756 34804 21758
rect 34748 21746 34804 21756
rect 34524 21588 34580 21644
rect 34524 21532 34692 21588
rect 34412 20750 34414 20802
rect 34466 20750 34468 20802
rect 34412 20692 34468 20750
rect 34524 20804 34580 20814
rect 34524 20710 34580 20748
rect 34636 20802 34692 21532
rect 34636 20750 34638 20802
rect 34690 20750 34692 20802
rect 34636 20738 34692 20750
rect 34412 20626 34468 20636
rect 34860 20244 34916 22094
rect 34972 20916 35028 22204
rect 35196 22484 35252 22494
rect 35196 22258 35252 22428
rect 35196 22206 35198 22258
rect 35250 22206 35252 22258
rect 35196 22194 35252 22206
rect 35532 22372 35588 22382
rect 35756 22372 35812 23102
rect 36204 23156 36260 23166
rect 36204 23062 36260 23100
rect 35588 22316 35812 22372
rect 35868 22932 35924 22942
rect 36316 22932 36372 24670
rect 36428 22932 36484 22942
rect 36316 22930 36484 22932
rect 36316 22878 36430 22930
rect 36482 22878 36484 22930
rect 36316 22876 36484 22878
rect 35084 21588 35140 21598
rect 35084 21494 35140 21532
rect 35532 21474 35588 22316
rect 35868 22260 35924 22876
rect 36428 22866 36484 22876
rect 35644 22204 35868 22260
rect 35644 22146 35700 22204
rect 35868 22166 35924 22204
rect 35644 22094 35646 22146
rect 35698 22094 35700 22146
rect 35644 22082 35700 22094
rect 36764 21812 36820 21822
rect 36876 21812 36932 30604
rect 37436 30434 37492 30828
rect 37660 30772 37716 32284
rect 37772 30996 37828 32510
rect 37884 31780 37940 34188
rect 37884 31714 37940 31724
rect 37996 34130 38052 34142
rect 37996 34078 37998 34130
rect 38050 34078 38052 34130
rect 37996 34020 38052 34078
rect 37884 30996 37940 31006
rect 37772 30994 37940 30996
rect 37772 30942 37886 30994
rect 37938 30942 37940 30994
rect 37772 30940 37940 30942
rect 37884 30930 37940 30940
rect 37436 30382 37438 30434
rect 37490 30382 37492 30434
rect 37436 30370 37492 30382
rect 37548 30716 37716 30772
rect 37324 30212 37380 30222
rect 37100 29986 37156 29998
rect 37100 29934 37102 29986
rect 37154 29934 37156 29986
rect 37100 28980 37156 29934
rect 37100 28914 37156 28924
rect 37212 29428 37268 29438
rect 37212 27186 37268 29372
rect 37212 27134 37214 27186
rect 37266 27134 37268 27186
rect 37212 27122 37268 27134
rect 37324 27076 37380 30156
rect 37436 28418 37492 28430
rect 37436 28366 37438 28418
rect 37490 28366 37492 28418
rect 37436 27858 37492 28366
rect 37436 27806 37438 27858
rect 37490 27806 37492 27858
rect 37436 27794 37492 27806
rect 37436 27300 37492 27310
rect 37436 27206 37492 27244
rect 37324 26908 37380 27020
rect 37324 26852 37492 26908
rect 37100 26516 37156 26526
rect 37100 26290 37156 26460
rect 37100 26238 37102 26290
rect 37154 26238 37156 26290
rect 37100 26226 37156 26238
rect 37324 25618 37380 25630
rect 37324 25566 37326 25618
rect 37378 25566 37380 25618
rect 37212 24722 37268 24734
rect 37212 24670 37214 24722
rect 37266 24670 37268 24722
rect 37212 24050 37268 24670
rect 37212 23998 37214 24050
rect 37266 23998 37268 24050
rect 37212 23986 37268 23998
rect 36988 23828 37044 23838
rect 36988 23734 37044 23772
rect 37212 23716 37268 23726
rect 37324 23716 37380 25566
rect 37436 25172 37492 26852
rect 37436 25106 37492 25116
rect 37436 24500 37492 24510
rect 37436 23938 37492 24444
rect 37436 23886 37438 23938
rect 37490 23886 37492 23938
rect 37436 23874 37492 23886
rect 37268 23660 37380 23716
rect 37212 23622 37268 23660
rect 37100 23268 37156 23278
rect 37100 22594 37156 23212
rect 37100 22542 37102 22594
rect 37154 22542 37156 22594
rect 37100 22530 37156 22542
rect 37436 22596 37492 22606
rect 37548 22596 37604 30716
rect 37884 30212 37940 30222
rect 37884 30118 37940 30156
rect 37996 29876 38052 33964
rect 38108 33908 38164 34972
rect 38220 34962 38276 34972
rect 38444 34356 38500 37660
rect 38556 37490 38612 38556
rect 38556 37438 38558 37490
rect 38610 37438 38612 37490
rect 38556 37426 38612 37438
rect 38556 37044 38612 37054
rect 38556 36482 38612 36988
rect 38556 36430 38558 36482
rect 38610 36430 38612 36482
rect 38556 36418 38612 36430
rect 38556 36258 38612 36270
rect 38556 36206 38558 36258
rect 38610 36206 38612 36258
rect 38556 35698 38612 36206
rect 38556 35646 38558 35698
rect 38610 35646 38612 35698
rect 38556 35634 38612 35646
rect 38668 35252 38724 39454
rect 38892 38836 38948 38846
rect 38892 37828 38948 38780
rect 39004 38050 39060 40124
rect 39452 39508 39508 39518
rect 39452 39506 40068 39508
rect 39452 39454 39454 39506
rect 39506 39454 40068 39506
rect 39452 39452 40068 39454
rect 39452 39442 39508 39452
rect 39452 39060 39508 39070
rect 39452 38966 39508 39004
rect 39116 38836 39172 38846
rect 39676 38836 39732 38846
rect 39116 38834 39396 38836
rect 39116 38782 39118 38834
rect 39170 38782 39396 38834
rect 39116 38780 39396 38782
rect 39116 38770 39172 38780
rect 39004 37998 39006 38050
rect 39058 37998 39060 38050
rect 39004 37986 39060 37998
rect 39228 38612 39284 38622
rect 38892 37772 39060 37828
rect 38892 37266 38948 37278
rect 38892 37214 38894 37266
rect 38946 37214 38948 37266
rect 38892 37156 38948 37214
rect 38892 37090 38948 37100
rect 38668 35186 38724 35196
rect 38668 34916 38724 34926
rect 39004 34916 39060 37772
rect 39228 37380 39284 38556
rect 39116 37324 39284 37380
rect 39116 35922 39172 37324
rect 39228 37156 39284 37166
rect 39228 36370 39284 37100
rect 39228 36318 39230 36370
rect 39282 36318 39284 36370
rect 39228 36306 39284 36318
rect 39340 36596 39396 38780
rect 39676 38742 39732 38780
rect 39116 35870 39118 35922
rect 39170 35870 39172 35922
rect 39116 35858 39172 35870
rect 39340 35698 39396 36540
rect 39452 38052 39508 38062
rect 39452 36484 39508 37996
rect 40012 38050 40068 39452
rect 41580 38834 41636 38846
rect 41580 38782 41582 38834
rect 41634 38782 41636 38834
rect 41132 38722 41188 38734
rect 41132 38670 41134 38722
rect 41186 38670 41188 38722
rect 40908 38612 40964 38622
rect 40908 38518 40964 38556
rect 40012 37998 40014 38050
rect 40066 37998 40068 38050
rect 40012 37986 40068 37998
rect 40908 38052 40964 38062
rect 40908 37958 40964 37996
rect 40348 37380 40404 37390
rect 40908 37380 40964 37390
rect 40348 37378 40964 37380
rect 40348 37326 40350 37378
rect 40402 37326 40910 37378
rect 40962 37326 40964 37378
rect 40348 37324 40964 37326
rect 40348 37314 40404 37324
rect 40908 37314 40964 37324
rect 40012 37268 40068 37278
rect 40012 37174 40068 37212
rect 39564 37154 39620 37166
rect 39564 37102 39566 37154
rect 39618 37102 39620 37154
rect 39564 37044 39620 37102
rect 40348 37156 40404 37166
rect 40684 37156 40740 37166
rect 40404 37100 40516 37156
rect 40348 37090 40404 37100
rect 39564 36978 39620 36988
rect 40460 37044 40516 37100
rect 39788 36484 39844 36494
rect 39452 36482 39732 36484
rect 39452 36430 39454 36482
rect 39506 36430 39732 36482
rect 39452 36428 39732 36430
rect 39452 36418 39508 36428
rect 39340 35646 39342 35698
rect 39394 35646 39396 35698
rect 39340 35634 39396 35646
rect 39452 35140 39508 35150
rect 39116 34916 39172 34926
rect 39004 34914 39172 34916
rect 39004 34862 39118 34914
rect 39170 34862 39172 34914
rect 39004 34860 39172 34862
rect 38668 34822 38724 34860
rect 38444 34300 38724 34356
rect 38332 34244 38388 34254
rect 38108 33842 38164 33852
rect 38220 34242 38388 34244
rect 38220 34190 38334 34242
rect 38386 34190 38388 34242
rect 38220 34188 38388 34190
rect 38108 33684 38164 33694
rect 38108 32786 38164 33628
rect 38220 33124 38276 34188
rect 38332 34178 38388 34188
rect 38332 33908 38388 33918
rect 38332 33234 38388 33852
rect 38668 33348 38724 34300
rect 39116 34244 39172 34860
rect 39452 34914 39508 35084
rect 39452 34862 39454 34914
rect 39506 34862 39508 34914
rect 39452 34850 39508 34862
rect 39676 34804 39732 36428
rect 39788 36390 39844 36428
rect 40124 36260 40180 36270
rect 40124 36166 40180 36204
rect 39900 36036 39956 36046
rect 39900 35924 39956 35980
rect 39900 35922 40180 35924
rect 39900 35870 39902 35922
rect 39954 35870 40180 35922
rect 39900 35868 40180 35870
rect 39900 35858 39956 35868
rect 39116 34178 39172 34188
rect 39340 34692 39396 34702
rect 39004 34132 39060 34142
rect 38892 34020 38948 34030
rect 38892 33926 38948 33964
rect 38668 33282 38724 33292
rect 38332 33182 38334 33234
rect 38386 33182 38388 33234
rect 38332 33170 38388 33182
rect 38220 33058 38276 33068
rect 38108 32734 38110 32786
rect 38162 32734 38164 32786
rect 38108 30436 38164 32734
rect 38332 32564 38388 32574
rect 38332 32470 38388 32508
rect 38780 32562 38836 32574
rect 38780 32510 38782 32562
rect 38834 32510 38836 32562
rect 38780 32340 38836 32510
rect 38780 32274 38836 32284
rect 38892 32452 38948 32462
rect 38892 31778 38948 32396
rect 39004 31948 39060 34076
rect 39116 33348 39172 33358
rect 39116 32786 39172 33292
rect 39116 32734 39118 32786
rect 39170 32734 39172 32786
rect 39116 32722 39172 32734
rect 39004 31892 39172 31948
rect 38892 31726 38894 31778
rect 38946 31726 38948 31778
rect 38108 30370 38164 30380
rect 38220 30996 38276 31006
rect 38220 30098 38276 30940
rect 38220 30046 38222 30098
rect 38274 30046 38276 30098
rect 38220 30034 38276 30046
rect 38668 30098 38724 30110
rect 38668 30046 38670 30098
rect 38722 30046 38724 30098
rect 37660 29820 38052 29876
rect 37660 26908 37716 29820
rect 38220 29540 38276 29550
rect 37772 29316 37828 29326
rect 37772 29314 38164 29316
rect 37772 29262 37774 29314
rect 37826 29262 38164 29314
rect 37772 29260 38164 29262
rect 37772 29250 37828 29260
rect 37772 29092 37828 29102
rect 37772 27300 37828 29036
rect 37772 27234 37828 27244
rect 37884 27860 37940 27870
rect 37884 27074 37940 27804
rect 38108 27748 38164 29260
rect 38220 28644 38276 29484
rect 38444 28644 38500 28654
rect 38220 28642 38612 28644
rect 38220 28590 38446 28642
rect 38498 28590 38612 28642
rect 38220 28588 38612 28590
rect 38444 28578 38500 28588
rect 38332 27858 38388 27870
rect 38332 27806 38334 27858
rect 38386 27806 38388 27858
rect 38108 27692 38276 27748
rect 37884 27022 37886 27074
rect 37938 27022 37940 27074
rect 37660 26852 37828 26908
rect 37772 26290 37828 26852
rect 37772 26238 37774 26290
rect 37826 26238 37828 26290
rect 37772 25620 37828 26238
rect 37884 26180 37940 27022
rect 38220 27076 38276 27692
rect 38332 27298 38388 27806
rect 38332 27246 38334 27298
rect 38386 27246 38388 27298
rect 38332 27234 38388 27246
rect 38108 26964 38164 27002
rect 38220 26982 38276 27020
rect 38556 27074 38612 28588
rect 38668 27636 38724 30046
rect 38892 30100 38948 31726
rect 39004 31668 39060 31678
rect 39004 30994 39060 31612
rect 39004 30942 39006 30994
rect 39058 30942 39060 30994
rect 39004 30930 39060 30942
rect 38892 30034 38948 30044
rect 39004 29988 39060 29998
rect 39116 29988 39172 31892
rect 39004 29986 39172 29988
rect 39004 29934 39006 29986
rect 39058 29934 39172 29986
rect 39004 29932 39172 29934
rect 39340 30210 39396 34636
rect 39452 34356 39508 34366
rect 39452 34262 39508 34300
rect 39676 34132 39732 34748
rect 39788 35252 39844 35262
rect 39788 34804 39844 35196
rect 40124 34914 40180 35868
rect 40124 34862 40126 34914
rect 40178 34862 40180 34914
rect 40124 34850 40180 34862
rect 40012 34804 40068 34814
rect 39788 34802 40012 34804
rect 39788 34750 39790 34802
rect 39842 34750 40012 34802
rect 39788 34748 40012 34750
rect 39788 34738 39844 34748
rect 40012 34244 40068 34748
rect 40460 34802 40516 36988
rect 40684 36370 40740 37100
rect 40684 36318 40686 36370
rect 40738 36318 40740 36370
rect 40684 36306 40740 36318
rect 41020 36370 41076 36382
rect 41020 36318 41022 36370
rect 41074 36318 41076 36370
rect 41020 35812 41076 36318
rect 41132 36260 41188 38670
rect 41356 38722 41412 38734
rect 41356 38670 41358 38722
rect 41410 38670 41412 38722
rect 41244 37380 41300 37390
rect 41244 37266 41300 37324
rect 41244 37214 41246 37266
rect 41298 37214 41300 37266
rect 41244 37202 41300 37214
rect 41356 37268 41412 38670
rect 41356 37202 41412 37212
rect 41356 37044 41412 37054
rect 41412 36988 41524 37044
rect 41356 36978 41412 36988
rect 41356 36260 41412 36270
rect 41132 36204 41356 36260
rect 41132 35812 41188 35822
rect 41020 35810 41188 35812
rect 41020 35758 41134 35810
rect 41186 35758 41188 35810
rect 41020 35756 41188 35758
rect 41020 34914 41076 35756
rect 41132 35746 41188 35756
rect 41020 34862 41022 34914
rect 41074 34862 41076 34914
rect 41020 34850 41076 34862
rect 40460 34750 40462 34802
rect 40514 34750 40516 34802
rect 40460 34356 40516 34750
rect 40460 34290 40516 34300
rect 41132 34692 41188 34702
rect 41132 34354 41188 34636
rect 41132 34302 41134 34354
rect 41186 34302 41188 34354
rect 41132 34290 41188 34302
rect 40012 34188 40292 34244
rect 39788 34132 39844 34142
rect 39676 34076 39788 34132
rect 39788 34038 39844 34076
rect 40236 34130 40292 34188
rect 40236 34078 40238 34130
rect 40290 34078 40292 34130
rect 40236 34066 40292 34078
rect 40908 34132 40964 34142
rect 41356 34132 41412 36204
rect 41468 35810 41524 36988
rect 41468 35758 41470 35810
rect 41522 35758 41524 35810
rect 41468 35746 41524 35758
rect 41468 35476 41524 35486
rect 41468 35026 41524 35420
rect 41468 34974 41470 35026
rect 41522 34974 41524 35026
rect 41468 34580 41524 34974
rect 41580 34804 41636 38782
rect 41804 38836 41860 38846
rect 41804 38834 41972 38836
rect 41804 38782 41806 38834
rect 41858 38782 41972 38834
rect 41804 38780 41972 38782
rect 41804 38770 41860 38780
rect 41692 38722 41748 38734
rect 41692 38670 41694 38722
rect 41746 38670 41748 38722
rect 41692 37490 41748 38670
rect 41692 37438 41694 37490
rect 41746 37438 41748 37490
rect 41692 37426 41748 37438
rect 41916 35924 41972 38780
rect 43148 38162 43204 38174
rect 43148 38110 43150 38162
rect 43202 38110 43204 38162
rect 42476 38050 42532 38062
rect 42476 37998 42478 38050
rect 42530 37998 42532 38050
rect 42028 37156 42084 37166
rect 42028 37062 42084 37100
rect 41916 34914 41972 35868
rect 41916 34862 41918 34914
rect 41970 34862 41972 34914
rect 41916 34850 41972 34862
rect 42364 36932 42420 36942
rect 42364 35588 42420 36876
rect 42476 36596 42532 37998
rect 42476 36530 42532 36540
rect 42700 38050 42756 38062
rect 42700 37998 42702 38050
rect 42754 37998 42756 38050
rect 42700 36484 42756 37998
rect 43148 37266 43204 38110
rect 43708 37940 43764 37950
rect 43148 37214 43150 37266
rect 43202 37214 43204 37266
rect 43148 37202 43204 37214
rect 43260 37938 43764 37940
rect 43260 37886 43710 37938
rect 43762 37886 43764 37938
rect 43260 37884 43764 37886
rect 42700 36418 42756 36428
rect 42812 37042 42868 37054
rect 42812 36990 42814 37042
rect 42866 36990 42868 37042
rect 42700 35698 42756 35710
rect 42700 35646 42702 35698
rect 42754 35646 42756 35698
rect 42700 35588 42756 35646
rect 42364 35586 42756 35588
rect 42364 35534 42366 35586
rect 42418 35534 42756 35586
rect 42364 35532 42756 35534
rect 41580 34738 41636 34748
rect 41468 34524 41860 34580
rect 41468 34132 41524 34142
rect 41356 34130 41524 34132
rect 41356 34078 41470 34130
rect 41522 34078 41524 34130
rect 41356 34076 41524 34078
rect 40908 34038 40964 34076
rect 41468 34066 41524 34076
rect 41804 34130 41860 34524
rect 41804 34078 41806 34130
rect 41858 34078 41860 34130
rect 41804 34066 41860 34078
rect 41356 33348 41412 33358
rect 41132 33346 41412 33348
rect 41132 33294 41358 33346
rect 41410 33294 41412 33346
rect 41132 33292 41412 33294
rect 40796 33236 40852 33246
rect 41020 33236 41076 33246
rect 40796 33234 41076 33236
rect 40796 33182 40798 33234
rect 40850 33182 41022 33234
rect 41074 33182 41076 33234
rect 40796 33180 41076 33182
rect 40796 33170 40852 33180
rect 41020 33170 41076 33180
rect 41020 32788 41076 32798
rect 41132 32788 41188 33292
rect 41356 33282 41412 33292
rect 41804 33346 41860 33358
rect 41804 33294 41806 33346
rect 41858 33294 41860 33346
rect 41020 32786 41188 32788
rect 41020 32734 41022 32786
rect 41074 32734 41188 32786
rect 41020 32732 41188 32734
rect 39564 32564 39620 32574
rect 39564 32470 39620 32508
rect 41020 31948 41076 32732
rect 41804 32450 41860 33294
rect 41804 32398 41806 32450
rect 41858 32398 41860 32450
rect 41804 32386 41860 32398
rect 42028 33122 42084 33134
rect 42028 33070 42030 33122
rect 42082 33070 42084 33122
rect 40908 31892 41076 31948
rect 41580 31892 41636 31902
rect 39452 31780 39508 31790
rect 39452 31666 39508 31724
rect 39452 31614 39454 31666
rect 39506 31614 39508 31666
rect 39452 31602 39508 31614
rect 39676 31778 39732 31790
rect 39676 31726 39678 31778
rect 39730 31726 39732 31778
rect 39564 31556 39620 31566
rect 39564 30994 39620 31500
rect 39564 30942 39566 30994
rect 39618 30942 39620 30994
rect 39564 30930 39620 30942
rect 39676 30884 39732 31726
rect 40236 31556 40292 31566
rect 40236 31462 40292 31500
rect 39900 30884 39956 30894
rect 39676 30882 39956 30884
rect 39676 30830 39902 30882
rect 39954 30830 39956 30882
rect 39676 30828 39956 30830
rect 39340 30158 39342 30210
rect 39394 30158 39396 30210
rect 39004 29876 39060 29932
rect 38780 29820 39060 29876
rect 38780 28084 38836 29820
rect 38780 28018 38836 28028
rect 38892 29652 38948 29662
rect 38668 27570 38724 27580
rect 38556 27022 38558 27074
rect 38610 27022 38612 27074
rect 38556 27010 38612 27022
rect 38892 27074 38948 29596
rect 39340 29428 39396 30158
rect 39900 29652 39956 30828
rect 39900 29586 39956 29596
rect 40796 30210 40852 30222
rect 40796 30158 40798 30210
rect 40850 30158 40852 30210
rect 39340 29362 39396 29372
rect 40124 29204 40180 29214
rect 40124 29202 40292 29204
rect 40124 29150 40126 29202
rect 40178 29150 40292 29202
rect 40124 29148 40292 29150
rect 40124 29138 40180 29148
rect 38892 27022 38894 27074
rect 38946 27022 38948 27074
rect 38892 27010 38948 27022
rect 39004 28980 39060 28990
rect 38108 26898 38164 26908
rect 39004 26964 39060 28924
rect 39676 28418 39732 28430
rect 39676 28366 39678 28418
rect 39730 28366 39732 28418
rect 39676 27860 39732 28366
rect 40012 27860 40068 27870
rect 39676 27804 40012 27860
rect 39564 27748 39620 27758
rect 39620 27692 39732 27748
rect 39564 27654 39620 27692
rect 39116 27636 39172 27646
rect 39116 27634 39508 27636
rect 39116 27582 39118 27634
rect 39170 27582 39508 27634
rect 39116 27580 39508 27582
rect 39116 27570 39172 27580
rect 39340 27412 39396 27422
rect 38780 26516 38836 26526
rect 38780 26290 38836 26460
rect 38780 26238 38782 26290
rect 38834 26238 38836 26290
rect 38780 26226 38836 26238
rect 38220 26180 38276 26190
rect 37884 26178 38276 26180
rect 37884 26126 38222 26178
rect 38274 26126 38276 26178
rect 37884 26124 38276 26126
rect 39004 26180 39060 26908
rect 39228 27076 39284 27086
rect 39228 26962 39284 27020
rect 39228 26910 39230 26962
rect 39282 26910 39284 26962
rect 39228 26898 39284 26910
rect 39116 26180 39172 26190
rect 39004 26178 39172 26180
rect 39004 26126 39118 26178
rect 39170 26126 39172 26178
rect 39004 26124 39172 26126
rect 38220 26114 38276 26124
rect 39116 26114 39172 26124
rect 37772 25554 37828 25564
rect 37772 25284 37828 25294
rect 37772 25282 38052 25284
rect 37772 25230 37774 25282
rect 37826 25230 38052 25282
rect 37772 25228 38052 25230
rect 37772 25218 37828 25228
rect 37436 22594 37604 22596
rect 37436 22542 37438 22594
rect 37490 22542 37604 22594
rect 37436 22540 37604 22542
rect 37660 25172 37716 25182
rect 37660 24164 37716 25116
rect 37436 22530 37492 22540
rect 37660 22258 37716 24108
rect 37884 24610 37940 24622
rect 37884 24558 37886 24610
rect 37938 24558 37940 24610
rect 37772 23940 37828 23950
rect 37772 23846 37828 23884
rect 37884 23828 37940 24558
rect 37884 23762 37940 23772
rect 37996 22484 38052 25228
rect 38108 25282 38164 25294
rect 38108 25230 38110 25282
rect 38162 25230 38164 25282
rect 38108 24500 38164 25230
rect 38444 25282 38500 25294
rect 38444 25230 38446 25282
rect 38498 25230 38500 25282
rect 38332 24724 38388 24734
rect 38332 24630 38388 24668
rect 38444 24500 38500 25230
rect 38108 24434 38164 24444
rect 38332 24444 38444 24500
rect 38332 23268 38388 24444
rect 38444 24434 38500 24444
rect 38780 25282 38836 25294
rect 39116 25284 39172 25294
rect 38780 25230 38782 25282
rect 38834 25230 38836 25282
rect 38780 24276 38836 25230
rect 38780 24210 38836 24220
rect 38892 25282 39172 25284
rect 38892 25230 39118 25282
rect 39170 25230 39172 25282
rect 38892 25228 39172 25230
rect 38444 24164 38500 24174
rect 38444 24070 38500 24108
rect 38780 23940 38836 23950
rect 38556 23938 38836 23940
rect 38556 23886 38782 23938
rect 38834 23886 38836 23938
rect 38556 23884 38836 23886
rect 38556 23716 38612 23884
rect 38780 23874 38836 23884
rect 38332 23212 38500 23268
rect 37660 22206 37662 22258
rect 37714 22206 37716 22258
rect 37660 22194 37716 22206
rect 37772 22428 38052 22484
rect 36092 21810 36932 21812
rect 36092 21758 36766 21810
rect 36818 21758 36932 21810
rect 36092 21756 36932 21758
rect 35980 21700 36036 21710
rect 35980 21606 36036 21644
rect 35532 21422 35534 21474
rect 35586 21422 35588 21474
rect 35532 21410 35588 21422
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 20916 35252 20926
rect 36092 20916 36148 21756
rect 36764 21746 36820 21756
rect 36204 21586 36260 21598
rect 36204 21534 36206 21586
rect 36258 21534 36260 21586
rect 36204 21364 36260 21534
rect 36204 21298 36260 21308
rect 37660 21586 37716 21598
rect 37660 21534 37662 21586
rect 37714 21534 37716 21586
rect 34972 20914 35252 20916
rect 34972 20862 35198 20914
rect 35250 20862 35252 20914
rect 34972 20860 35252 20862
rect 34860 20178 34916 20188
rect 34524 20020 34580 20030
rect 35084 20020 35140 20030
rect 34300 20018 34580 20020
rect 34300 19966 34526 20018
rect 34578 19966 34580 20018
rect 34300 19964 34580 19966
rect 34076 19618 34132 19628
rect 34188 19794 34244 19806
rect 34188 19742 34190 19794
rect 34242 19742 34244 19794
rect 34076 19012 34132 19022
rect 33740 17602 33796 17612
rect 33852 19010 34132 19012
rect 33852 18958 34078 19010
rect 34130 18958 34132 19010
rect 33852 18956 34132 18958
rect 33740 16772 33796 16782
rect 33740 16098 33796 16716
rect 33740 16046 33742 16098
rect 33794 16046 33796 16098
rect 33740 16034 33796 16046
rect 33852 15540 33908 18956
rect 34076 18946 34132 18956
rect 34076 17668 34132 17678
rect 34188 17668 34244 19742
rect 34076 17666 34244 17668
rect 34076 17614 34078 17666
rect 34130 17614 34244 17666
rect 34076 17612 34244 17614
rect 34076 17602 34132 17612
rect 34188 16772 34244 17612
rect 34300 16884 34356 19964
rect 34524 19954 34580 19964
rect 34636 20018 35140 20020
rect 34636 19966 35086 20018
rect 35138 19966 35140 20018
rect 34636 19964 35140 19966
rect 34636 19794 34692 19964
rect 35084 19954 35140 19964
rect 34636 19742 34638 19794
rect 34690 19742 34692 19794
rect 34636 19730 34692 19742
rect 34748 19794 34804 19806
rect 35196 19796 35252 20860
rect 35644 20860 36260 20916
rect 35644 20802 35700 20860
rect 35644 20750 35646 20802
rect 35698 20750 35700 20802
rect 35644 20738 35700 20750
rect 35980 20692 36036 20702
rect 35980 20598 36036 20636
rect 35756 20356 35812 20366
rect 34748 19742 34750 19794
rect 34802 19742 34804 19794
rect 34412 19124 34468 19134
rect 34412 17890 34468 19068
rect 34524 19122 34580 19134
rect 34524 19070 34526 19122
rect 34578 19070 34580 19122
rect 34524 18340 34580 19070
rect 34748 19124 34804 19742
rect 34748 19058 34804 19068
rect 34972 19740 35252 19796
rect 35532 20018 35588 20030
rect 35532 19966 35534 20018
rect 35586 19966 35588 20018
rect 34972 18900 35028 19740
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35532 19348 35588 19966
rect 35308 19292 35588 19348
rect 34636 18844 35028 18900
rect 35084 19234 35140 19246
rect 35084 19182 35086 19234
rect 35138 19182 35140 19234
rect 34636 18450 34692 18844
rect 34636 18398 34638 18450
rect 34690 18398 34692 18450
rect 34636 18386 34692 18398
rect 34748 18452 34804 18462
rect 34524 18274 34580 18284
rect 34748 18338 34804 18396
rect 34748 18286 34750 18338
rect 34802 18286 34804 18338
rect 34412 17838 34414 17890
rect 34466 17838 34468 17890
rect 34412 17826 34468 17838
rect 34748 17444 34804 18286
rect 34972 18452 35028 18462
rect 34972 18116 35028 18396
rect 34972 18050 35028 18060
rect 35084 17892 35140 19182
rect 35308 18452 35364 19292
rect 35644 19234 35700 19246
rect 35644 19182 35646 19234
rect 35698 19182 35700 19234
rect 35308 18386 35364 18396
rect 35420 19124 35476 19134
rect 35420 18450 35476 19068
rect 35420 18398 35422 18450
rect 35474 18398 35476 18450
rect 35420 18386 35476 18398
rect 35532 19012 35588 19022
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35084 17826 35140 17836
rect 34972 17778 35028 17790
rect 34972 17726 34974 17778
rect 35026 17726 35028 17778
rect 34972 17668 35028 17726
rect 34972 17556 35028 17612
rect 35420 17668 35476 17678
rect 35532 17668 35588 18956
rect 35644 18676 35700 19182
rect 35756 19012 35812 20300
rect 36092 20132 36148 20142
rect 36092 20038 36148 20076
rect 35980 20018 36036 20030
rect 35980 19966 35982 20018
rect 36034 19966 36036 20018
rect 35756 18946 35812 18956
rect 35868 19124 35924 19134
rect 35644 18610 35700 18620
rect 35868 18452 35924 19068
rect 35420 17666 35588 17668
rect 35420 17614 35422 17666
rect 35474 17614 35588 17666
rect 35420 17612 35588 17614
rect 35644 18396 35924 18452
rect 35420 17602 35476 17612
rect 35308 17556 35364 17566
rect 34972 17500 35308 17556
rect 35308 17490 35364 17500
rect 34748 17388 34916 17444
rect 34748 16884 34804 16894
rect 34300 16828 34468 16884
rect 33964 16660 34020 16670
rect 33964 16658 34132 16660
rect 33964 16606 33966 16658
rect 34018 16606 34132 16658
rect 33964 16604 34132 16606
rect 33964 16594 34020 16604
rect 33852 15474 33908 15484
rect 33628 15092 33796 15148
rect 33292 14578 33348 14588
rect 33180 14532 33236 14542
rect 33180 14438 33236 14476
rect 32956 14420 33012 14430
rect 32956 14326 33012 14364
rect 32620 13692 32900 13748
rect 33628 13748 33684 13758
rect 32508 12962 32564 12974
rect 32508 12910 32510 12962
rect 32562 12910 32564 12962
rect 32508 12628 32564 12910
rect 32508 12562 32564 12572
rect 32284 12460 32452 12516
rect 32172 12180 32228 12190
rect 32060 12124 32172 12180
rect 32172 12114 32228 12124
rect 32172 11508 32228 11518
rect 32172 11414 32228 11452
rect 32284 11284 32340 12460
rect 32508 12404 32564 12414
rect 32396 12348 32508 12404
rect 32396 12178 32452 12348
rect 32508 12338 32564 12348
rect 32396 12126 32398 12178
rect 32450 12126 32452 12178
rect 32396 12114 32452 12126
rect 32620 11788 32676 13692
rect 33628 13654 33684 13692
rect 33068 13636 33124 13646
rect 32732 13634 33124 13636
rect 32732 13582 33070 13634
rect 33122 13582 33124 13634
rect 32732 13580 33124 13582
rect 32732 12964 32788 13580
rect 33068 13570 33124 13580
rect 33740 13188 33796 15092
rect 33852 14756 33908 14766
rect 33852 14662 33908 14700
rect 33964 13860 34020 13870
rect 33964 13766 34020 13804
rect 33628 13132 33796 13188
rect 33628 12964 33684 13132
rect 32732 12870 32788 12908
rect 33516 12962 33684 12964
rect 33516 12910 33630 12962
rect 33682 12910 33684 12962
rect 33516 12908 33684 12910
rect 33180 12850 33236 12862
rect 33180 12798 33182 12850
rect 33234 12798 33236 12850
rect 33180 12740 33236 12798
rect 33180 12674 33236 12684
rect 32844 12180 32900 12190
rect 33068 12180 33124 12190
rect 32900 12178 33124 12180
rect 32900 12126 33070 12178
rect 33122 12126 33124 12178
rect 32900 12124 33124 12126
rect 32844 12114 32900 12124
rect 33068 12114 33124 12124
rect 33180 12180 33236 12190
rect 33068 11956 33124 11966
rect 32620 11732 33012 11788
rect 32284 11228 32676 11284
rect 32620 9940 32676 11228
rect 32956 11172 33012 11732
rect 32956 11106 33012 11116
rect 31724 9268 31780 9278
rect 31724 9174 31780 9212
rect 31276 8930 31668 8932
rect 31276 8878 31278 8930
rect 31330 8878 31668 8930
rect 31276 8876 31668 8878
rect 31276 8866 31332 8876
rect 30716 8418 30772 8428
rect 30604 8372 30660 8382
rect 30604 8148 30660 8316
rect 31836 8372 31892 8382
rect 30044 8082 30100 8092
rect 30156 8146 30660 8148
rect 30156 8094 30606 8146
rect 30658 8094 30660 8146
rect 30156 8092 30660 8094
rect 30156 7586 30212 8092
rect 30156 7534 30158 7586
rect 30210 7534 30212 7586
rect 30156 7522 30212 7534
rect 29484 6690 29652 6692
rect 29484 6638 29486 6690
rect 29538 6638 29652 6690
rect 29484 6636 29652 6638
rect 30156 7364 30212 7374
rect 30156 6692 30212 7308
rect 29484 6626 29540 6636
rect 30156 6598 30212 6636
rect 30604 6690 30660 8092
rect 30828 8258 30884 8270
rect 30828 8206 30830 8258
rect 30882 8206 30884 8258
rect 30828 8148 30884 8206
rect 31276 8260 31332 8270
rect 31276 8166 31332 8204
rect 31836 8258 31892 8316
rect 31836 8206 31838 8258
rect 31890 8206 31892 8258
rect 31836 8194 31892 8206
rect 30828 8082 30884 8092
rect 31948 8148 32004 9884
rect 32396 9938 32676 9940
rect 32396 9886 32622 9938
rect 32674 9886 32676 9938
rect 32396 9884 32676 9886
rect 32060 9828 32116 9838
rect 32060 9734 32116 9772
rect 32060 9268 32116 9278
rect 32060 9174 32116 9212
rect 32396 9266 32452 9884
rect 32620 9874 32676 9884
rect 33068 9828 33124 11900
rect 33180 11508 33236 12124
rect 33516 12068 33572 12908
rect 33628 12898 33684 12908
rect 33740 12964 33796 12974
rect 33628 12628 33684 12638
rect 33628 12178 33684 12572
rect 33628 12126 33630 12178
rect 33682 12126 33684 12178
rect 33628 12114 33684 12126
rect 33740 12290 33796 12908
rect 33740 12238 33742 12290
rect 33794 12238 33796 12290
rect 33404 12012 33572 12068
rect 33404 11956 33460 12012
rect 33740 11956 33796 12238
rect 33964 12962 34020 12974
rect 33964 12910 33966 12962
rect 34018 12910 34020 12962
rect 33404 11890 33460 11900
rect 33516 11900 33796 11956
rect 33852 12180 33908 12190
rect 33180 10834 33236 11452
rect 33180 10782 33182 10834
rect 33234 10782 33236 10834
rect 33180 10770 33236 10782
rect 33292 11732 33348 11742
rect 33292 10834 33348 11676
rect 33516 11396 33572 11900
rect 33292 10782 33294 10834
rect 33346 10782 33348 10834
rect 33292 10770 33348 10782
rect 33404 11394 33572 11396
rect 33404 11342 33518 11394
rect 33570 11342 33572 11394
rect 33404 11340 33572 11342
rect 33404 10834 33460 11340
rect 33516 11330 33572 11340
rect 33740 11732 33796 11742
rect 33404 10782 33406 10834
rect 33458 10782 33460 10834
rect 33404 10770 33460 10782
rect 33516 11172 33572 11182
rect 33404 10612 33460 10622
rect 33292 9828 33348 9838
rect 33068 9826 33348 9828
rect 33068 9774 33294 9826
rect 33346 9774 33348 9826
rect 33068 9772 33348 9774
rect 33292 9762 33348 9772
rect 32956 9714 33012 9726
rect 32956 9662 32958 9714
rect 33010 9662 33012 9714
rect 32956 9604 33012 9662
rect 32396 9214 32398 9266
rect 32450 9214 32452 9266
rect 32396 9202 32452 9214
rect 32508 9548 33012 9604
rect 31948 8082 32004 8092
rect 32396 7700 32452 7710
rect 32508 7700 32564 9548
rect 33404 9266 33460 10556
rect 33404 9214 33406 9266
rect 33458 9214 33460 9266
rect 33404 9202 33460 9214
rect 33180 9044 33236 9054
rect 33516 9044 33572 11116
rect 33628 10498 33684 10510
rect 33628 10446 33630 10498
rect 33682 10446 33684 10498
rect 33628 10276 33684 10446
rect 33740 10500 33796 11676
rect 33852 10724 33908 12124
rect 33964 11506 34020 12910
rect 34076 12852 34132 16604
rect 34188 15314 34244 16716
rect 34300 16658 34356 16670
rect 34300 16606 34302 16658
rect 34354 16606 34356 16658
rect 34300 16548 34356 16606
rect 34300 16482 34356 16492
rect 34188 15262 34190 15314
rect 34242 15262 34244 15314
rect 34188 15250 34244 15262
rect 34412 16324 34468 16828
rect 34412 15314 34468 16268
rect 34412 15262 34414 15314
rect 34466 15262 34468 15314
rect 34412 15250 34468 15262
rect 34524 16882 34804 16884
rect 34524 16830 34750 16882
rect 34802 16830 34804 16882
rect 34524 16828 34804 16830
rect 34524 15148 34580 16828
rect 34748 16818 34804 16828
rect 34860 16660 34916 17388
rect 35196 16772 35252 16782
rect 34748 16604 34916 16660
rect 35084 16770 35252 16772
rect 35084 16718 35198 16770
rect 35250 16718 35252 16770
rect 35084 16716 35252 16718
rect 34524 15092 34692 15148
rect 34188 14532 34244 14542
rect 34188 14530 34356 14532
rect 34188 14478 34190 14530
rect 34242 14478 34356 14530
rect 34188 14476 34356 14478
rect 34188 14466 34244 14476
rect 34188 12852 34244 12862
rect 34076 12850 34244 12852
rect 34076 12798 34190 12850
rect 34242 12798 34244 12850
rect 34076 12796 34244 12798
rect 34188 12786 34244 12796
rect 34076 12404 34132 12414
rect 34076 12066 34132 12348
rect 34076 12014 34078 12066
rect 34130 12014 34132 12066
rect 34076 12002 34132 12014
rect 34300 11788 34356 14476
rect 34412 13746 34468 13758
rect 34412 13694 34414 13746
rect 34466 13694 34468 13746
rect 34412 12068 34468 13694
rect 34636 13076 34692 15092
rect 34412 12002 34468 12012
rect 34524 13020 34692 13076
rect 33964 11454 33966 11506
rect 34018 11454 34020 11506
rect 33964 11442 34020 11454
rect 34076 11732 34356 11788
rect 33852 10668 34020 10724
rect 33852 10500 33908 10510
rect 33740 10498 33908 10500
rect 33740 10446 33854 10498
rect 33906 10446 33908 10498
rect 33740 10444 33908 10446
rect 33852 10434 33908 10444
rect 33964 10276 34020 10668
rect 33628 10220 34020 10276
rect 33628 9828 33684 10220
rect 33628 9762 33684 9772
rect 33740 9826 33796 9838
rect 33740 9774 33742 9826
rect 33794 9774 33796 9826
rect 33180 9042 33572 9044
rect 33180 8990 33182 9042
rect 33234 8990 33572 9042
rect 33180 8988 33572 8990
rect 33180 8978 33236 8988
rect 33628 8484 33684 8494
rect 32396 7698 32564 7700
rect 32396 7646 32398 7698
rect 32450 7646 32564 7698
rect 32396 7644 32564 7646
rect 32844 8148 32900 8158
rect 32396 7634 32452 7644
rect 30604 6638 30606 6690
rect 30658 6638 30660 6690
rect 30604 6626 30660 6638
rect 32844 6690 32900 8092
rect 33628 7474 33684 8428
rect 33628 7422 33630 7474
rect 33682 7422 33684 7474
rect 33628 7410 33684 7422
rect 33740 6914 33796 9774
rect 33964 9716 34020 9726
rect 34076 9716 34132 11732
rect 34524 11394 34580 13020
rect 34748 12628 34804 16604
rect 34860 16098 34916 16110
rect 34860 16046 34862 16098
rect 34914 16046 34916 16098
rect 34860 15202 34916 16046
rect 35084 15988 35140 16716
rect 35196 16706 35252 16716
rect 35532 16660 35588 16670
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35420 16100 35476 16110
rect 35532 16100 35588 16604
rect 35420 16098 35588 16100
rect 35420 16046 35422 16098
rect 35474 16046 35588 16098
rect 35420 16044 35588 16046
rect 35420 16034 35476 16044
rect 35084 15932 35252 15988
rect 34860 15150 34862 15202
rect 34914 15150 34916 15202
rect 34860 15138 34916 15150
rect 34972 15876 35028 15886
rect 34860 14644 34916 14654
rect 34860 14530 34916 14588
rect 34860 14478 34862 14530
rect 34914 14478 34916 14530
rect 34860 13972 34916 14478
rect 34972 14418 35028 15820
rect 34972 14366 34974 14418
rect 35026 14366 35028 14418
rect 34972 14354 35028 14366
rect 35084 15314 35140 15326
rect 35084 15262 35086 15314
rect 35138 15262 35140 15314
rect 34972 13972 35028 13982
rect 34860 13916 34972 13972
rect 34972 13878 35028 13916
rect 35084 13748 35140 15262
rect 35196 15092 35252 15932
rect 35644 15428 35700 18396
rect 35980 18338 36036 19966
rect 36092 19236 36148 19246
rect 36092 19142 36148 19180
rect 35980 18286 35982 18338
rect 36034 18286 36036 18338
rect 35980 18274 36036 18286
rect 35868 18228 35924 18238
rect 35868 17780 35924 18172
rect 35756 17778 35924 17780
rect 35756 17726 35870 17778
rect 35922 17726 35924 17778
rect 35756 17724 35924 17726
rect 35756 16882 35812 17724
rect 35868 17714 35924 17724
rect 36204 17668 36260 20860
rect 36316 20690 36372 20702
rect 36316 20638 36318 20690
rect 36370 20638 36372 20690
rect 36316 17890 36372 20638
rect 36988 20690 37044 20702
rect 36988 20638 36990 20690
rect 37042 20638 37044 20690
rect 36764 20244 36820 20254
rect 36764 20018 36820 20188
rect 36764 19966 36766 20018
rect 36818 19966 36820 20018
rect 36764 19954 36820 19966
rect 36988 19346 37044 20638
rect 37660 20356 37716 21534
rect 37660 20290 37716 20300
rect 36988 19294 36990 19346
rect 37042 19294 37044 19346
rect 36316 17838 36318 17890
rect 36370 17838 36372 17890
rect 36316 17826 36372 17838
rect 36428 19122 36484 19134
rect 36428 19070 36430 19122
rect 36482 19070 36484 19122
rect 36428 17780 36484 19070
rect 36988 19124 37044 19294
rect 36988 19058 37044 19068
rect 37100 20018 37156 20030
rect 37100 19966 37102 20018
rect 37154 19966 37156 20018
rect 36540 19012 36596 19022
rect 36540 18918 36596 18956
rect 37100 19012 37156 19966
rect 37436 19796 37492 19806
rect 37436 19234 37492 19740
rect 37436 19182 37438 19234
rect 37490 19182 37492 19234
rect 37436 19170 37492 19182
rect 37548 19684 37604 19694
rect 37100 18946 37156 18956
rect 36652 18452 36708 18462
rect 36652 18358 36708 18396
rect 37436 18340 37492 18350
rect 37436 18246 37492 18284
rect 36428 17714 36484 17724
rect 36540 17890 36596 17902
rect 36540 17838 36542 17890
rect 36594 17838 36596 17890
rect 35980 17612 36372 17668
rect 35980 17106 36036 17612
rect 36316 17556 36372 17612
rect 36428 17556 36484 17566
rect 36316 17500 36428 17556
rect 36428 17462 36484 17500
rect 35980 17054 35982 17106
rect 36034 17054 36036 17106
rect 35980 17042 36036 17054
rect 35756 16830 35758 16882
rect 35810 16830 35812 16882
rect 35756 16818 35812 16830
rect 36316 16994 36372 17006
rect 36316 16942 36318 16994
rect 36370 16942 36372 16994
rect 36316 16772 36372 16942
rect 36540 16996 36596 17838
rect 37436 17780 37492 17790
rect 37436 17686 37492 17724
rect 36988 17556 37044 17566
rect 36988 17462 37044 17500
rect 36540 16882 36596 16940
rect 36540 16830 36542 16882
rect 36594 16830 36596 16882
rect 36540 16818 36596 16830
rect 37548 17106 37604 19628
rect 37548 17054 37550 17106
rect 37602 17054 37604 17106
rect 36316 16706 36372 16716
rect 35756 16210 35812 16222
rect 35756 16158 35758 16210
rect 35810 16158 35812 16210
rect 35756 16100 35812 16158
rect 35756 16034 35812 16044
rect 37324 15540 37380 15550
rect 37324 15446 37380 15484
rect 35868 15428 35924 15438
rect 35644 15426 35924 15428
rect 35644 15374 35870 15426
rect 35922 15374 35924 15426
rect 35644 15372 35924 15374
rect 35868 15362 35924 15372
rect 35532 15316 35588 15326
rect 35532 15222 35588 15260
rect 37548 15148 37604 17054
rect 37772 17108 37828 22428
rect 37884 22260 37940 22270
rect 37884 19684 37940 22204
rect 37996 22036 38052 22428
rect 38220 22258 38276 22270
rect 38220 22206 38222 22258
rect 38274 22206 38276 22258
rect 37996 21980 38164 22036
rect 37996 21812 38052 21822
rect 37996 21718 38052 21756
rect 38108 21700 38164 21980
rect 38108 21634 38164 21644
rect 37884 19234 37940 19628
rect 37996 20802 38052 20814
rect 37996 20750 37998 20802
rect 38050 20750 38052 20802
rect 37996 19460 38052 20750
rect 38108 20578 38164 20590
rect 38108 20526 38110 20578
rect 38162 20526 38164 20578
rect 38108 20018 38164 20526
rect 38220 20132 38276 22206
rect 38444 21812 38500 23212
rect 38556 23042 38612 23660
rect 38556 22990 38558 23042
rect 38610 22990 38612 23042
rect 38556 22978 38612 22990
rect 38444 21746 38500 21756
rect 38668 22484 38724 22494
rect 38220 20066 38276 20076
rect 38108 19966 38110 20018
rect 38162 19966 38164 20018
rect 38108 19954 38164 19966
rect 38668 19796 38724 22428
rect 38892 22484 38948 25228
rect 39116 25218 39172 25228
rect 39340 24724 39396 27356
rect 39452 27188 39508 27580
rect 39564 27188 39620 27198
rect 39452 27186 39620 27188
rect 39452 27134 39566 27186
rect 39618 27134 39620 27186
rect 39452 27132 39620 27134
rect 39564 27122 39620 27132
rect 39676 27076 39732 27692
rect 40012 27746 40068 27804
rect 40012 27694 40014 27746
rect 40066 27694 40068 27746
rect 40012 27682 40068 27694
rect 40124 27858 40180 27870
rect 40124 27806 40126 27858
rect 40178 27806 40180 27858
rect 39676 27010 39732 27020
rect 40012 27188 40068 27198
rect 40012 27074 40068 27132
rect 40012 27022 40014 27074
rect 40066 27022 40068 27074
rect 40012 27010 40068 27022
rect 40124 26964 40180 27806
rect 40236 27076 40292 29148
rect 40796 29092 40852 30158
rect 40796 29026 40852 29036
rect 40684 28642 40740 28654
rect 40684 28590 40686 28642
rect 40738 28590 40740 28642
rect 40684 27748 40740 28590
rect 40684 27682 40740 27692
rect 40348 27076 40404 27086
rect 40236 27074 40404 27076
rect 40236 27022 40350 27074
rect 40402 27022 40404 27074
rect 40236 27020 40404 27022
rect 40348 27010 40404 27020
rect 40124 26898 40180 26908
rect 40684 26850 40740 26862
rect 40684 26798 40686 26850
rect 40738 26798 40740 26850
rect 40124 26628 40180 26638
rect 39676 26516 39732 26526
rect 39676 26422 39732 26460
rect 40124 25620 40180 26572
rect 40124 25526 40180 25564
rect 40460 25394 40516 25406
rect 40460 25342 40462 25394
rect 40514 25342 40516 25394
rect 39676 25282 39732 25294
rect 39676 25230 39678 25282
rect 39730 25230 39732 25282
rect 39676 24834 39732 25230
rect 39676 24782 39678 24834
rect 39730 24782 39732 24834
rect 39452 24724 39508 24734
rect 39340 24722 39508 24724
rect 39340 24670 39454 24722
rect 39506 24670 39508 24722
rect 39340 24668 39508 24670
rect 39452 24658 39508 24668
rect 39116 24612 39172 24622
rect 39116 24518 39172 24556
rect 39116 24276 39172 24286
rect 39116 23940 39172 24220
rect 39116 23874 39172 23884
rect 39004 23828 39060 23838
rect 39004 23154 39060 23772
rect 39004 23102 39006 23154
rect 39058 23102 39060 23154
rect 39004 23090 39060 23102
rect 38892 22418 38948 22428
rect 39116 20802 39172 20814
rect 39116 20750 39118 20802
rect 39170 20750 39172 20802
rect 38780 19908 38836 19918
rect 39116 19908 39172 20750
rect 39228 20692 39284 20702
rect 39228 20690 39396 20692
rect 39228 20638 39230 20690
rect 39282 20638 39396 20690
rect 39228 20636 39396 20638
rect 39228 20626 39284 20636
rect 39228 20020 39284 20030
rect 39228 19926 39284 19964
rect 38780 19906 39172 19908
rect 38780 19854 38782 19906
rect 38834 19854 39172 19906
rect 38780 19852 39172 19854
rect 38780 19842 38836 19852
rect 38668 19730 38724 19740
rect 37996 19404 38388 19460
rect 37884 19182 37886 19234
rect 37938 19182 37940 19234
rect 37884 19170 37940 19182
rect 38220 19236 38276 19246
rect 38220 19010 38276 19180
rect 38220 18958 38222 19010
rect 38274 18958 38276 19010
rect 37884 18676 37940 18686
rect 37884 17778 37940 18620
rect 38220 17780 38276 18958
rect 38332 18450 38388 19404
rect 38892 19236 38948 19246
rect 38892 19142 38948 19180
rect 38332 18398 38334 18450
rect 38386 18398 38388 18450
rect 38332 18340 38388 18398
rect 38332 18116 38388 18284
rect 38332 18050 38388 18060
rect 38444 19124 38500 19134
rect 37884 17726 37886 17778
rect 37938 17726 37940 17778
rect 37884 17714 37940 17726
rect 37996 17724 38276 17780
rect 37772 17042 37828 17052
rect 37660 15540 37716 15550
rect 37660 15446 37716 15484
rect 37436 15092 37604 15148
rect 37996 15092 38052 17724
rect 38444 17666 38500 19068
rect 38668 19012 38724 19022
rect 38668 19010 38836 19012
rect 38668 18958 38670 19010
rect 38722 18958 38836 19010
rect 38668 18956 38836 18958
rect 38668 18946 38724 18956
rect 38444 17614 38446 17666
rect 38498 17614 38500 17666
rect 38444 17602 38500 17614
rect 38556 18564 38612 18574
rect 38556 17444 38612 18508
rect 38780 18564 38836 18956
rect 38892 18564 38948 18574
rect 38780 18562 38948 18564
rect 38780 18510 38894 18562
rect 38946 18510 38948 18562
rect 38780 18508 38948 18510
rect 38780 18340 38836 18508
rect 38892 18498 38948 18508
rect 38780 18274 38836 18284
rect 39004 18452 39060 19852
rect 39340 19460 39396 20636
rect 39564 20018 39620 20030
rect 39564 19966 39566 20018
rect 39618 19966 39620 20018
rect 39564 19796 39620 19966
rect 39564 19730 39620 19740
rect 38332 17388 38612 17444
rect 38892 18228 38948 18238
rect 38892 17444 38948 18172
rect 39004 17556 39060 18396
rect 39116 19404 39396 19460
rect 39116 18228 39172 19404
rect 39340 19292 39620 19348
rect 39340 19234 39396 19292
rect 39340 19182 39342 19234
rect 39394 19182 39396 19234
rect 39340 19170 39396 19182
rect 39452 18452 39508 18462
rect 39452 18358 39508 18396
rect 39116 18162 39172 18172
rect 39228 18116 39284 18126
rect 39116 17556 39172 17566
rect 39004 17554 39172 17556
rect 39004 17502 39118 17554
rect 39170 17502 39172 17554
rect 39004 17500 39172 17502
rect 39116 17490 39172 17500
rect 38892 17388 39060 17444
rect 38220 17332 38276 17342
rect 38220 16098 38276 17276
rect 38220 16046 38222 16098
rect 38274 16046 38276 16098
rect 38220 16034 38276 16046
rect 38108 15428 38164 15438
rect 38108 15334 38164 15372
rect 38332 15148 38388 17388
rect 38556 17108 38612 17118
rect 38556 15986 38612 17052
rect 38556 15934 38558 15986
rect 38610 15934 38612 15986
rect 38556 15922 38612 15934
rect 38892 16996 38948 17006
rect 38892 15540 38948 16940
rect 38892 15474 38948 15484
rect 39004 16210 39060 17388
rect 39004 16158 39006 16210
rect 39058 16158 39060 16210
rect 38332 15092 38500 15148
rect 35196 15036 35588 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35532 14756 35588 15036
rect 34860 13692 35140 13748
rect 35196 14700 35588 14756
rect 34860 13188 34916 13692
rect 35196 13636 35252 14700
rect 35532 14532 35588 14542
rect 35532 14438 35588 14476
rect 36988 14418 37044 14430
rect 36988 14366 36990 14418
rect 37042 14366 37044 14418
rect 36988 14196 37044 14366
rect 37324 14308 37380 14318
rect 36988 14130 37044 14140
rect 37212 14306 37380 14308
rect 37212 14254 37326 14306
rect 37378 14254 37380 14306
rect 37212 14252 37380 14254
rect 35420 13860 35476 13870
rect 35420 13766 35476 13804
rect 35308 13748 35364 13758
rect 35308 13654 35364 13692
rect 34860 13122 34916 13132
rect 34972 13580 35252 13636
rect 36316 13634 36372 13646
rect 36316 13582 36318 13634
rect 36370 13582 36372 13634
rect 34636 12572 34804 12628
rect 34860 12962 34916 12974
rect 34860 12910 34862 12962
rect 34914 12910 34916 12962
rect 34636 11506 34692 12572
rect 34636 11454 34638 11506
rect 34690 11454 34692 11506
rect 34636 11442 34692 11454
rect 34860 12292 34916 12910
rect 34524 11342 34526 11394
rect 34578 11342 34580 11394
rect 34524 10612 34580 11342
rect 34524 10546 34580 10556
rect 34636 9828 34692 9838
rect 34860 9828 34916 12236
rect 34972 12178 35028 13580
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 13188 35252 13198
rect 35196 12404 35252 13132
rect 35420 12964 35476 12974
rect 35420 12962 35812 12964
rect 35420 12910 35422 12962
rect 35474 12910 35812 12962
rect 35420 12908 35812 12910
rect 35420 12898 35476 12908
rect 35196 12348 35700 12404
rect 35644 12290 35700 12348
rect 35756 12402 35812 12908
rect 36316 12962 36372 13582
rect 36316 12910 36318 12962
rect 36370 12910 36372 12962
rect 36316 12898 36372 12910
rect 35756 12350 35758 12402
rect 35810 12350 35812 12402
rect 35756 12338 35812 12350
rect 35644 12238 35646 12290
rect 35698 12238 35700 12290
rect 35644 12226 35700 12238
rect 36540 12290 36596 12302
rect 36540 12238 36542 12290
rect 36594 12238 36596 12290
rect 34972 12126 34974 12178
rect 35026 12126 35028 12178
rect 34972 11844 35028 12126
rect 35532 12180 35588 12190
rect 35532 12086 35588 12124
rect 36540 12180 36596 12238
rect 36540 12114 36596 12124
rect 36652 12292 36708 12302
rect 36652 12178 36708 12236
rect 36652 12126 36654 12178
rect 36706 12126 36708 12178
rect 36652 12114 36708 12126
rect 36988 12292 37044 12302
rect 34972 11778 35028 11788
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 36988 11282 37044 12236
rect 37212 12068 37268 14252
rect 37324 14242 37380 14252
rect 37324 13860 37380 13870
rect 37324 13074 37380 13804
rect 37324 13022 37326 13074
rect 37378 13022 37380 13074
rect 37324 13010 37380 13022
rect 37212 11394 37268 12012
rect 37212 11342 37214 11394
rect 37266 11342 37268 11394
rect 37212 11330 37268 11342
rect 36988 11230 36990 11282
rect 37042 11230 37044 11282
rect 36988 11218 37044 11230
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 34692 9772 34916 9828
rect 35084 9826 35140 9838
rect 35084 9774 35086 9826
rect 35138 9774 35140 9826
rect 34636 9734 34692 9772
rect 33964 9714 34132 9716
rect 33964 9662 33966 9714
rect 34018 9662 34132 9714
rect 33964 9660 34132 9662
rect 33964 9650 34020 9660
rect 34860 9042 34916 9054
rect 34860 8990 34862 9042
rect 34914 8990 34916 9042
rect 34076 8148 34132 8158
rect 34132 8092 34356 8148
rect 34076 8054 34132 8092
rect 33964 7476 34020 7486
rect 33964 7382 34020 7420
rect 34300 7474 34356 8092
rect 34300 7422 34302 7474
rect 34354 7422 34356 7474
rect 34300 7410 34356 7422
rect 34860 7364 34916 8990
rect 35084 8370 35140 9774
rect 35980 9826 36036 9838
rect 35980 9774 35982 9826
rect 36034 9774 36036 9826
rect 35420 9044 35476 9054
rect 35420 9042 35588 9044
rect 35420 8990 35422 9042
rect 35474 8990 35588 9042
rect 35420 8988 35588 8990
rect 35420 8978 35476 8988
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35084 8318 35086 8370
rect 35138 8318 35140 8370
rect 35084 8306 35140 8318
rect 35532 8372 35588 8988
rect 35532 8306 35588 8316
rect 35756 8260 35812 8270
rect 35756 8166 35812 8204
rect 35532 7700 35588 7710
rect 35980 7700 36036 9774
rect 37436 9268 37492 15092
rect 37996 15026 38052 15036
rect 37772 14418 37828 14430
rect 37772 14366 37774 14418
rect 37826 14366 37828 14418
rect 37772 14308 37828 14366
rect 37548 14252 37772 14308
rect 37548 12962 37604 14252
rect 37772 14242 37828 14252
rect 38108 14308 38164 14318
rect 38108 14306 38388 14308
rect 38108 14254 38110 14306
rect 38162 14254 38388 14306
rect 38108 14252 38388 14254
rect 38108 14242 38164 14252
rect 38220 14084 38276 14094
rect 37996 13860 38052 13870
rect 37996 13858 38164 13860
rect 37996 13806 37998 13858
rect 38050 13806 38164 13858
rect 37996 13804 38164 13806
rect 37996 13794 38052 13804
rect 37660 13748 37716 13758
rect 37660 13746 37828 13748
rect 37660 13694 37662 13746
rect 37714 13694 37828 13746
rect 37660 13692 37828 13694
rect 37660 13682 37716 13692
rect 37772 13300 37828 13692
rect 37548 12910 37550 12962
rect 37602 12910 37604 12962
rect 37548 12898 37604 12910
rect 37660 13244 38052 13300
rect 37660 12516 37716 13244
rect 37996 13074 38052 13244
rect 37996 13022 37998 13074
rect 38050 13022 38052 13074
rect 37996 13010 38052 13022
rect 37436 9202 37492 9212
rect 37548 12460 37716 12516
rect 37884 12964 37940 12974
rect 37548 9156 37604 12460
rect 37884 12404 37940 12908
rect 37660 12292 37716 12302
rect 37660 12198 37716 12236
rect 37772 11396 37828 11406
rect 37884 11396 37940 12348
rect 37772 11394 37940 11396
rect 37772 11342 37774 11394
rect 37826 11342 37940 11394
rect 37772 11340 37940 11342
rect 37996 12852 38052 12862
rect 37996 11394 38052 12796
rect 38108 12180 38164 13804
rect 38220 13746 38276 14028
rect 38220 13694 38222 13746
rect 38274 13694 38276 13746
rect 38220 12292 38276 13694
rect 38332 12964 38388 14252
rect 38444 14306 38500 15092
rect 38668 15092 38724 15102
rect 38668 14532 38724 15036
rect 38444 14254 38446 14306
rect 38498 14254 38500 14306
rect 38444 13748 38500 14254
rect 38444 13682 38500 13692
rect 38556 14530 38724 14532
rect 38556 14478 38670 14530
rect 38722 14478 38724 14530
rect 38556 14476 38724 14478
rect 38332 12898 38388 12908
rect 38556 12852 38612 14476
rect 38668 14466 38724 14476
rect 39004 14530 39060 16158
rect 39004 14478 39006 14530
rect 39058 14478 39060 14530
rect 39004 14466 39060 14478
rect 38780 13972 38836 13982
rect 38780 13878 38836 13916
rect 39228 13860 39284 18060
rect 39564 17220 39620 19292
rect 39676 18116 39732 24782
rect 40236 25284 40292 25294
rect 40236 24834 40292 25228
rect 40236 24782 40238 24834
rect 40290 24782 40292 24834
rect 40236 24770 40292 24782
rect 40012 24724 40068 24734
rect 40068 24668 40180 24724
rect 40012 24658 40068 24668
rect 39788 24388 39844 24398
rect 39788 23828 39844 24332
rect 39788 22482 39844 23772
rect 39788 22430 39790 22482
rect 39842 22430 39844 22482
rect 39788 22418 39844 22430
rect 40012 21812 40068 21822
rect 39900 20130 39956 20142
rect 39900 20078 39902 20130
rect 39954 20078 39956 20130
rect 39676 18050 39732 18060
rect 39788 20020 39844 20030
rect 39788 19234 39844 19964
rect 39788 19182 39790 19234
rect 39842 19182 39844 19234
rect 39452 16884 39508 16894
rect 39452 16790 39508 16828
rect 39564 16212 39620 17164
rect 39676 17892 39732 17902
rect 39676 16994 39732 17836
rect 39676 16942 39678 16994
rect 39730 16942 39732 16994
rect 39676 16930 39732 16942
rect 39788 16996 39844 19182
rect 39900 19908 39956 20078
rect 39900 19124 39956 19852
rect 39900 19058 39956 19068
rect 40012 18452 40068 21756
rect 40012 18386 40068 18396
rect 40012 17108 40068 17118
rect 40124 17108 40180 24668
rect 40236 23940 40292 23950
rect 40236 22370 40292 23884
rect 40460 23938 40516 25342
rect 40684 25396 40740 26798
rect 40684 25330 40740 25340
rect 40908 25620 40964 31892
rect 41580 31220 41636 31836
rect 41916 31220 41972 31230
rect 41580 31218 41972 31220
rect 41580 31166 41582 31218
rect 41634 31166 41918 31218
rect 41970 31166 41972 31218
rect 41580 31164 41972 31166
rect 41020 30884 41076 30894
rect 41020 30882 41188 30884
rect 41020 30830 41022 30882
rect 41074 30830 41188 30882
rect 41020 30828 41188 30830
rect 41020 30818 41076 30828
rect 41020 30210 41076 30222
rect 41020 30158 41022 30210
rect 41074 30158 41076 30210
rect 41020 30100 41076 30158
rect 41020 30034 41076 30044
rect 41020 29428 41076 29438
rect 41132 29428 41188 30828
rect 41468 30212 41524 30222
rect 41076 29372 41188 29428
rect 41356 29540 41412 29550
rect 41020 29334 41076 29372
rect 41020 27860 41076 27870
rect 41020 27766 41076 27804
rect 41244 27188 41300 27198
rect 41244 26908 41300 27132
rect 41356 27076 41412 29484
rect 41468 29426 41524 30156
rect 41468 29374 41470 29426
rect 41522 29374 41524 29426
rect 41468 28868 41524 29374
rect 41468 28802 41524 28812
rect 41356 26982 41412 27020
rect 40908 25506 40964 25564
rect 40908 25454 40910 25506
rect 40962 25454 40964 25506
rect 40908 25396 40964 25454
rect 40908 25330 40964 25340
rect 41132 26852 41300 26908
rect 41132 24724 41188 26852
rect 41580 26516 41636 31164
rect 41916 31154 41972 31164
rect 42028 30996 42084 33070
rect 42364 31948 42420 35532
rect 42700 34914 42756 34926
rect 42700 34862 42702 34914
rect 42754 34862 42756 34914
rect 42700 34468 42756 34862
rect 42700 34402 42756 34412
rect 42700 33348 42756 33358
rect 42812 33348 42868 36990
rect 43036 36596 43092 36606
rect 43036 36484 43092 36540
rect 43036 36482 43204 36484
rect 43036 36430 43038 36482
rect 43090 36430 43204 36482
rect 43036 36428 43204 36430
rect 43036 36418 43092 36428
rect 43036 35924 43092 35934
rect 43036 35830 43092 35868
rect 42756 33292 42868 33348
rect 42700 33254 42756 33292
rect 42028 30930 42084 30940
rect 42140 31892 42420 31948
rect 42700 32562 42756 32574
rect 42700 32510 42702 32562
rect 42754 32510 42756 32562
rect 41692 30884 41748 30894
rect 41748 30828 41860 30884
rect 41692 30818 41748 30828
rect 41692 30210 41748 30222
rect 41692 30158 41694 30210
rect 41746 30158 41748 30210
rect 41692 28980 41748 30158
rect 41804 29540 41860 30828
rect 42140 30212 42196 31892
rect 42700 31780 42756 32510
rect 43148 32562 43204 36428
rect 43260 36482 43316 37884
rect 43708 37874 43764 37884
rect 44156 37268 44212 37278
rect 44156 37174 44212 37212
rect 43820 37156 43876 37166
rect 43372 37044 43428 37054
rect 43372 36594 43428 36988
rect 43372 36542 43374 36594
rect 43426 36542 43428 36594
rect 43372 36530 43428 36542
rect 43260 36430 43262 36482
rect 43314 36430 43316 36482
rect 43260 35700 43316 36430
rect 43484 36484 43540 36494
rect 43484 36390 43540 36428
rect 43484 35700 43540 35710
rect 43260 35698 43540 35700
rect 43260 35646 43486 35698
rect 43538 35646 43540 35698
rect 43260 35644 43540 35646
rect 43260 35476 43316 35644
rect 43484 35634 43540 35644
rect 43260 35410 43316 35420
rect 43148 32510 43150 32562
rect 43202 32510 43204 32562
rect 43148 32498 43204 32510
rect 43260 33346 43316 33358
rect 43260 33294 43262 33346
rect 43314 33294 43316 33346
rect 43260 32340 43316 33294
rect 43260 32274 43316 32284
rect 42700 31714 42756 31724
rect 42252 31108 42308 31118
rect 42252 31106 42532 31108
rect 42252 31054 42254 31106
rect 42306 31054 42532 31106
rect 42252 31052 42532 31054
rect 42252 31042 42308 31052
rect 42140 30146 42196 30156
rect 42364 29988 42420 29998
rect 41804 29474 41860 29484
rect 41916 29986 42420 29988
rect 41916 29934 42366 29986
rect 42418 29934 42420 29986
rect 41916 29932 42420 29934
rect 41916 29538 41972 29932
rect 42364 29922 42420 29932
rect 41916 29486 41918 29538
rect 41970 29486 41972 29538
rect 41916 29474 41972 29486
rect 42252 29428 42308 29438
rect 41692 28914 41748 28924
rect 42028 29426 42308 29428
rect 42028 29374 42254 29426
rect 42306 29374 42308 29426
rect 42028 29372 42308 29374
rect 42028 28756 42084 29372
rect 42252 29362 42308 29372
rect 41692 28700 42084 28756
rect 41692 27188 41748 28700
rect 42476 28644 42532 31052
rect 43596 31106 43652 31118
rect 43596 31054 43598 31106
rect 43650 31054 43652 31106
rect 43260 30882 43316 30894
rect 43260 30830 43262 30882
rect 43314 30830 43316 30882
rect 43260 30324 43316 30830
rect 42812 30098 42868 30110
rect 42812 30046 42814 30098
rect 42866 30046 42868 30098
rect 42812 29652 42868 30046
rect 42812 29586 42868 29596
rect 42924 29538 42980 29550
rect 42924 29486 42926 29538
rect 42978 29486 42980 29538
rect 42700 29426 42756 29438
rect 42700 29374 42702 29426
rect 42754 29374 42756 29426
rect 42700 28754 42756 29374
rect 42700 28702 42702 28754
rect 42754 28702 42756 28754
rect 42700 28690 42756 28702
rect 42812 29092 42868 29102
rect 41916 28642 42532 28644
rect 41916 28590 42478 28642
rect 42530 28590 42532 28642
rect 41916 28588 42532 28590
rect 41692 27122 41748 27132
rect 41804 28418 41860 28430
rect 41804 28366 41806 28418
rect 41858 28366 41860 28418
rect 41804 27074 41860 28366
rect 41916 27858 41972 28588
rect 42476 28578 42532 28588
rect 42812 28420 42868 29036
rect 42924 28644 42980 29486
rect 42924 28578 42980 28588
rect 43036 29428 43092 29438
rect 42812 28364 42980 28420
rect 41916 27806 41918 27858
rect 41970 27806 41972 27858
rect 41916 27794 41972 27806
rect 42924 27858 42980 28364
rect 42924 27806 42926 27858
rect 42978 27806 42980 27858
rect 42924 27794 42980 27806
rect 42812 27746 42868 27758
rect 42812 27694 42814 27746
rect 42866 27694 42868 27746
rect 41804 27022 41806 27074
rect 41858 27022 41860 27074
rect 41804 27010 41860 27022
rect 42588 27076 42644 27086
rect 41580 26450 41636 26460
rect 41356 25506 41412 25518
rect 42476 25508 42532 25518
rect 41356 25454 41358 25506
rect 41410 25454 41412 25506
rect 41244 24724 41300 24734
rect 41132 24722 41300 24724
rect 41132 24670 41246 24722
rect 41298 24670 41300 24722
rect 41132 24668 41300 24670
rect 41244 24658 41300 24668
rect 40908 24610 40964 24622
rect 40908 24558 40910 24610
rect 40962 24558 40964 24610
rect 40908 24164 40964 24558
rect 40908 24098 40964 24108
rect 40460 23886 40462 23938
rect 40514 23886 40516 23938
rect 40460 23874 40516 23886
rect 41132 23940 41188 23950
rect 41132 23846 41188 23884
rect 40796 23828 40852 23838
rect 40796 23734 40852 23772
rect 41356 22482 41412 25454
rect 42028 25506 42532 25508
rect 42028 25454 42478 25506
rect 42530 25454 42532 25506
rect 42028 25452 42532 25454
rect 41692 25396 41748 25406
rect 41468 25284 41524 25294
rect 41468 25190 41524 25228
rect 41356 22430 41358 22482
rect 41410 22430 41412 22482
rect 41356 22418 41412 22430
rect 41580 23714 41636 23726
rect 41580 23662 41582 23714
rect 41634 23662 41636 23714
rect 40236 22318 40238 22370
rect 40290 22318 40292 22370
rect 40236 20020 40292 22318
rect 40236 19236 40292 19964
rect 40572 22148 40628 22158
rect 41580 22148 41636 23662
rect 40572 22146 41636 22148
rect 40572 22094 40574 22146
rect 40626 22094 41636 22146
rect 40572 22092 41636 22094
rect 40348 19906 40404 19918
rect 40348 19854 40350 19906
rect 40402 19854 40404 19906
rect 40348 19684 40404 19854
rect 40572 19908 40628 22092
rect 41132 21700 41188 21710
rect 41132 21606 41188 21644
rect 41468 21700 41524 21710
rect 41468 21606 41524 21644
rect 41692 21476 41748 25340
rect 41916 25394 41972 25406
rect 41916 25342 41918 25394
rect 41970 25342 41972 25394
rect 41916 25284 41972 25342
rect 41916 25218 41972 25228
rect 41916 24834 41972 24846
rect 41916 24782 41918 24834
rect 41970 24782 41972 24834
rect 41804 24722 41860 24734
rect 41804 24670 41806 24722
rect 41858 24670 41860 24722
rect 41804 24052 41860 24670
rect 41916 24276 41972 24782
rect 41916 24210 41972 24220
rect 41916 24052 41972 24062
rect 41804 24050 41972 24052
rect 41804 23998 41918 24050
rect 41970 23998 41972 24050
rect 41804 23996 41972 23998
rect 41916 23986 41972 23996
rect 42028 23378 42084 25452
rect 42476 25442 42532 25452
rect 42028 23326 42030 23378
rect 42082 23326 42084 23378
rect 42028 23314 42084 23326
rect 42140 25284 42196 25294
rect 42140 22820 42196 25228
rect 42588 24722 42644 27020
rect 42812 27074 42868 27694
rect 42812 27022 42814 27074
rect 42866 27022 42868 27074
rect 42812 27010 42868 27022
rect 43036 26908 43092 29372
rect 43148 28644 43204 28654
rect 43260 28644 43316 30268
rect 43484 30436 43540 30446
rect 43148 28642 43316 28644
rect 43148 28590 43150 28642
rect 43202 28590 43316 28642
rect 43148 28588 43316 28590
rect 43372 29652 43428 29662
rect 43372 28644 43428 29596
rect 43484 28868 43540 30380
rect 43596 30212 43652 31054
rect 43596 30146 43652 30156
rect 43596 29540 43652 29550
rect 43596 29426 43652 29484
rect 43596 29374 43598 29426
rect 43650 29374 43652 29426
rect 43596 29362 43652 29374
rect 43596 28868 43652 28878
rect 43484 28866 43652 28868
rect 43484 28814 43598 28866
rect 43650 28814 43652 28866
rect 43484 28812 43652 28814
rect 43596 28802 43652 28812
rect 43708 28756 43764 28766
rect 43708 28644 43764 28700
rect 43372 28588 43764 28644
rect 43148 28578 43204 28588
rect 43820 28532 43876 37100
rect 44828 36372 44884 36382
rect 44828 35810 44884 36316
rect 44828 35758 44830 35810
rect 44882 35758 44884 35810
rect 44828 35746 44884 35758
rect 44940 35924 44996 35934
rect 44716 35586 44772 35598
rect 44716 35534 44718 35586
rect 44770 35534 44772 35586
rect 44716 35028 44772 35534
rect 43932 34972 44772 35028
rect 43932 34802 43988 34972
rect 43932 34750 43934 34802
rect 43986 34750 43988 34802
rect 43932 32340 43988 34750
rect 44044 34804 44100 34814
rect 44044 34020 44100 34748
rect 44044 32562 44100 33964
rect 44828 34690 44884 34702
rect 44828 34638 44830 34690
rect 44882 34638 44884 34690
rect 44828 34020 44884 34638
rect 44940 34242 44996 35868
rect 45164 34804 45220 34814
rect 45164 34710 45220 34748
rect 44940 34190 44942 34242
rect 44994 34190 44996 34242
rect 44940 34178 44996 34190
rect 45388 34132 45444 34142
rect 45388 34038 45444 34076
rect 44828 33954 44884 33964
rect 44156 33908 44212 33918
rect 44156 33346 44212 33852
rect 45948 33908 46004 33918
rect 45948 33814 46004 33852
rect 44156 33294 44158 33346
rect 44210 33294 44212 33346
rect 44156 33282 44212 33294
rect 44044 32510 44046 32562
rect 44098 32510 44100 32562
rect 44044 32498 44100 32510
rect 45836 33124 45892 33134
rect 43932 32274 43988 32284
rect 45164 32340 45220 32350
rect 45164 32246 45220 32284
rect 45612 31892 45668 31902
rect 44940 31554 44996 31566
rect 44940 31502 44942 31554
rect 44994 31502 44996 31554
rect 44940 31444 44996 31502
rect 44828 31388 44940 31444
rect 44828 30772 44884 31388
rect 44940 31378 44996 31388
rect 45052 30996 45108 31006
rect 45052 30994 45556 30996
rect 45052 30942 45054 30994
rect 45106 30942 45556 30994
rect 45052 30940 45556 30942
rect 45052 30930 45108 30940
rect 44828 30706 44884 30716
rect 44940 30884 44996 30894
rect 44828 30324 44884 30334
rect 44268 30212 44324 30222
rect 43708 28476 43876 28532
rect 43932 29426 43988 29438
rect 43932 29374 43934 29426
rect 43986 29374 43988 29426
rect 43932 28532 43988 29374
rect 44268 29316 44324 30156
rect 44828 30098 44884 30268
rect 44828 30046 44830 30098
rect 44882 30046 44884 30098
rect 44828 30034 44884 30046
rect 44940 29426 44996 30828
rect 45164 30772 45220 30782
rect 45164 30210 45220 30716
rect 45164 30158 45166 30210
rect 45218 30158 45220 30210
rect 45164 30146 45220 30158
rect 45500 30436 45556 30940
rect 44940 29374 44942 29426
rect 44994 29374 44996 29426
rect 44940 29362 44996 29374
rect 45388 30100 45444 30110
rect 44492 29316 44548 29326
rect 44268 29260 44492 29316
rect 43708 27412 43764 28476
rect 43932 28466 43988 28476
rect 44156 28530 44212 28542
rect 44156 28478 44158 28530
rect 44210 28478 44212 28530
rect 44156 28420 44212 28478
rect 44492 28420 44548 29260
rect 45388 28866 45444 30044
rect 45500 30098 45556 30380
rect 45500 30046 45502 30098
rect 45554 30046 45556 30098
rect 45500 30034 45556 30046
rect 45500 29652 45556 29662
rect 45612 29652 45668 31836
rect 45724 30884 45780 30894
rect 45724 30790 45780 30828
rect 45836 30210 45892 33068
rect 45836 30158 45838 30210
rect 45890 30158 45892 30210
rect 45836 30146 45892 30158
rect 45500 29650 45668 29652
rect 45500 29598 45502 29650
rect 45554 29598 45668 29650
rect 45500 29596 45668 29598
rect 45500 29586 45556 29596
rect 45948 29316 46004 29326
rect 45948 29222 46004 29260
rect 45388 28814 45390 28866
rect 45442 28814 45444 28866
rect 45388 28802 45444 28814
rect 45612 28980 45668 28990
rect 44156 28364 44548 28420
rect 43708 27346 43764 27356
rect 43820 28308 43876 28318
rect 43036 26852 43204 26908
rect 42588 24670 42590 24722
rect 42642 24670 42644 24722
rect 42588 24658 42644 24670
rect 42924 24722 42980 24734
rect 42924 24670 42926 24722
rect 42978 24670 42980 24722
rect 42028 22764 42196 22820
rect 42364 24108 42644 24164
rect 41916 21476 41972 21486
rect 41692 21474 41972 21476
rect 41692 21422 41918 21474
rect 41970 21422 41972 21474
rect 41692 21420 41972 21422
rect 41132 20916 41188 20926
rect 41132 20914 41860 20916
rect 41132 20862 41134 20914
rect 41186 20862 41860 20914
rect 41132 20860 41860 20862
rect 41132 20850 41188 20860
rect 41804 20130 41860 20860
rect 41804 20078 41806 20130
rect 41858 20078 41860 20130
rect 41804 20066 41860 20078
rect 40572 19842 40628 19852
rect 41020 20018 41076 20030
rect 41020 19966 41022 20018
rect 41074 19966 41076 20018
rect 40348 19618 40404 19628
rect 40908 19684 40964 19694
rect 41020 19684 41076 19966
rect 41356 20020 41412 20030
rect 41916 20020 41972 21420
rect 42028 20244 42084 22764
rect 42140 22372 42196 22382
rect 42364 22372 42420 24108
rect 42140 22370 42420 22372
rect 42140 22318 42142 22370
rect 42194 22318 42420 22370
rect 42140 22316 42420 22318
rect 42140 22306 42196 22316
rect 42140 20692 42196 20702
rect 42140 20598 42196 20636
rect 42028 20178 42084 20188
rect 42140 20020 42196 20030
rect 41916 20018 42196 20020
rect 41916 19966 42142 20018
rect 42194 19966 42196 20018
rect 41916 19964 42196 19966
rect 41356 19908 41412 19964
rect 41356 19906 41636 19908
rect 41356 19854 41358 19906
rect 41410 19854 41636 19906
rect 41356 19852 41636 19854
rect 41356 19842 41412 19852
rect 40964 19628 41076 19684
rect 40908 19618 40964 19628
rect 40236 19170 40292 19180
rect 40460 19460 40516 19470
rect 40012 17106 40292 17108
rect 40012 17054 40014 17106
rect 40066 17054 40292 17106
rect 40012 17052 40292 17054
rect 40012 17042 40068 17052
rect 39900 16996 39956 17006
rect 39788 16940 39900 16996
rect 39900 16930 39956 16940
rect 39564 16156 40068 16212
rect 39452 16100 39508 16110
rect 39564 16100 39620 16156
rect 39452 16098 39620 16100
rect 39452 16046 39454 16098
rect 39506 16046 39620 16098
rect 39452 16044 39620 16046
rect 39452 16034 39508 16044
rect 39788 15986 39844 15998
rect 39788 15934 39790 15986
rect 39842 15934 39844 15986
rect 39340 15428 39396 15438
rect 39340 14532 39396 15372
rect 39676 15428 39732 15438
rect 39788 15428 39844 15934
rect 40012 15538 40068 16156
rect 40012 15486 40014 15538
rect 40066 15486 40068 15538
rect 40012 15474 40068 15486
rect 40124 16098 40180 16110
rect 40124 16046 40126 16098
rect 40178 16046 40180 16098
rect 40124 15988 40180 16046
rect 39676 15426 39844 15428
rect 39676 15374 39678 15426
rect 39730 15374 39844 15426
rect 39676 15372 39844 15374
rect 39676 15362 39732 15372
rect 39340 14438 39396 14476
rect 39340 13860 39396 13870
rect 39284 13858 39396 13860
rect 39284 13806 39342 13858
rect 39394 13806 39396 13858
rect 39284 13804 39396 13806
rect 39228 13766 39284 13804
rect 39340 13794 39396 13804
rect 39900 13858 39956 13870
rect 39900 13806 39902 13858
rect 39954 13806 39956 13858
rect 39116 13524 39172 13534
rect 39116 13522 39508 13524
rect 39116 13470 39118 13522
rect 39170 13470 39508 13522
rect 39116 13468 39508 13470
rect 39116 13458 39172 13468
rect 38780 12964 38836 12974
rect 38556 12786 38612 12796
rect 38668 12850 38724 12862
rect 38668 12798 38670 12850
rect 38722 12798 38724 12850
rect 38668 12292 38724 12798
rect 38220 12236 38388 12292
rect 38108 12114 38164 12124
rect 37996 11342 37998 11394
rect 38050 11342 38052 11394
rect 37772 11330 37828 11340
rect 37996 11330 38052 11342
rect 38332 11394 38388 12236
rect 38332 11342 38334 11394
rect 38386 11342 38388 11394
rect 38332 11330 38388 11342
rect 38444 12180 38500 12190
rect 38444 11172 38500 12124
rect 38332 11116 38500 11172
rect 38556 12068 38612 12078
rect 37548 9062 37604 9100
rect 37884 9156 37940 9166
rect 37884 8258 37940 9100
rect 37884 8206 37886 8258
rect 37938 8206 37940 8258
rect 37884 8194 37940 8206
rect 38332 8260 38388 11116
rect 38444 9714 38500 9726
rect 38444 9662 38446 9714
rect 38498 9662 38500 9714
rect 38444 9268 38500 9662
rect 38556 9492 38612 12012
rect 38668 11394 38724 12236
rect 38668 11342 38670 11394
rect 38722 11342 38724 11394
rect 38668 11330 38724 11342
rect 38780 9826 38836 12908
rect 38780 9774 38782 9826
rect 38834 9774 38836 9826
rect 38780 9762 38836 9774
rect 39340 9826 39396 9838
rect 39340 9774 39342 9826
rect 39394 9774 39396 9826
rect 38556 9426 38612 9436
rect 38556 9268 38612 9278
rect 38444 9266 38612 9268
rect 38444 9214 38558 9266
rect 38610 9214 38612 9266
rect 38444 9212 38612 9214
rect 38556 9202 38612 9212
rect 38556 8932 38612 8942
rect 38444 8260 38500 8270
rect 38332 8258 38500 8260
rect 38332 8206 38446 8258
rect 38498 8206 38500 8258
rect 38332 8204 38500 8206
rect 38444 8194 38500 8204
rect 35532 7698 36036 7700
rect 35532 7646 35534 7698
rect 35586 7646 36036 7698
rect 35532 7644 36036 7646
rect 36092 8034 36148 8046
rect 36092 7982 36094 8034
rect 36146 7982 36148 8034
rect 35532 7634 35588 7644
rect 34860 7298 34916 7308
rect 35644 7474 35700 7486
rect 35644 7422 35646 7474
rect 35698 7422 35700 7474
rect 35644 7364 35700 7422
rect 36092 7476 36148 7982
rect 38556 7698 38612 8876
rect 38556 7646 38558 7698
rect 38610 7646 38612 7698
rect 38556 7634 38612 7646
rect 36204 7476 36260 7486
rect 36092 7420 36204 7476
rect 36204 7382 36260 7420
rect 35644 7298 35700 7308
rect 39340 7250 39396 9774
rect 39452 9714 39508 13468
rect 39900 13300 39956 13806
rect 39900 13234 39956 13244
rect 40124 12964 40180 15932
rect 40236 15314 40292 17052
rect 40236 15262 40238 15314
rect 40290 15262 40292 15314
rect 40236 15250 40292 15262
rect 40460 15148 40516 19404
rect 41580 18674 41636 19852
rect 42140 19348 42196 19964
rect 42140 19282 42196 19292
rect 41580 18622 41582 18674
rect 41634 18622 41636 18674
rect 41580 18610 41636 18622
rect 41356 18564 41412 18574
rect 41356 18470 41412 18508
rect 42028 18450 42084 18462
rect 42028 18398 42030 18450
rect 42082 18398 42084 18450
rect 42028 17220 42084 18398
rect 42028 17154 42084 17164
rect 42252 17780 42308 17790
rect 42364 17780 42420 22316
rect 42476 23940 42532 23950
rect 42476 22370 42532 23884
rect 42588 23938 42644 24108
rect 42588 23886 42590 23938
rect 42642 23886 42644 23938
rect 42588 23874 42644 23886
rect 42476 22318 42478 22370
rect 42530 22318 42532 22370
rect 42476 21586 42532 22318
rect 42476 21534 42478 21586
rect 42530 21534 42532 21586
rect 42476 21522 42532 21534
rect 42588 23154 42644 23166
rect 42588 23102 42590 23154
rect 42642 23102 42644 23154
rect 42588 22372 42644 23102
rect 42924 23156 42980 24670
rect 43036 23940 43092 23950
rect 43036 23846 43092 23884
rect 43036 23156 43092 23166
rect 42924 23100 43036 23156
rect 43036 23090 43092 23100
rect 42476 20692 42532 20702
rect 42588 20692 42644 22316
rect 42700 21700 42756 21710
rect 42700 20802 42756 21644
rect 42700 20750 42702 20802
rect 42754 20750 42756 20802
rect 42700 20738 42756 20750
rect 42532 20636 42644 20692
rect 42476 20578 42532 20636
rect 42476 20526 42478 20578
rect 42530 20526 42532 20578
rect 42476 18450 42532 20526
rect 42812 20132 42868 20142
rect 42812 20038 42868 20076
rect 42700 20018 42756 20030
rect 42700 19966 42702 20018
rect 42754 19966 42756 20018
rect 42588 19124 42644 19134
rect 42588 19030 42644 19068
rect 42476 18398 42478 18450
rect 42530 18398 42532 18450
rect 42476 18386 42532 18398
rect 42588 17892 42644 17902
rect 42700 17892 42756 19966
rect 42588 17890 42756 17892
rect 42588 17838 42590 17890
rect 42642 17838 42756 17890
rect 42588 17836 42756 17838
rect 42588 17826 42644 17836
rect 42308 17724 42420 17780
rect 41244 16884 41300 16894
rect 40348 15092 40516 15148
rect 40684 16098 40740 16110
rect 40684 16046 40686 16098
rect 40738 16046 40740 16098
rect 40684 15148 40740 16046
rect 41244 16098 41300 16828
rect 41244 16046 41246 16098
rect 41298 16046 41300 16098
rect 40796 15876 40852 15886
rect 40796 15782 40852 15820
rect 40684 15092 40964 15148
rect 40348 13972 40404 15092
rect 40348 13906 40404 13916
rect 40908 13970 40964 15092
rect 40908 13918 40910 13970
rect 40962 13918 40964 13970
rect 40908 13906 40964 13918
rect 41132 14532 41188 14542
rect 41132 13746 41188 14476
rect 41132 13694 41134 13746
rect 41186 13694 41188 13746
rect 41132 13682 41188 13694
rect 40908 13300 40964 13310
rect 40236 12964 40292 12974
rect 40684 12964 40740 12974
rect 40180 12962 40292 12964
rect 40180 12910 40238 12962
rect 40290 12910 40292 12962
rect 40180 12908 40292 12910
rect 40124 12870 40180 12908
rect 40236 12898 40292 12908
rect 40348 12962 40740 12964
rect 40348 12910 40686 12962
rect 40738 12910 40740 12962
rect 40348 12908 40740 12910
rect 39676 12852 39732 12862
rect 39900 12852 39956 12862
rect 39676 12850 39956 12852
rect 39676 12798 39678 12850
rect 39730 12798 39902 12850
rect 39954 12798 39956 12850
rect 39676 12796 39956 12798
rect 39676 12786 39732 12796
rect 39900 12786 39956 12796
rect 40236 12404 40292 12414
rect 40348 12404 40404 12908
rect 40684 12898 40740 12908
rect 40908 12850 40964 13244
rect 40908 12798 40910 12850
rect 40962 12798 40964 12850
rect 40908 12786 40964 12798
rect 41244 12852 41300 16046
rect 41916 16100 41972 16110
rect 41916 16006 41972 16044
rect 41356 15314 41412 15326
rect 41356 15262 41358 15314
rect 41410 15262 41412 15314
rect 41356 15092 41412 15262
rect 42252 15314 42308 17724
rect 42252 15262 42254 15314
rect 42306 15262 42308 15314
rect 42252 15250 42308 15262
rect 42364 16884 42420 16894
rect 41356 15026 41412 15036
rect 42364 14308 42420 16828
rect 42924 16098 42980 16110
rect 42924 16046 42926 16098
rect 42978 16046 42980 16098
rect 42924 15148 42980 16046
rect 42924 15092 43092 15148
rect 43036 14754 43092 15092
rect 43036 14702 43038 14754
rect 43090 14702 43092 14754
rect 43036 14690 43092 14702
rect 43148 14308 43204 26852
rect 43820 26514 43876 28252
rect 43820 26462 43822 26514
rect 43874 26462 43876 26514
rect 43820 26450 43876 26462
rect 44044 28308 44100 28318
rect 44044 27858 44100 28252
rect 44044 27806 44046 27858
rect 44098 27806 44100 27858
rect 43484 25508 43540 25518
rect 43372 25506 43540 25508
rect 43372 25454 43486 25506
rect 43538 25454 43540 25506
rect 43372 25452 43540 25454
rect 43372 21362 43428 25452
rect 43484 25442 43540 25452
rect 44044 24948 44100 27806
rect 44492 27746 44548 28364
rect 44492 27694 44494 27746
rect 44546 27694 44548 27746
rect 44492 27682 44548 27694
rect 44604 28756 44660 28766
rect 44604 27188 44660 28700
rect 45612 28642 45668 28924
rect 45612 28590 45614 28642
rect 45666 28590 45668 28642
rect 44828 28530 44884 28542
rect 44828 28478 44830 28530
rect 44882 28478 44884 28530
rect 44828 28308 44884 28478
rect 44940 28532 44996 28542
rect 44940 28438 44996 28476
rect 45052 28530 45108 28542
rect 45052 28478 45054 28530
rect 45106 28478 45108 28530
rect 44828 28242 44884 28252
rect 44604 27132 44884 27188
rect 44156 26964 44212 26974
rect 44156 26514 44212 26908
rect 44156 26462 44158 26514
rect 44210 26462 44212 26514
rect 44156 26450 44212 26462
rect 44716 26964 44772 26974
rect 44044 24892 44324 24948
rect 44268 24836 44324 24892
rect 44492 24836 44548 24846
rect 44268 24780 44492 24836
rect 44492 24742 44548 24780
rect 44044 24722 44100 24734
rect 44716 24724 44772 26908
rect 44828 25506 44884 27132
rect 45052 26964 45108 28478
rect 45052 26898 45108 26908
rect 45612 26908 45668 28590
rect 45612 26852 45780 26908
rect 44828 25454 44830 25506
rect 44882 25454 44884 25506
rect 44828 25442 44884 25454
rect 45276 25618 45332 25630
rect 45276 25566 45278 25618
rect 45330 25566 45332 25618
rect 45052 24836 45108 24846
rect 45276 24836 45332 25566
rect 45108 24780 45332 24836
rect 45052 24770 45108 24780
rect 44044 24670 44046 24722
rect 44098 24670 44100 24722
rect 44044 24612 44100 24670
rect 44044 24546 44100 24556
rect 44604 24722 44772 24724
rect 44604 24670 44718 24722
rect 44770 24670 44772 24722
rect 44604 24668 44772 24670
rect 44604 24388 44660 24668
rect 44716 24658 44772 24668
rect 44940 24724 44996 24734
rect 44828 24612 44884 24622
rect 44828 24498 44884 24556
rect 44828 24446 44830 24498
rect 44882 24446 44884 24498
rect 44828 24434 44884 24446
rect 44156 24332 44660 24388
rect 44156 23938 44212 24332
rect 44940 24276 44996 24668
rect 44156 23886 44158 23938
rect 44210 23886 44212 23938
rect 44156 23874 44212 23886
rect 44828 24220 44996 24276
rect 45500 24722 45556 24734
rect 45500 24670 45502 24722
rect 45554 24670 45556 24722
rect 44828 23938 44884 24220
rect 45276 24050 45332 24062
rect 45276 23998 45278 24050
rect 45330 23998 45332 24050
rect 44828 23886 44830 23938
rect 44882 23886 44884 23938
rect 44828 23874 44884 23886
rect 44940 23940 44996 23950
rect 45276 23940 45332 23998
rect 44996 23884 45332 23940
rect 44492 23828 44548 23838
rect 44492 23266 44548 23772
rect 44492 23214 44494 23266
rect 44546 23214 44548 23266
rect 44492 23202 44548 23214
rect 44716 23604 44772 23614
rect 43484 22372 43540 22382
rect 43484 22278 43540 22316
rect 43596 21700 43652 21710
rect 43596 21586 43652 21644
rect 43596 21534 43598 21586
rect 43650 21534 43652 21586
rect 43596 21522 43652 21534
rect 44716 21586 44772 23548
rect 44940 23154 44996 23884
rect 45500 23380 45556 24670
rect 45724 24722 45780 26852
rect 45724 24670 45726 24722
rect 45778 24670 45780 24722
rect 45724 24658 45780 24670
rect 45948 24500 46004 24510
rect 45948 23938 46004 24444
rect 45948 23886 45950 23938
rect 46002 23886 46004 23938
rect 45948 23874 46004 23886
rect 45724 23714 45780 23726
rect 45724 23662 45726 23714
rect 45778 23662 45780 23714
rect 45724 23380 45780 23662
rect 44940 23102 44942 23154
rect 44994 23102 44996 23154
rect 44940 23090 44996 23102
rect 45276 23324 45780 23380
rect 45164 21700 45220 21710
rect 45276 21700 45332 23324
rect 45500 23156 45556 23166
rect 45500 23062 45556 23100
rect 45164 21698 45332 21700
rect 45164 21646 45166 21698
rect 45218 21646 45332 21698
rect 45164 21644 45332 21646
rect 45164 21634 45220 21644
rect 44716 21534 44718 21586
rect 44770 21534 44772 21586
rect 44716 21522 44772 21534
rect 43372 21310 43374 21362
rect 43426 21310 43428 21362
rect 43372 21298 43428 21310
rect 43260 20132 43316 20142
rect 43260 20038 43316 20076
rect 44044 20018 44100 20030
rect 44044 19966 44046 20018
rect 44098 19966 44100 20018
rect 44044 19458 44100 19966
rect 44044 19406 44046 19458
rect 44098 19406 44100 19458
rect 44044 19394 44100 19406
rect 44940 20018 44996 20030
rect 44940 19966 44942 20018
rect 44994 19966 44996 20018
rect 43596 18452 43652 18462
rect 43484 16996 43540 17006
rect 43372 16884 43428 16894
rect 43372 15986 43428 16828
rect 43484 16882 43540 16940
rect 43484 16830 43486 16882
rect 43538 16830 43540 16882
rect 43484 16818 43540 16830
rect 43596 16098 43652 18396
rect 44940 18452 44996 19966
rect 44940 18386 44996 18396
rect 45052 18562 45108 18574
rect 45052 18510 45054 18562
rect 45106 18510 45108 18562
rect 44380 17220 44436 17230
rect 44380 16882 44436 17164
rect 44380 16830 44382 16882
rect 44434 16830 44436 16882
rect 44380 16818 44436 16830
rect 45052 16884 45108 18510
rect 45948 18452 46004 18462
rect 45948 18358 46004 18396
rect 45052 16818 45108 16828
rect 45500 16772 45556 16782
rect 43596 16046 43598 16098
rect 43650 16046 43652 16098
rect 43596 16034 43652 16046
rect 45276 16770 45556 16772
rect 45276 16718 45502 16770
rect 45554 16718 45556 16770
rect 45276 16716 45556 16718
rect 45276 16100 45332 16716
rect 45500 16706 45556 16716
rect 43372 15934 43374 15986
rect 43426 15934 43428 15986
rect 43372 15922 43428 15934
rect 42364 14306 42756 14308
rect 42364 14254 42366 14306
rect 42418 14254 42756 14306
rect 42364 14252 42756 14254
rect 42364 14242 42420 14252
rect 42700 13746 42756 14252
rect 43148 14242 43204 14252
rect 45276 15092 45332 16044
rect 45388 15092 45444 15102
rect 45276 15090 45444 15092
rect 45276 15038 45390 15090
rect 45442 15038 45444 15090
rect 45276 15036 45444 15038
rect 45276 13858 45332 15036
rect 45388 15026 45444 15036
rect 45276 13806 45278 13858
rect 45330 13806 45332 13858
rect 45276 13794 45332 13806
rect 42700 13694 42702 13746
rect 42754 13694 42756 13746
rect 42700 13682 42756 13694
rect 43708 13748 43764 13758
rect 43708 13654 43764 13692
rect 42140 12962 42196 12974
rect 42140 12910 42142 12962
rect 42194 12910 42196 12962
rect 41356 12852 41412 12862
rect 41244 12850 41412 12852
rect 41244 12798 41358 12850
rect 41410 12798 41412 12850
rect 41244 12796 41412 12798
rect 40236 12402 40404 12404
rect 40236 12350 40238 12402
rect 40290 12350 40404 12402
rect 40236 12348 40404 12350
rect 41132 12404 41188 12414
rect 41356 12404 41412 12796
rect 41132 12402 41412 12404
rect 41132 12350 41134 12402
rect 41186 12350 41412 12402
rect 41132 12348 41412 12350
rect 41804 12404 41860 12442
rect 40236 12338 40292 12348
rect 41132 12338 41188 12348
rect 41804 12338 41860 12348
rect 41804 12180 41860 12190
rect 41580 11282 41636 11294
rect 41580 11230 41582 11282
rect 41634 11230 41636 11282
rect 41580 11172 41636 11230
rect 41580 11106 41636 11116
rect 39900 9828 39956 9838
rect 39900 9734 39956 9772
rect 40684 9826 40740 9838
rect 40684 9774 40686 9826
rect 40738 9774 40740 9826
rect 39452 9662 39454 9714
rect 39506 9662 39508 9714
rect 39452 9650 39508 9662
rect 40684 8428 40740 9774
rect 41580 9826 41636 9838
rect 41580 9774 41582 9826
rect 41634 9774 41636 9826
rect 41580 9268 41636 9774
rect 41580 9202 41636 9212
rect 41244 9156 41300 9166
rect 41244 9062 41300 9100
rect 41804 9154 41860 12124
rect 42028 12178 42084 12190
rect 42028 12126 42030 12178
rect 42082 12126 42084 12178
rect 42028 11172 42084 12126
rect 42140 11620 42196 12910
rect 43036 12964 43092 12974
rect 43036 12870 43092 12908
rect 45836 12964 45892 12974
rect 45836 12402 45892 12908
rect 45836 12350 45838 12402
rect 45890 12350 45892 12402
rect 45836 12338 45892 12350
rect 42364 12180 42420 12190
rect 42364 12086 42420 12124
rect 42812 12178 42868 12190
rect 42812 12126 42814 12178
rect 42866 12126 42868 12178
rect 42700 12068 42756 12078
rect 42812 12068 42868 12126
rect 42756 12012 42868 12068
rect 42700 12002 42756 12012
rect 42476 11620 42532 11630
rect 42140 11618 42532 11620
rect 42140 11566 42478 11618
rect 42530 11566 42532 11618
rect 42140 11564 42532 11566
rect 42476 11554 42532 11564
rect 42028 11106 42084 11116
rect 43372 9268 43428 9278
rect 43372 9174 43428 9212
rect 41804 9102 41806 9154
rect 41858 9102 41860 9154
rect 41804 9090 41860 9102
rect 41580 8932 41636 8942
rect 41580 8838 41636 8876
rect 40684 8372 40964 8428
rect 40908 8258 40964 8372
rect 40908 8206 40910 8258
rect 40962 8206 40964 8258
rect 40908 8194 40964 8206
rect 39340 7198 39342 7250
rect 39394 7198 39396 7250
rect 39340 7186 39396 7198
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 33740 6862 33742 6914
rect 33794 6862 33796 6914
rect 33740 6850 33796 6862
rect 32844 6638 32846 6690
rect 32898 6638 32900 6690
rect 32844 6626 32900 6638
rect 29148 6526 29150 6578
rect 29202 6526 29204 6578
rect 29148 6514 29204 6526
rect 28812 5742 28814 5794
rect 28866 5742 28868 5794
rect 28812 5730 28868 5742
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 28588 5070 28590 5122
rect 28642 5070 28644 5122
rect 28588 5058 28644 5070
rect 24892 4958 24894 5010
rect 24946 4958 24948 5010
rect 24892 4946 24948 4958
rect 24668 4398 24670 4450
rect 24722 4398 24724 4450
rect 24668 4386 24724 4398
rect 24108 4286 24110 4338
rect 24162 4286 24164 4338
rect 24108 4274 24164 4286
rect 20300 4172 20916 4228
rect 21196 4116 21252 4126
rect 21196 4022 21252 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 19852 3502 19854 3554
rect 19906 3502 19908 3554
rect 19852 3490 19908 3502
rect 19516 3390 19518 3442
rect 19570 3390 19572 3442
rect 19516 3378 19572 3390
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
<< via2 >>
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 1708 43762 1764 43764
rect 1708 43710 1710 43762
rect 1710 43710 1762 43762
rect 1762 43710 1764 43762
rect 1708 43708 1764 43710
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 1708 42530 1764 42532
rect 1708 42478 1710 42530
rect 1710 42478 1762 42530
rect 1762 42478 1764 42530
rect 1708 42476 1764 42478
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 11900 40572 11956 40628
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 7644 39340 7700 39396
rect 2044 36316 2100 36372
rect 1708 34300 1764 34356
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 5180 36092 5236 36148
rect 4844 35868 4900 35924
rect 3164 35644 3220 35700
rect 3836 35698 3892 35700
rect 3836 35646 3838 35698
rect 3838 35646 3890 35698
rect 3890 35646 3892 35698
rect 3836 35644 3892 35646
rect 3500 35420 3556 35476
rect 3052 35026 3108 35028
rect 3052 34974 3054 35026
rect 3054 34974 3106 35026
rect 3106 34974 3108 35026
rect 3052 34972 3108 34974
rect 4508 35698 4564 35700
rect 4508 35646 4510 35698
rect 4510 35646 4562 35698
rect 4562 35646 4564 35698
rect 4508 35644 4564 35646
rect 2492 34300 2548 34356
rect 2156 33516 2212 33572
rect 2044 33180 2100 33236
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4956 35084 5012 35140
rect 4396 34690 4452 34692
rect 4396 34638 4398 34690
rect 4398 34638 4450 34690
rect 4450 34638 4452 34690
rect 4396 34636 4452 34638
rect 4284 33852 4340 33908
rect 4172 33570 4228 33572
rect 4172 33518 4174 33570
rect 4174 33518 4226 33570
rect 4226 33518 4228 33570
rect 4172 33516 4228 33518
rect 4060 33404 4116 33460
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 5404 34972 5460 35028
rect 5516 36204 5572 36260
rect 5516 35644 5572 35700
rect 5964 36092 6020 36148
rect 5628 35532 5684 35588
rect 6300 36370 6356 36372
rect 6300 36318 6302 36370
rect 6302 36318 6354 36370
rect 6354 36318 6356 36370
rect 6300 36316 6356 36318
rect 6972 36258 7028 36260
rect 6972 36206 6974 36258
rect 6974 36206 7026 36258
rect 7026 36206 7028 36258
rect 6972 36204 7028 36206
rect 6748 36092 6804 36148
rect 6748 35922 6804 35924
rect 6748 35870 6750 35922
rect 6750 35870 6802 35922
rect 6802 35870 6804 35922
rect 6748 35868 6804 35870
rect 11452 40236 11508 40292
rect 12124 40124 12180 40180
rect 9212 38892 9268 38948
rect 11228 39004 11284 39060
rect 9436 36482 9492 36484
rect 9436 36430 9438 36482
rect 9438 36430 9490 36482
rect 9490 36430 9492 36482
rect 9436 36428 9492 36430
rect 9660 36370 9716 36372
rect 9660 36318 9662 36370
rect 9662 36318 9714 36370
rect 9714 36318 9716 36370
rect 9660 36316 9716 36318
rect 10108 36316 10164 36372
rect 7980 36092 8036 36148
rect 6076 35084 6132 35140
rect 6188 35420 6244 35476
rect 5068 34690 5124 34692
rect 5068 34638 5070 34690
rect 5070 34638 5122 34690
rect 5122 34638 5124 34690
rect 5068 34636 5124 34638
rect 5964 34636 6020 34692
rect 5292 33906 5348 33908
rect 5292 33854 5294 33906
rect 5294 33854 5346 33906
rect 5346 33854 5348 33906
rect 5292 33852 5348 33854
rect 4844 33292 4900 33348
rect 3724 33234 3780 33236
rect 3724 33182 3726 33234
rect 3726 33182 3778 33234
rect 3778 33182 3780 33234
rect 3724 33180 3780 33182
rect 3724 32956 3780 33012
rect 3836 32732 3892 32788
rect 5628 33346 5684 33348
rect 5628 33294 5630 33346
rect 5630 33294 5682 33346
rect 5682 33294 5684 33346
rect 5628 33292 5684 33294
rect 6076 33852 6132 33908
rect 6636 33852 6692 33908
rect 6188 33404 6244 33460
rect 4844 32956 4900 33012
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 3948 31666 4004 31668
rect 3948 31614 3950 31666
rect 3950 31614 4002 31666
rect 4002 31614 4004 31666
rect 3948 31612 4004 31614
rect 2492 31500 2548 31556
rect 3836 31554 3892 31556
rect 3836 31502 3838 31554
rect 3838 31502 3890 31554
rect 3890 31502 3892 31554
rect 3836 31500 3892 31502
rect 5404 32786 5460 32788
rect 5404 32734 5406 32786
rect 5406 32734 5458 32786
rect 5458 32734 5460 32786
rect 5404 32732 5460 32734
rect 6972 32732 7028 32788
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 2268 30156 2324 30212
rect 3724 30210 3780 30212
rect 3724 30158 3726 30210
rect 3726 30158 3778 30210
rect 3778 30158 3780 30210
rect 3724 30156 3780 30158
rect 3836 30098 3892 30100
rect 3836 30046 3838 30098
rect 3838 30046 3890 30098
rect 3890 30046 3892 30098
rect 3836 30044 3892 30046
rect 5516 31612 5572 31668
rect 5404 30044 5460 30100
rect 5068 29596 5124 29652
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 1820 28588 1876 28644
rect 2268 28588 2324 28644
rect 5628 29650 5684 29652
rect 5628 29598 5630 29650
rect 5630 29598 5682 29650
rect 5682 29598 5684 29650
rect 5628 29596 5684 29598
rect 4284 28028 4340 28084
rect 4732 27916 4788 27972
rect 1932 27580 1988 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 1932 27186 1988 27188
rect 1932 27134 1934 27186
rect 1934 27134 1986 27186
rect 1986 27134 1988 27186
rect 1932 27132 1988 27134
rect 4284 27074 4340 27076
rect 4284 27022 4286 27074
rect 4286 27022 4338 27074
rect 4338 27022 4340 27074
rect 4284 27020 4340 27022
rect 2380 26908 2436 26964
rect 3164 26908 3220 26964
rect 1932 26236 1988 26292
rect 4620 26962 4676 26964
rect 4620 26910 4622 26962
rect 4622 26910 4674 26962
rect 4674 26910 4676 26962
rect 4620 26908 4676 26910
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 5628 28642 5684 28644
rect 5628 28590 5630 28642
rect 5630 28590 5682 28642
rect 5682 28590 5684 28642
rect 5628 28588 5684 28590
rect 6636 27970 6692 27972
rect 6636 27918 6638 27970
rect 6638 27918 6690 27970
rect 6690 27918 6692 27970
rect 6636 27916 6692 27918
rect 5068 26012 5124 26068
rect 4844 25788 4900 25844
rect 2716 25676 2772 25732
rect 4620 25730 4676 25732
rect 4620 25678 4622 25730
rect 4622 25678 4674 25730
rect 4674 25678 4676 25730
rect 4620 25676 4676 25678
rect 2828 25564 2884 25620
rect 1820 24610 1876 24612
rect 1820 24558 1822 24610
rect 1822 24558 1874 24610
rect 1874 24558 1876 24610
rect 1820 24556 1876 24558
rect 2044 24220 2100 24276
rect 4284 25564 4340 25620
rect 4732 25394 4788 25396
rect 4732 25342 4734 25394
rect 4734 25342 4786 25394
rect 4786 25342 4788 25394
rect 4732 25340 4788 25342
rect 6972 26012 7028 26068
rect 6188 25788 6244 25844
rect 5852 25228 5908 25284
rect 6636 25452 6692 25508
rect 7756 35474 7812 35476
rect 7756 35422 7758 35474
rect 7758 35422 7810 35474
rect 7810 35422 7812 35474
rect 7756 35420 7812 35422
rect 7868 35084 7924 35140
rect 10892 36316 10948 36372
rect 11676 38946 11732 38948
rect 11676 38894 11678 38946
rect 11678 38894 11730 38946
rect 11730 38894 11732 38946
rect 11676 38892 11732 38894
rect 12908 40348 12964 40404
rect 12796 40236 12852 40292
rect 12572 38892 12628 38948
rect 12908 39228 12964 39284
rect 12796 37996 12852 38052
rect 13580 42028 13636 42084
rect 13692 41186 13748 41188
rect 13692 41134 13694 41186
rect 13694 41134 13746 41186
rect 13746 41134 13748 41186
rect 13692 41132 13748 41134
rect 13468 40236 13524 40292
rect 13692 40348 13748 40404
rect 13468 38892 13524 38948
rect 13020 37436 13076 37492
rect 13692 39228 13748 39284
rect 17388 42028 17444 42084
rect 16044 41858 16100 41860
rect 16044 41806 16046 41858
rect 16046 41806 16098 41858
rect 16098 41806 16100 41858
rect 16044 41804 16100 41806
rect 22876 43484 22932 43540
rect 19852 42588 19908 42644
rect 20188 42476 20244 42532
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19516 42140 19572 42196
rect 17948 41804 18004 41860
rect 16044 40572 16100 40628
rect 15148 40460 15204 40516
rect 14588 40348 14644 40404
rect 14364 40124 14420 40180
rect 14364 39618 14420 39620
rect 14364 39566 14366 39618
rect 14366 39566 14418 39618
rect 14418 39566 14420 39618
rect 14364 39564 14420 39566
rect 15036 40236 15092 40292
rect 15932 40236 15988 40292
rect 15372 39452 15428 39508
rect 14364 38892 14420 38948
rect 13804 38722 13860 38724
rect 13804 38670 13806 38722
rect 13806 38670 13858 38722
rect 13858 38670 13860 38722
rect 13804 38668 13860 38670
rect 15260 39394 15316 39396
rect 15260 39342 15262 39394
rect 15262 39342 15314 39394
rect 15314 39342 15316 39394
rect 15260 39340 15316 39342
rect 15036 38780 15092 38836
rect 11116 36428 11172 36484
rect 10780 36204 10836 36260
rect 8540 35532 8596 35588
rect 8204 35308 8260 35364
rect 8204 34748 8260 34804
rect 9212 35138 9268 35140
rect 9212 35086 9214 35138
rect 9214 35086 9266 35138
rect 9266 35086 9268 35138
rect 9212 35084 9268 35086
rect 8540 34748 8596 34804
rect 9884 34748 9940 34804
rect 8316 34636 8372 34692
rect 9548 33906 9604 33908
rect 9548 33854 9550 33906
rect 9550 33854 9602 33906
rect 9602 33854 9604 33906
rect 9548 33852 9604 33854
rect 9548 33180 9604 33236
rect 8652 33068 8708 33124
rect 8540 32786 8596 32788
rect 8540 32734 8542 32786
rect 8542 32734 8594 32786
rect 8594 32734 8596 32786
rect 8540 32732 8596 32734
rect 7420 31164 7476 31220
rect 8316 31500 8372 31556
rect 8204 31218 8260 31220
rect 8204 31166 8206 31218
rect 8206 31166 8258 31218
rect 8258 31166 8260 31218
rect 8204 31164 8260 31166
rect 9212 31500 9268 31556
rect 7756 26236 7812 26292
rect 8204 26290 8260 26292
rect 8204 26238 8206 26290
rect 8206 26238 8258 26290
rect 8258 26238 8260 26290
rect 8204 26236 8260 26238
rect 8092 25788 8148 25844
rect 7756 25506 7812 25508
rect 7756 25454 7758 25506
rect 7758 25454 7810 25506
rect 7810 25454 7812 25506
rect 7756 25452 7812 25454
rect 4284 24780 4340 24836
rect 6972 24834 7028 24836
rect 6972 24782 6974 24834
rect 6974 24782 7026 24834
rect 7026 24782 7028 24834
rect 6972 24780 7028 24782
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 2380 22988 2436 23044
rect 1708 21532 1764 21588
rect 1708 20130 1764 20132
rect 1708 20078 1710 20130
rect 1710 20078 1762 20130
rect 1762 20078 1764 20130
rect 1708 20076 1764 20078
rect 1820 20860 1876 20916
rect 2716 22876 2772 22932
rect 1932 20188 1988 20244
rect 1708 18508 1764 18564
rect 2044 19740 2100 19796
rect 1932 19068 1988 19124
rect 1820 18844 1876 18900
rect 1708 18172 1764 18228
rect 1708 17724 1764 17780
rect 1708 17388 1764 17444
rect 5852 24610 5908 24612
rect 5852 24558 5854 24610
rect 5854 24558 5906 24610
rect 5906 24558 5908 24610
rect 5852 24556 5908 24558
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4732 22370 4788 22372
rect 4732 22318 4734 22370
rect 4734 22318 4786 22370
rect 4786 22318 4788 22370
rect 4732 22316 4788 22318
rect 4284 22092 4340 22148
rect 4956 23324 5012 23380
rect 6188 23772 6244 23828
rect 5852 23378 5908 23380
rect 5852 23326 5854 23378
rect 5854 23326 5906 23378
rect 5906 23326 5908 23378
rect 5852 23324 5908 23326
rect 6636 23714 6692 23716
rect 6636 23662 6638 23714
rect 6638 23662 6690 23714
rect 6690 23662 6692 23714
rect 6636 23660 6692 23662
rect 6412 23324 6468 23380
rect 6972 23436 7028 23492
rect 6860 23212 6916 23268
rect 5964 22370 6020 22372
rect 5964 22318 5966 22370
rect 5966 22318 6018 22370
rect 6018 22318 6020 22370
rect 5964 22316 6020 22318
rect 6412 22316 6468 22372
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4284 20412 4340 20468
rect 3164 20188 3220 20244
rect 2268 19234 2324 19236
rect 2268 19182 2270 19234
rect 2270 19182 2322 19234
rect 2322 19182 2324 19234
rect 2268 19180 2324 19182
rect 2156 18732 2212 18788
rect 2156 18508 2212 18564
rect 2268 18338 2324 18340
rect 2268 18286 2270 18338
rect 2270 18286 2322 18338
rect 2322 18286 2324 18338
rect 2268 18284 2324 18286
rect 2044 17442 2100 17444
rect 2044 17390 2046 17442
rect 2046 17390 2098 17442
rect 2098 17390 2100 17442
rect 2044 17388 2100 17390
rect 2156 16268 2212 16324
rect 1820 15148 1876 15204
rect 2940 19404 2996 19460
rect 2604 19122 2660 19124
rect 2604 19070 2606 19122
rect 2606 19070 2658 19122
rect 2658 19070 2660 19122
rect 2604 19068 2660 19070
rect 4172 19852 4228 19908
rect 3500 19516 3556 19572
rect 2380 17836 2436 17892
rect 3836 19010 3892 19012
rect 3836 18958 3838 19010
rect 3838 18958 3890 19010
rect 3890 18958 3892 19010
rect 3836 18956 3892 18958
rect 3388 18450 3444 18452
rect 3388 18398 3390 18450
rect 3390 18398 3442 18450
rect 3442 18398 3444 18450
rect 3388 18396 3444 18398
rect 4060 17890 4116 17892
rect 4060 17838 4062 17890
rect 4062 17838 4114 17890
rect 4114 17838 4116 17890
rect 4060 17836 4116 17838
rect 3500 17666 3556 17668
rect 3500 17614 3502 17666
rect 3502 17614 3554 17666
rect 3554 17614 3556 17666
rect 3500 17612 3556 17614
rect 3612 17554 3668 17556
rect 3612 17502 3614 17554
rect 3614 17502 3666 17554
rect 3666 17502 3668 17554
rect 3612 17500 3668 17502
rect 2716 17442 2772 17444
rect 2716 17390 2718 17442
rect 2718 17390 2770 17442
rect 2770 17390 2772 17442
rect 2716 17388 2772 17390
rect 4172 17164 4228 17220
rect 2380 16828 2436 16884
rect 3500 16322 3556 16324
rect 3500 16270 3502 16322
rect 3502 16270 3554 16322
rect 3554 16270 3556 16322
rect 3500 16268 3556 16270
rect 3500 15202 3556 15204
rect 3500 15150 3502 15202
rect 3502 15150 3554 15202
rect 3554 15150 3556 15202
rect 3500 15148 3556 15150
rect 3724 13916 3780 13972
rect 5068 20578 5124 20580
rect 5068 20526 5070 20578
rect 5070 20526 5122 20578
rect 5122 20526 5124 20578
rect 5068 20524 5124 20526
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4508 19458 4564 19460
rect 4508 19406 4510 19458
rect 4510 19406 4562 19458
rect 4562 19406 4564 19458
rect 4508 19404 4564 19406
rect 7084 22258 7140 22260
rect 7084 22206 7086 22258
rect 7086 22206 7138 22258
rect 7138 22206 7140 22258
rect 7084 22204 7140 22206
rect 6300 20802 6356 20804
rect 6300 20750 6302 20802
rect 6302 20750 6354 20802
rect 6354 20750 6356 20802
rect 6300 20748 6356 20750
rect 5964 20412 6020 20468
rect 6636 20578 6692 20580
rect 6636 20526 6638 20578
rect 6638 20526 6690 20578
rect 6690 20526 6692 20578
rect 6636 20524 6692 20526
rect 5628 19852 5684 19908
rect 4844 19404 4900 19460
rect 4620 19346 4676 19348
rect 4620 19294 4622 19346
rect 4622 19294 4674 19346
rect 4674 19294 4676 19346
rect 4620 19292 4676 19294
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4620 17778 4676 17780
rect 4620 17726 4622 17778
rect 4622 17726 4674 17778
rect 4674 17726 4676 17778
rect 4620 17724 4676 17726
rect 6860 20412 6916 20468
rect 6076 19292 6132 19348
rect 7644 23378 7700 23380
rect 7644 23326 7646 23378
rect 7646 23326 7698 23378
rect 7698 23326 7700 23378
rect 7644 23324 7700 23326
rect 8540 26124 8596 26180
rect 8652 26236 8708 26292
rect 9212 26012 9268 26068
rect 8428 24834 8484 24836
rect 8428 24782 8430 24834
rect 8430 24782 8482 24834
rect 8482 24782 8484 24834
rect 8428 24780 8484 24782
rect 7980 24556 8036 24612
rect 8876 24556 8932 24612
rect 8652 23826 8708 23828
rect 8652 23774 8654 23826
rect 8654 23774 8706 23826
rect 8706 23774 8708 23826
rect 8652 23772 8708 23774
rect 8988 23772 9044 23828
rect 9548 28418 9604 28420
rect 9548 28366 9550 28418
rect 9550 28366 9602 28418
rect 9602 28366 9604 28418
rect 9548 28364 9604 28366
rect 9548 27020 9604 27076
rect 11228 36204 11284 36260
rect 12908 36092 12964 36148
rect 13692 36594 13748 36596
rect 13692 36542 13694 36594
rect 13694 36542 13746 36594
rect 13746 36542 13748 36594
rect 13692 36540 13748 36542
rect 14252 37436 14308 37492
rect 14700 37490 14756 37492
rect 14700 37438 14702 37490
rect 14702 37438 14754 37490
rect 14754 37438 14756 37490
rect 14700 37436 14756 37438
rect 14588 37212 14644 37268
rect 14364 35980 14420 36036
rect 13020 34972 13076 35028
rect 10556 33404 10612 33460
rect 10332 33234 10388 33236
rect 10332 33182 10334 33234
rect 10334 33182 10386 33234
rect 10386 33182 10388 33234
rect 10332 33180 10388 33182
rect 10108 33122 10164 33124
rect 10108 33070 10110 33122
rect 10110 33070 10162 33122
rect 10162 33070 10164 33122
rect 10108 33068 10164 33070
rect 10556 32396 10612 32452
rect 10444 31554 10500 31556
rect 10444 31502 10446 31554
rect 10446 31502 10498 31554
rect 10498 31502 10500 31554
rect 10444 31500 10500 31502
rect 10108 28530 10164 28532
rect 10108 28478 10110 28530
rect 10110 28478 10162 28530
rect 10162 28478 10164 28530
rect 10108 28476 10164 28478
rect 9884 27356 9940 27412
rect 10444 28364 10500 28420
rect 10220 28082 10276 28084
rect 10220 28030 10222 28082
rect 10222 28030 10274 28082
rect 10274 28030 10276 28082
rect 10220 28028 10276 28030
rect 9996 26962 10052 26964
rect 9996 26910 9998 26962
rect 9998 26910 10050 26962
rect 10050 26910 10052 26962
rect 9996 26908 10052 26910
rect 11340 33404 11396 33460
rect 12796 33516 12852 33572
rect 13356 33404 13412 33460
rect 11676 32620 11732 32676
rect 11564 32450 11620 32452
rect 11564 32398 11566 32450
rect 11566 32398 11618 32450
rect 11618 32398 11620 32450
rect 11564 32396 11620 32398
rect 11564 31778 11620 31780
rect 11564 31726 11566 31778
rect 11566 31726 11618 31778
rect 11618 31726 11620 31778
rect 11564 31724 11620 31726
rect 11228 31612 11284 31668
rect 10780 30156 10836 30212
rect 12012 32396 12068 32452
rect 12572 32562 12628 32564
rect 12572 32510 12574 32562
rect 12574 32510 12626 32562
rect 12626 32510 12628 32562
rect 12572 32508 12628 32510
rect 12908 32172 12964 32228
rect 12236 31724 12292 31780
rect 11900 31666 11956 31668
rect 11900 31614 11902 31666
rect 11902 31614 11954 31666
rect 11954 31614 11956 31666
rect 11900 31612 11956 31614
rect 12236 30940 12292 30996
rect 11676 29036 11732 29092
rect 12124 30210 12180 30212
rect 12124 30158 12126 30210
rect 12126 30158 12178 30210
rect 12178 30158 12180 30210
rect 12124 30156 12180 30158
rect 11452 28476 11508 28532
rect 11788 27020 11844 27076
rect 10220 26402 10276 26404
rect 10220 26350 10222 26402
rect 10222 26350 10274 26402
rect 10274 26350 10276 26402
rect 10220 26348 10276 26350
rect 9996 26290 10052 26292
rect 9996 26238 9998 26290
rect 9998 26238 10050 26290
rect 10050 26238 10052 26290
rect 9996 26236 10052 26238
rect 9996 26012 10052 26068
rect 8540 22988 8596 23044
rect 9660 23826 9716 23828
rect 9660 23774 9662 23826
rect 9662 23774 9714 23826
rect 9714 23774 9716 23826
rect 9660 23772 9716 23774
rect 9996 24668 10052 24724
rect 9436 23212 9492 23268
rect 9884 23212 9940 23268
rect 7420 21698 7476 21700
rect 7420 21646 7422 21698
rect 7422 21646 7474 21698
rect 7474 21646 7476 21698
rect 7420 21644 7476 21646
rect 8428 22370 8484 22372
rect 8428 22318 8430 22370
rect 8430 22318 8482 22370
rect 8482 22318 8484 22370
rect 8428 22316 8484 22318
rect 8204 22146 8260 22148
rect 8204 22094 8206 22146
rect 8206 22094 8258 22146
rect 8258 22094 8260 22146
rect 8204 22092 8260 22094
rect 8092 21810 8148 21812
rect 8092 21758 8094 21810
rect 8094 21758 8146 21810
rect 8146 21758 8148 21810
rect 8092 21756 8148 21758
rect 7532 21532 7588 21588
rect 7532 20748 7588 20804
rect 7644 20412 7700 20468
rect 9884 20524 9940 20580
rect 4956 18732 5012 18788
rect 4956 18396 5012 18452
rect 5180 18172 5236 18228
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 6412 20018 6468 20020
rect 6412 19966 6414 20018
rect 6414 19966 6466 20018
rect 6466 19966 6468 20018
rect 6412 19964 6468 19966
rect 7196 19404 7252 19460
rect 6748 19292 6804 19348
rect 6636 19122 6692 19124
rect 6636 19070 6638 19122
rect 6638 19070 6690 19122
rect 6690 19070 6692 19122
rect 6636 19068 6692 19070
rect 6076 17666 6132 17668
rect 6076 17614 6078 17666
rect 6078 17614 6130 17666
rect 6130 17614 6132 17666
rect 6076 17612 6132 17614
rect 5628 17164 5684 17220
rect 6748 18284 6804 18340
rect 6412 18226 6468 18228
rect 6412 18174 6414 18226
rect 6414 18174 6466 18226
rect 6466 18174 6468 18226
rect 6412 18172 6468 18174
rect 8876 20018 8932 20020
rect 8876 19966 8878 20018
rect 8878 19966 8930 20018
rect 8930 19966 8932 20018
rect 8876 19964 8932 19966
rect 8764 19740 8820 19796
rect 7308 18172 7364 18228
rect 8092 17836 8148 17892
rect 6188 17164 6244 17220
rect 10220 21756 10276 21812
rect 10220 21308 10276 21364
rect 10556 25116 10612 25172
rect 11116 26962 11172 26964
rect 11116 26910 11118 26962
rect 11118 26910 11170 26962
rect 11170 26910 11172 26962
rect 11116 26908 11172 26910
rect 11004 26348 11060 26404
rect 11676 26348 11732 26404
rect 10892 25340 10948 25396
rect 10780 25228 10836 25284
rect 11340 24834 11396 24836
rect 11340 24782 11342 24834
rect 11342 24782 11394 24834
rect 11394 24782 11396 24834
rect 11340 24780 11396 24782
rect 10780 24332 10836 24388
rect 10444 23436 10500 23492
rect 10444 23154 10500 23156
rect 10444 23102 10446 23154
rect 10446 23102 10498 23154
rect 10498 23102 10500 23154
rect 10444 23100 10500 23102
rect 10668 23266 10724 23268
rect 10668 23214 10670 23266
rect 10670 23214 10722 23266
rect 10722 23214 10724 23266
rect 10668 23212 10724 23214
rect 10780 23100 10836 23156
rect 11900 24556 11956 24612
rect 12012 24108 12068 24164
rect 11900 23548 11956 23604
rect 11004 21586 11060 21588
rect 11004 21534 11006 21586
rect 11006 21534 11058 21586
rect 11058 21534 11060 21586
rect 11004 21532 11060 21534
rect 10556 20914 10612 20916
rect 10556 20862 10558 20914
rect 10558 20862 10610 20914
rect 10610 20862 10612 20914
rect 10556 20860 10612 20862
rect 11004 20578 11060 20580
rect 11004 20526 11006 20578
rect 11006 20526 11058 20578
rect 11058 20526 11060 20578
rect 11004 20524 11060 20526
rect 11676 22540 11732 22596
rect 13916 33404 13972 33460
rect 13692 32508 13748 32564
rect 13580 32172 13636 32228
rect 13692 31948 13748 32004
rect 13580 31612 13636 31668
rect 13356 30156 13412 30212
rect 12796 30044 12852 30100
rect 13468 30044 13524 30100
rect 12348 27468 12404 27524
rect 14588 35084 14644 35140
rect 14476 34972 14532 35028
rect 15148 37324 15204 37380
rect 15036 36988 15092 37044
rect 15260 36988 15316 37044
rect 15372 38892 15428 38948
rect 15148 36876 15204 36932
rect 15596 39618 15652 39620
rect 15596 39566 15598 39618
rect 15598 39566 15650 39618
rect 15650 39566 15652 39618
rect 15596 39564 15652 39566
rect 15484 38780 15540 38836
rect 15596 38050 15652 38052
rect 15596 37998 15598 38050
rect 15598 37998 15650 38050
rect 15650 37998 15652 38050
rect 15596 37996 15652 37998
rect 15708 37266 15764 37268
rect 15708 37214 15710 37266
rect 15710 37214 15762 37266
rect 15762 37214 15764 37266
rect 15708 37212 15764 37214
rect 14476 32844 14532 32900
rect 14924 33404 14980 33460
rect 14700 32508 14756 32564
rect 14476 31554 14532 31556
rect 14476 31502 14478 31554
rect 14478 31502 14530 31554
rect 14530 31502 14532 31554
rect 14476 31500 14532 31502
rect 13916 29484 13972 29540
rect 14140 29260 14196 29316
rect 14140 29036 14196 29092
rect 13244 27244 13300 27300
rect 13692 27356 13748 27412
rect 12684 27132 12740 27188
rect 12460 25564 12516 25620
rect 13804 27244 13860 27300
rect 15036 33292 15092 33348
rect 15036 31948 15092 32004
rect 15484 36594 15540 36596
rect 15484 36542 15486 36594
rect 15486 36542 15538 36594
rect 15538 36542 15540 36594
rect 15484 36540 15540 36542
rect 15260 36370 15316 36372
rect 15260 36318 15262 36370
rect 15262 36318 15314 36370
rect 15314 36318 15316 36370
rect 15260 36316 15316 36318
rect 15372 36258 15428 36260
rect 15372 36206 15374 36258
rect 15374 36206 15426 36258
rect 15426 36206 15428 36258
rect 15372 36204 15428 36206
rect 15596 35420 15652 35476
rect 15372 34914 15428 34916
rect 15372 34862 15374 34914
rect 15374 34862 15426 34914
rect 15426 34862 15428 34914
rect 15372 34860 15428 34862
rect 15596 34242 15652 34244
rect 15596 34190 15598 34242
rect 15598 34190 15650 34242
rect 15650 34190 15652 34242
rect 15596 34188 15652 34190
rect 15372 31666 15428 31668
rect 15372 31614 15374 31666
rect 15374 31614 15426 31666
rect 15426 31614 15428 31666
rect 15372 31612 15428 31614
rect 15036 31106 15092 31108
rect 15036 31054 15038 31106
rect 15038 31054 15090 31106
rect 15090 31054 15092 31106
rect 15036 31052 15092 31054
rect 14924 29596 14980 29652
rect 15372 31276 15428 31332
rect 14924 29036 14980 29092
rect 14812 27244 14868 27300
rect 15820 36764 15876 36820
rect 16492 40460 16548 40516
rect 16156 40236 16212 40292
rect 16268 38834 16324 38836
rect 16268 38782 16270 38834
rect 16270 38782 16322 38834
rect 16322 38782 16324 38834
rect 16268 38780 16324 38782
rect 16492 38220 16548 38276
rect 16380 37212 16436 37268
rect 16492 36988 16548 37044
rect 17388 40402 17444 40404
rect 17388 40350 17390 40402
rect 17390 40350 17442 40402
rect 17442 40350 17444 40402
rect 17388 40348 17444 40350
rect 18508 41132 18564 41188
rect 19404 41132 19460 41188
rect 17948 40684 18004 40740
rect 17500 39564 17556 39620
rect 16716 38946 16772 38948
rect 16716 38894 16718 38946
rect 16718 38894 16770 38946
rect 16770 38894 16772 38946
rect 16716 38892 16772 38894
rect 16828 38780 16884 38836
rect 17388 38722 17444 38724
rect 17388 38670 17390 38722
rect 17390 38670 17442 38722
rect 17442 38670 17444 38722
rect 17388 38668 17444 38670
rect 17724 37324 17780 37380
rect 17836 38780 17892 38836
rect 19628 41132 19684 41188
rect 19836 40794 19892 40796
rect 19628 40684 19684 40740
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19180 39676 19236 39732
rect 17836 37266 17892 37268
rect 17836 37214 17838 37266
rect 17838 37214 17890 37266
rect 17890 37214 17892 37266
rect 17836 37212 17892 37214
rect 16604 37100 16660 37156
rect 17388 37154 17444 37156
rect 17388 37102 17390 37154
rect 17390 37102 17442 37154
rect 17442 37102 17444 37154
rect 17388 37100 17444 37102
rect 17612 36764 17668 36820
rect 16492 36092 16548 36148
rect 16604 35980 16660 36036
rect 16156 34242 16212 34244
rect 16156 34190 16158 34242
rect 16158 34190 16210 34242
rect 16210 34190 16212 34242
rect 16156 34188 16212 34190
rect 16044 33628 16100 33684
rect 15820 33516 15876 33572
rect 16156 32844 16212 32900
rect 15484 30156 15540 30212
rect 12796 25282 12852 25284
rect 12796 25230 12798 25282
rect 12798 25230 12850 25282
rect 12850 25230 12852 25282
rect 12796 25228 12852 25230
rect 14028 25116 14084 25172
rect 12348 24834 12404 24836
rect 12348 24782 12350 24834
rect 12350 24782 12402 24834
rect 12402 24782 12404 24834
rect 12348 24780 12404 24782
rect 14476 24892 14532 24948
rect 13244 24722 13300 24724
rect 13244 24670 13246 24722
rect 13246 24670 13298 24722
rect 13298 24670 13300 24722
rect 13244 24668 13300 24670
rect 13020 23884 13076 23940
rect 14252 23884 14308 23940
rect 12796 23548 12852 23604
rect 12572 23436 12628 23492
rect 12908 23436 12964 23492
rect 12236 22540 12292 22596
rect 11676 21756 11732 21812
rect 10108 19516 10164 19572
rect 8988 18396 9044 18452
rect 9212 17554 9268 17556
rect 9212 17502 9214 17554
rect 9214 17502 9266 17554
rect 9266 17502 9268 17554
rect 9212 17500 9268 17502
rect 8428 17106 8484 17108
rect 8428 17054 8430 17106
rect 8430 17054 8482 17106
rect 8482 17054 8484 17106
rect 8428 17052 8484 17054
rect 8540 17164 8596 17220
rect 5516 16268 5572 16324
rect 6076 16828 6132 16884
rect 9660 17948 9716 18004
rect 9548 17164 9604 17220
rect 8204 16716 8260 16772
rect 9100 16882 9156 16884
rect 9100 16830 9102 16882
rect 9102 16830 9154 16882
rect 9154 16830 9156 16882
rect 9100 16828 9156 16830
rect 8988 16716 9044 16772
rect 9660 16716 9716 16772
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 5068 15314 5124 15316
rect 5068 15262 5070 15314
rect 5070 15262 5122 15314
rect 5122 15262 5124 15314
rect 5068 15260 5124 15262
rect 4844 14530 4900 14532
rect 4844 14478 4846 14530
rect 4846 14478 4898 14530
rect 4898 14478 4900 14530
rect 4844 14476 4900 14478
rect 5964 15260 6020 15316
rect 7308 15148 7364 15204
rect 7980 14530 8036 14532
rect 7980 14478 7982 14530
rect 7982 14478 8034 14530
rect 8034 14478 8036 14530
rect 7980 14476 8036 14478
rect 9100 15538 9156 15540
rect 9100 15486 9102 15538
rect 9102 15486 9154 15538
rect 9154 15486 9156 15538
rect 9100 15484 9156 15486
rect 8540 15202 8596 15204
rect 8540 15150 8542 15202
rect 8542 15150 8594 15202
rect 8594 15150 8596 15202
rect 8540 15148 8596 15150
rect 9660 15148 9716 15204
rect 10444 20076 10500 20132
rect 10556 19964 10612 20020
rect 12796 22204 12852 22260
rect 12460 22092 12516 22148
rect 11788 21532 11844 21588
rect 11340 20914 11396 20916
rect 11340 20862 11342 20914
rect 11342 20862 11394 20914
rect 11394 20862 11396 20914
rect 11340 20860 11396 20862
rect 10780 19516 10836 19572
rect 10668 19404 10724 19460
rect 10332 18450 10388 18452
rect 10332 18398 10334 18450
rect 10334 18398 10386 18450
rect 10386 18398 10388 18450
rect 10332 18396 10388 18398
rect 9996 16604 10052 16660
rect 10444 17948 10500 18004
rect 10668 17890 10724 17892
rect 10668 17838 10670 17890
rect 10670 17838 10722 17890
rect 10722 17838 10724 17890
rect 10668 17836 10724 17838
rect 11676 20130 11732 20132
rect 11676 20078 11678 20130
rect 11678 20078 11730 20130
rect 11730 20078 11732 20130
rect 11676 20076 11732 20078
rect 11452 20018 11508 20020
rect 11452 19966 11454 20018
rect 11454 19966 11506 20018
rect 11506 19966 11508 20018
rect 11452 19964 11508 19966
rect 11116 19794 11172 19796
rect 11116 19742 11118 19794
rect 11118 19742 11170 19794
rect 11170 19742 11172 19794
rect 11116 19740 11172 19742
rect 11340 19740 11396 19796
rect 10668 16828 10724 16884
rect 12012 19852 12068 19908
rect 12236 19852 12292 19908
rect 12348 19964 12404 20020
rect 11788 19516 11844 19572
rect 11564 17948 11620 18004
rect 11676 17612 11732 17668
rect 11564 17388 11620 17444
rect 11676 17276 11732 17332
rect 10220 15484 10276 15540
rect 11452 16770 11508 16772
rect 11452 16718 11454 16770
rect 11454 16718 11506 16770
rect 11506 16718 11508 16770
rect 11452 16716 11508 16718
rect 9884 14700 9940 14756
rect 10556 14588 10612 14644
rect 9548 14476 9604 14532
rect 1820 12684 1876 12740
rect 1820 11452 1876 11508
rect 3612 13468 3668 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 3500 12738 3556 12740
rect 3500 12686 3502 12738
rect 3502 12686 3554 12738
rect 3554 12686 3556 12738
rect 3500 12684 3556 12686
rect 5628 14252 5684 14308
rect 5292 13970 5348 13972
rect 5292 13918 5294 13970
rect 5294 13918 5346 13970
rect 5346 13918 5348 13970
rect 5292 13916 5348 13918
rect 7196 14306 7252 14308
rect 7196 14254 7198 14306
rect 7198 14254 7250 14306
rect 7250 14254 7252 14306
rect 7196 14252 7252 14254
rect 5068 13468 5124 13524
rect 12348 18844 12404 18900
rect 15148 24668 15204 24724
rect 14700 23938 14756 23940
rect 14700 23886 14702 23938
rect 14702 23886 14754 23938
rect 14754 23886 14756 23938
rect 14700 23884 14756 23886
rect 14364 23436 14420 23492
rect 14924 23436 14980 23492
rect 14476 23212 14532 23268
rect 13580 22146 13636 22148
rect 13580 22094 13582 22146
rect 13582 22094 13634 22146
rect 13634 22094 13636 22146
rect 13580 22092 13636 22094
rect 13916 23100 13972 23156
rect 13020 21868 13076 21924
rect 13132 21698 13188 21700
rect 13132 21646 13134 21698
rect 13134 21646 13186 21698
rect 13186 21646 13188 21698
rect 13132 21644 13188 21646
rect 13804 21868 13860 21924
rect 13580 21026 13636 21028
rect 13580 20974 13582 21026
rect 13582 20974 13634 21026
rect 13634 20974 13636 21026
rect 13580 20972 13636 20974
rect 13468 20860 13524 20916
rect 12572 20076 12628 20132
rect 12124 17612 12180 17668
rect 12124 16994 12180 16996
rect 12124 16942 12126 16994
rect 12126 16942 12178 16994
rect 12178 16942 12180 16994
rect 12124 16940 12180 16942
rect 12236 17500 12292 17556
rect 12796 20018 12852 20020
rect 12796 19966 12798 20018
rect 12798 19966 12850 20018
rect 12850 19966 12852 20018
rect 12796 19964 12852 19966
rect 13692 19964 13748 20020
rect 13580 19906 13636 19908
rect 13580 19854 13582 19906
rect 13582 19854 13634 19906
rect 13634 19854 13636 19906
rect 13580 19852 13636 19854
rect 13580 19628 13636 19684
rect 12796 19404 12852 19460
rect 12684 19180 12740 19236
rect 13468 19404 13524 19460
rect 13356 19068 13412 19124
rect 12796 18674 12852 18676
rect 12796 18622 12798 18674
rect 12798 18622 12850 18674
rect 12850 18622 12852 18674
rect 12796 18620 12852 18622
rect 13020 18732 13076 18788
rect 12908 18508 12964 18564
rect 13692 19292 13748 19348
rect 15036 23212 15092 23268
rect 14028 21644 14084 21700
rect 14700 21868 14756 21924
rect 14364 21474 14420 21476
rect 14364 21422 14366 21474
rect 14366 21422 14418 21474
rect 14418 21422 14420 21474
rect 14364 21420 14420 21422
rect 13804 19852 13860 19908
rect 13804 19180 13860 19236
rect 14140 20748 14196 20804
rect 13580 18956 13636 19012
rect 13804 19010 13860 19012
rect 13804 18958 13806 19010
rect 13806 18958 13858 19010
rect 13858 18958 13860 19010
rect 13804 18956 13860 18958
rect 12236 16492 12292 16548
rect 11788 15484 11844 15540
rect 12572 16604 12628 16660
rect 12684 16828 12740 16884
rect 12684 15986 12740 15988
rect 12684 15934 12686 15986
rect 12686 15934 12738 15986
rect 12738 15934 12740 15986
rect 12684 15932 12740 15934
rect 12572 15314 12628 15316
rect 12572 15262 12574 15314
rect 12574 15262 12626 15314
rect 12626 15262 12628 15314
rect 12572 15260 12628 15262
rect 8316 13692 8372 13748
rect 10332 13746 10388 13748
rect 10332 13694 10334 13746
rect 10334 13694 10386 13746
rect 10386 13694 10388 13746
rect 10332 13692 10388 13694
rect 6076 12684 6132 12740
rect 7308 12684 7364 12740
rect 4060 12124 4116 12180
rect 3612 11564 3668 11620
rect 3724 11900 3780 11956
rect 3500 11452 3556 11508
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 3724 10332 3780 10388
rect 2492 9996 2548 10052
rect 2044 9548 2100 9604
rect 1932 8988 1988 9044
rect 2940 9660 2996 9716
rect 5404 11954 5460 11956
rect 5404 11902 5406 11954
rect 5406 11902 5458 11954
rect 5458 11902 5460 11954
rect 5404 11900 5460 11902
rect 4844 11340 4900 11396
rect 4060 9996 4116 10052
rect 5292 11564 5348 11620
rect 5628 11394 5684 11396
rect 5628 11342 5630 11394
rect 5630 11342 5682 11394
rect 5682 11342 5684 11394
rect 5628 11340 5684 11342
rect 6076 11340 6132 11396
rect 6076 10556 6132 10612
rect 5180 10332 5236 10388
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4172 9772 4228 9828
rect 4172 9602 4228 9604
rect 4172 9550 4174 9602
rect 4174 9550 4226 9602
rect 4226 9550 4228 9602
rect 4172 9548 4228 9550
rect 4956 9714 5012 9716
rect 4956 9662 4958 9714
rect 4958 9662 5010 9714
rect 5010 9662 5012 9714
rect 4956 9660 5012 9662
rect 8540 12738 8596 12740
rect 8540 12686 8542 12738
rect 8542 12686 8594 12738
rect 8594 12686 8596 12738
rect 8540 12684 8596 12686
rect 12572 14700 12628 14756
rect 11900 14642 11956 14644
rect 11900 14590 11902 14642
rect 11902 14590 11954 14642
rect 11954 14590 11956 14642
rect 11900 14588 11956 14590
rect 11564 12236 11620 12292
rect 7980 11900 8036 11956
rect 8876 12178 8932 12180
rect 8876 12126 8878 12178
rect 8878 12126 8930 12178
rect 8930 12126 8932 12178
rect 8876 12124 8932 12126
rect 9548 11954 9604 11956
rect 9548 11902 9550 11954
rect 9550 11902 9602 11954
rect 9602 11902 9604 11954
rect 9548 11900 9604 11902
rect 9660 11564 9716 11620
rect 8428 11452 8484 11508
rect 6188 10332 6244 10388
rect 6636 10556 6692 10612
rect 4844 8988 4900 9044
rect 5516 9772 5572 9828
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4284 6860 4340 6916
rect 5964 9042 6020 9044
rect 5964 8990 5966 9042
rect 5966 8990 6018 9042
rect 6018 8990 6020 9042
rect 5964 8988 6020 8990
rect 8428 10610 8484 10612
rect 8428 10558 8430 10610
rect 8430 10558 8482 10610
rect 8482 10558 8484 10610
rect 8428 10556 8484 10558
rect 11340 11676 11396 11732
rect 11004 11618 11060 11620
rect 11004 11566 11006 11618
rect 11006 11566 11058 11618
rect 11058 11566 11060 11618
rect 11004 11564 11060 11566
rect 10332 11170 10388 11172
rect 10332 11118 10334 11170
rect 10334 11118 10386 11170
rect 10386 11118 10388 11170
rect 10332 11116 10388 11118
rect 10668 11116 10724 11172
rect 9100 10610 9156 10612
rect 9100 10558 9102 10610
rect 9102 10558 9154 10610
rect 9154 10558 9156 10610
rect 9100 10556 9156 10558
rect 9996 10610 10052 10612
rect 9996 10558 9998 10610
rect 9998 10558 10050 10610
rect 10050 10558 10052 10610
rect 9996 10556 10052 10558
rect 9884 10332 9940 10388
rect 12348 12124 12404 12180
rect 12348 11676 12404 11732
rect 12012 11394 12068 11396
rect 12012 11342 12014 11394
rect 12014 11342 12066 11394
rect 12066 11342 12068 11394
rect 12012 11340 12068 11342
rect 12236 10780 12292 10836
rect 12460 11116 12516 11172
rect 13244 18396 13300 18452
rect 12908 18338 12964 18340
rect 12908 18286 12910 18338
rect 12910 18286 12962 18338
rect 12962 18286 12964 18338
rect 12908 18284 12964 18286
rect 12908 17500 12964 17556
rect 13692 17666 13748 17668
rect 13692 17614 13694 17666
rect 13694 17614 13746 17666
rect 13746 17614 13748 17666
rect 13692 17612 13748 17614
rect 13580 17554 13636 17556
rect 13580 17502 13582 17554
rect 13582 17502 13634 17554
rect 13634 17502 13636 17554
rect 13580 17500 13636 17502
rect 13132 17052 13188 17108
rect 12908 16940 12964 16996
rect 14028 19068 14084 19124
rect 14924 21756 14980 21812
rect 15036 21868 15092 21924
rect 14812 20748 14868 20804
rect 15372 25116 15428 25172
rect 15372 23884 15428 23940
rect 15708 31106 15764 31108
rect 15708 31054 15710 31106
rect 15710 31054 15762 31106
rect 15762 31054 15764 31106
rect 15708 31052 15764 31054
rect 15820 30044 15876 30100
rect 16044 30994 16100 30996
rect 16044 30942 16046 30994
rect 16046 30942 16098 30994
rect 16098 30942 16100 30994
rect 16044 30940 16100 30942
rect 16828 34242 16884 34244
rect 16828 34190 16830 34242
rect 16830 34190 16882 34242
rect 16882 34190 16884 34242
rect 16828 34188 16884 34190
rect 16940 33516 16996 33572
rect 16604 31836 16660 31892
rect 16940 32284 16996 32340
rect 16380 30828 16436 30884
rect 16828 31052 16884 31108
rect 15932 29484 15988 29540
rect 15820 28476 15876 28532
rect 16268 26908 16324 26964
rect 15708 23938 15764 23940
rect 15708 23886 15710 23938
rect 15710 23886 15762 23938
rect 15762 23886 15764 23938
rect 15708 23884 15764 23886
rect 15372 23436 15428 23492
rect 15372 21980 15428 22036
rect 15708 23660 15764 23716
rect 14924 20972 14980 21028
rect 14924 20636 14980 20692
rect 14028 18674 14084 18676
rect 14028 18622 14030 18674
rect 14030 18622 14082 18674
rect 14082 18622 14084 18674
rect 14028 18620 14084 18622
rect 14252 19740 14308 19796
rect 14476 19404 14532 19460
rect 14700 18450 14756 18452
rect 14700 18398 14702 18450
rect 14702 18398 14754 18450
rect 14754 18398 14756 18450
rect 14700 18396 14756 18398
rect 13916 16828 13972 16884
rect 13580 15986 13636 15988
rect 13580 15934 13582 15986
rect 13582 15934 13634 15986
rect 13634 15934 13636 15986
rect 13580 15932 13636 15934
rect 14364 16322 14420 16324
rect 14364 16270 14366 16322
rect 14366 16270 14418 16322
rect 14418 16270 14420 16322
rect 14364 16268 14420 16270
rect 14588 15148 14644 15204
rect 13244 13692 13300 13748
rect 13020 13244 13076 13300
rect 12908 12850 12964 12852
rect 12908 12798 12910 12850
rect 12910 12798 12962 12850
rect 12962 12798 12964 12850
rect 12908 12796 12964 12798
rect 13692 12962 13748 12964
rect 13692 12910 13694 12962
rect 13694 12910 13746 12962
rect 13746 12910 13748 12962
rect 13692 12908 13748 12910
rect 13468 12236 13524 12292
rect 12908 11676 12964 11732
rect 13916 13244 13972 13300
rect 14252 12962 14308 12964
rect 14252 12910 14254 12962
rect 14254 12910 14306 12962
rect 14306 12910 14308 12962
rect 14252 12908 14308 12910
rect 14028 12796 14084 12852
rect 13804 11340 13860 11396
rect 13468 10780 13524 10836
rect 13132 10386 13188 10388
rect 13132 10334 13134 10386
rect 13134 10334 13186 10386
rect 13186 10334 13188 10386
rect 13132 10332 13188 10334
rect 13468 9996 13524 10052
rect 12572 9714 12628 9716
rect 12572 9662 12574 9714
rect 12574 9662 12626 9714
rect 12626 9662 12628 9714
rect 12572 9660 12628 9662
rect 13916 11004 13972 11060
rect 13916 10610 13972 10612
rect 13916 10558 13918 10610
rect 13918 10558 13970 10610
rect 13970 10558 13972 10610
rect 13916 10556 13972 10558
rect 15036 18060 15092 18116
rect 14924 13916 14980 13972
rect 15260 20130 15316 20132
rect 15260 20078 15262 20130
rect 15262 20078 15314 20130
rect 15314 20078 15316 20130
rect 15260 20076 15316 20078
rect 15372 18956 15428 19012
rect 15708 23436 15764 23492
rect 15596 23154 15652 23156
rect 15596 23102 15598 23154
rect 15598 23102 15650 23154
rect 15650 23102 15652 23154
rect 15596 23100 15652 23102
rect 16492 29650 16548 29652
rect 16492 29598 16494 29650
rect 16494 29598 16546 29650
rect 16546 29598 16548 29650
rect 16492 29596 16548 29598
rect 16716 29484 16772 29540
rect 16828 28530 16884 28532
rect 16828 28478 16830 28530
rect 16830 28478 16882 28530
rect 16882 28478 16884 28530
rect 16828 28476 16884 28478
rect 16492 27804 16548 27860
rect 19404 39618 19460 39620
rect 19404 39566 19406 39618
rect 19406 39566 19458 39618
rect 19458 39566 19460 39618
rect 19404 39564 19460 39566
rect 21980 42754 22036 42756
rect 21980 42702 21982 42754
rect 21982 42702 22034 42754
rect 22034 42702 22036 42754
rect 21980 42700 22036 42702
rect 20412 42530 20468 42532
rect 20412 42478 20414 42530
rect 20414 42478 20466 42530
rect 20466 42478 20468 42530
rect 20412 42476 20468 42478
rect 20748 41020 20804 41076
rect 20636 40348 20692 40404
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19068 38220 19124 38276
rect 19180 38108 19236 38164
rect 18844 37996 18900 38052
rect 20188 38162 20244 38164
rect 20188 38110 20190 38162
rect 20190 38110 20242 38162
rect 20242 38110 20244 38162
rect 20188 38108 20244 38110
rect 21308 40572 21364 40628
rect 20972 38946 21028 38948
rect 20972 38894 20974 38946
rect 20974 38894 21026 38946
rect 21026 38894 21028 38946
rect 20972 38892 21028 38894
rect 21644 40348 21700 40404
rect 21756 39340 21812 39396
rect 19852 37826 19908 37828
rect 19852 37774 19854 37826
rect 19854 37774 19906 37826
rect 19906 37774 19908 37826
rect 19852 37772 19908 37774
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19628 36988 19684 37044
rect 20412 37324 20468 37380
rect 19740 36428 19796 36484
rect 19516 36316 19572 36372
rect 20076 37100 20132 37156
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 22092 42028 22148 42084
rect 22092 39730 22148 39732
rect 22092 39678 22094 39730
rect 22094 39678 22146 39730
rect 22146 39678 22148 39730
rect 22092 39676 22148 39678
rect 25340 43538 25396 43540
rect 25340 43486 25342 43538
rect 25342 43486 25394 43538
rect 25394 43486 25396 43538
rect 25340 43484 25396 43486
rect 22428 42028 22484 42084
rect 22204 39340 22260 39396
rect 23324 42588 23380 42644
rect 23436 42028 23492 42084
rect 25564 42028 25620 42084
rect 25676 42476 25732 42532
rect 24108 41916 24164 41972
rect 22876 41074 22932 41076
rect 22876 41022 22878 41074
rect 22878 41022 22930 41074
rect 22930 41022 22932 41074
rect 22876 41020 22932 41022
rect 26124 42700 26180 42756
rect 25788 41916 25844 41972
rect 26460 41970 26516 41972
rect 26460 41918 26462 41970
rect 26462 41918 26514 41970
rect 26514 41918 26516 41970
rect 26460 41916 26516 41918
rect 23996 40908 24052 40964
rect 22764 40460 22820 40516
rect 23884 40402 23940 40404
rect 23884 40350 23886 40402
rect 23886 40350 23938 40402
rect 23938 40350 23940 40402
rect 23884 40348 23940 40350
rect 22204 38834 22260 38836
rect 22204 38782 22206 38834
rect 22206 38782 22258 38834
rect 22258 38782 22260 38834
rect 22204 38780 22260 38782
rect 21308 37938 21364 37940
rect 21308 37886 21310 37938
rect 21310 37886 21362 37938
rect 21362 37886 21364 37938
rect 21308 37884 21364 37886
rect 22428 38220 22484 38276
rect 21644 37826 21700 37828
rect 21644 37774 21646 37826
rect 21646 37774 21698 37826
rect 21698 37774 21700 37826
rect 21644 37772 21700 37774
rect 21644 37436 21700 37492
rect 21084 37100 21140 37156
rect 21308 36988 21364 37044
rect 21644 36482 21700 36484
rect 21644 36430 21646 36482
rect 21646 36430 21698 36482
rect 21698 36430 21700 36482
rect 21644 36428 21700 36430
rect 21868 36316 21924 36372
rect 18284 35474 18340 35476
rect 18284 35422 18286 35474
rect 18286 35422 18338 35474
rect 18338 35422 18340 35474
rect 18284 35420 18340 35422
rect 17500 34076 17556 34132
rect 18172 34076 18228 34132
rect 17612 33628 17668 33684
rect 17276 33346 17332 33348
rect 17276 33294 17278 33346
rect 17278 33294 17330 33346
rect 17330 33294 17332 33346
rect 17276 33292 17332 33294
rect 17276 32172 17332 32228
rect 17612 31778 17668 31780
rect 17612 31726 17614 31778
rect 17614 31726 17666 31778
rect 17666 31726 17668 31778
rect 17612 31724 17668 31726
rect 18732 31948 18788 32004
rect 17948 31612 18004 31668
rect 17612 30882 17668 30884
rect 17612 30830 17614 30882
rect 17614 30830 17666 30882
rect 17666 30830 17668 30882
rect 17612 30828 17668 30830
rect 17388 30156 17444 30212
rect 17052 27692 17108 27748
rect 16604 27634 16660 27636
rect 16604 27582 16606 27634
rect 16606 27582 16658 27634
rect 16658 27582 16660 27634
rect 16604 27580 16660 27582
rect 16492 27186 16548 27188
rect 16492 27134 16494 27186
rect 16494 27134 16546 27186
rect 16546 27134 16548 27186
rect 16492 27132 16548 27134
rect 17052 26962 17108 26964
rect 17052 26910 17054 26962
rect 17054 26910 17106 26962
rect 17106 26910 17108 26962
rect 17052 26908 17108 26910
rect 16940 26796 16996 26852
rect 16716 24108 16772 24164
rect 17836 29986 17892 29988
rect 17836 29934 17838 29986
rect 17838 29934 17890 29986
rect 17890 29934 17892 29986
rect 17836 29932 17892 29934
rect 17724 29596 17780 29652
rect 18508 29484 18564 29540
rect 17388 28476 17444 28532
rect 18284 28028 18340 28084
rect 17500 27858 17556 27860
rect 17500 27806 17502 27858
rect 17502 27806 17554 27858
rect 17554 27806 17556 27858
rect 17500 27804 17556 27806
rect 17500 27132 17556 27188
rect 17164 24332 17220 24388
rect 18284 27634 18340 27636
rect 18284 27582 18286 27634
rect 18286 27582 18338 27634
rect 18338 27582 18340 27634
rect 18284 27580 18340 27582
rect 18620 27634 18676 27636
rect 18620 27582 18622 27634
rect 18622 27582 18674 27634
rect 18674 27582 18676 27634
rect 18620 27580 18676 27582
rect 18732 27244 18788 27300
rect 18620 26908 18676 26964
rect 18956 31724 19012 31780
rect 20412 35644 20468 35700
rect 21532 35698 21588 35700
rect 21532 35646 21534 35698
rect 21534 35646 21586 35698
rect 21586 35646 21588 35698
rect 21532 35644 21588 35646
rect 22316 36988 22372 37044
rect 22092 36876 22148 36932
rect 22092 36316 22148 36372
rect 22204 35810 22260 35812
rect 22204 35758 22206 35810
rect 22206 35758 22258 35810
rect 22258 35758 22260 35810
rect 22204 35756 22260 35758
rect 20860 34636 20916 34692
rect 21756 34636 21812 34692
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19292 34076 19348 34132
rect 19292 33852 19348 33908
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20300 32508 20356 32564
rect 19292 32396 19348 32452
rect 19404 31836 19460 31892
rect 17948 26460 18004 26516
rect 18620 26124 18676 26180
rect 18508 26066 18564 26068
rect 18508 26014 18510 26066
rect 18510 26014 18562 26066
rect 18562 26014 18564 26066
rect 18508 26012 18564 26014
rect 17612 25900 17668 25956
rect 17724 25394 17780 25396
rect 17724 25342 17726 25394
rect 17726 25342 17778 25394
rect 17778 25342 17780 25394
rect 17724 25340 17780 25342
rect 15708 22764 15764 22820
rect 15708 22482 15764 22484
rect 15708 22430 15710 22482
rect 15710 22430 15762 22482
rect 15762 22430 15764 22482
rect 15708 22428 15764 22430
rect 16604 22988 16660 23044
rect 16492 22428 16548 22484
rect 15708 21980 15764 22036
rect 16044 21980 16100 22036
rect 16156 21586 16212 21588
rect 16156 21534 16158 21586
rect 16158 21534 16210 21586
rect 16210 21534 16212 21586
rect 16156 21532 16212 21534
rect 17164 21868 17220 21924
rect 16492 21644 16548 21700
rect 16828 21698 16884 21700
rect 16828 21646 16830 21698
rect 16830 21646 16882 21698
rect 16882 21646 16884 21698
rect 16828 21644 16884 21646
rect 16044 20690 16100 20692
rect 16044 20638 16046 20690
rect 16046 20638 16098 20690
rect 16098 20638 16100 20690
rect 16044 20636 16100 20638
rect 15708 19740 15764 19796
rect 15932 20524 15988 20580
rect 15708 19292 15764 19348
rect 15596 18732 15652 18788
rect 15932 18844 15988 18900
rect 15484 18620 15540 18676
rect 15484 18172 15540 18228
rect 15708 18284 15764 18340
rect 15372 17612 15428 17668
rect 15932 17388 15988 17444
rect 17836 22316 17892 22372
rect 18172 23660 18228 23716
rect 18620 24722 18676 24724
rect 18620 24670 18622 24722
rect 18622 24670 18674 24722
rect 18674 24670 18676 24722
rect 18620 24668 18676 24670
rect 18620 24108 18676 24164
rect 18508 23212 18564 23268
rect 17948 23100 18004 23156
rect 18172 21980 18228 22036
rect 18396 22204 18452 22260
rect 17836 21756 17892 21812
rect 17500 21586 17556 21588
rect 17500 21534 17502 21586
rect 17502 21534 17554 21586
rect 17554 21534 17556 21586
rect 17500 21532 17556 21534
rect 17388 21308 17444 21364
rect 16828 20860 16884 20916
rect 16716 20018 16772 20020
rect 16716 19966 16718 20018
rect 16718 19966 16770 20018
rect 16770 19966 16772 20018
rect 16716 19964 16772 19966
rect 16716 19740 16772 19796
rect 16380 18956 16436 19012
rect 16380 18620 16436 18676
rect 16716 19122 16772 19124
rect 16716 19070 16718 19122
rect 16718 19070 16770 19122
rect 16770 19070 16772 19122
rect 16716 19068 16772 19070
rect 16828 18956 16884 19012
rect 17164 20802 17220 20804
rect 17164 20750 17166 20802
rect 17166 20750 17218 20802
rect 17218 20750 17220 20802
rect 17164 20748 17220 20750
rect 18396 21532 18452 21588
rect 18060 21308 18116 21364
rect 18284 21420 18340 21476
rect 17276 20690 17332 20692
rect 17276 20638 17278 20690
rect 17278 20638 17330 20690
rect 17330 20638 17332 20690
rect 17276 20636 17332 20638
rect 17388 20578 17444 20580
rect 17388 20526 17390 20578
rect 17390 20526 17442 20578
rect 17442 20526 17444 20578
rect 17388 20524 17444 20526
rect 17388 20130 17444 20132
rect 17388 20078 17390 20130
rect 17390 20078 17442 20130
rect 17442 20078 17444 20130
rect 17388 20076 17444 20078
rect 17612 19404 17668 19460
rect 17948 19122 18004 19124
rect 17948 19070 17950 19122
rect 17950 19070 18002 19122
rect 18002 19070 18004 19122
rect 17948 19068 18004 19070
rect 18172 19740 18228 19796
rect 18060 18732 18116 18788
rect 16604 17724 16660 17780
rect 17836 18508 17892 18564
rect 16268 17052 16324 17108
rect 16828 18172 16884 18228
rect 17612 18284 17668 18340
rect 16380 16882 16436 16884
rect 16380 16830 16382 16882
rect 16382 16830 16434 16882
rect 16434 16830 16436 16882
rect 16380 16828 16436 16830
rect 17388 17442 17444 17444
rect 17388 17390 17390 17442
rect 17390 17390 17442 17442
rect 17442 17390 17444 17442
rect 17388 17388 17444 17390
rect 15932 16604 15988 16660
rect 16604 16604 16660 16660
rect 18172 18450 18228 18452
rect 18172 18398 18174 18450
rect 18174 18398 18226 18450
rect 18226 18398 18228 18450
rect 18172 18396 18228 18398
rect 17948 18172 18004 18228
rect 17836 18060 17892 18116
rect 18060 17106 18116 17108
rect 18060 17054 18062 17106
rect 18062 17054 18114 17106
rect 18114 17054 18116 17106
rect 18060 17052 18116 17054
rect 17724 16604 17780 16660
rect 17388 16044 17444 16100
rect 17500 16156 17556 16212
rect 16268 15484 16324 15540
rect 16828 15538 16884 15540
rect 16828 15486 16830 15538
rect 16830 15486 16882 15538
rect 16882 15486 16884 15538
rect 16828 15484 16884 15486
rect 17500 15484 17556 15540
rect 15260 15372 15316 15428
rect 18172 15820 18228 15876
rect 16828 14700 16884 14756
rect 18620 19628 18676 19684
rect 18508 19292 18564 19348
rect 18508 18562 18564 18564
rect 18508 18510 18510 18562
rect 18510 18510 18562 18562
rect 18562 18510 18564 18562
rect 18508 18508 18564 18510
rect 18396 17500 18452 17556
rect 18844 25116 18900 25172
rect 19852 31778 19908 31780
rect 19852 31726 19854 31778
rect 19854 31726 19906 31778
rect 19906 31726 19908 31778
rect 19852 31724 19908 31726
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20412 32450 20468 32452
rect 20412 32398 20414 32450
rect 20414 32398 20466 32450
rect 20466 32398 20468 32450
rect 20412 32396 20468 32398
rect 20412 32172 20468 32228
rect 21644 33292 21700 33348
rect 21420 33180 21476 33236
rect 21420 32562 21476 32564
rect 21420 32510 21422 32562
rect 21422 32510 21474 32562
rect 21474 32510 21476 32562
rect 21420 32508 21476 32510
rect 21196 32060 21252 32116
rect 20972 31948 21028 32004
rect 20748 31164 20804 31220
rect 19516 30210 19572 30212
rect 19516 30158 19518 30210
rect 19518 30158 19570 30210
rect 19570 30158 19572 30210
rect 19516 30156 19572 30158
rect 19180 27804 19236 27860
rect 19628 29932 19684 29988
rect 20188 30156 20244 30212
rect 19404 29260 19460 29316
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20300 29708 20356 29764
rect 19964 28418 20020 28420
rect 19964 28366 19966 28418
rect 19966 28366 20018 28418
rect 20018 28366 20020 28418
rect 19964 28364 20020 28366
rect 20188 29260 20244 29316
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19516 27356 19572 27412
rect 19404 27074 19460 27076
rect 19404 27022 19406 27074
rect 19406 27022 19458 27074
rect 19458 27022 19460 27074
rect 19404 27020 19460 27022
rect 19292 26684 19348 26740
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20860 29426 20916 29428
rect 20860 29374 20862 29426
rect 20862 29374 20914 29426
rect 20914 29374 20916 29426
rect 20860 29372 20916 29374
rect 20860 28364 20916 28420
rect 20524 27074 20580 27076
rect 20524 27022 20526 27074
rect 20526 27022 20578 27074
rect 20578 27022 20580 27074
rect 20524 27020 20580 27022
rect 20748 28028 20804 28084
rect 18956 18844 19012 18900
rect 19852 25506 19908 25508
rect 19852 25454 19854 25506
rect 19854 25454 19906 25506
rect 19906 25454 19908 25506
rect 19852 25452 19908 25454
rect 19404 25116 19460 25172
rect 18284 14588 18340 14644
rect 18732 17500 18788 17556
rect 14812 13746 14868 13748
rect 14812 13694 14814 13746
rect 14814 13694 14866 13746
rect 14866 13694 14868 13746
rect 14812 13692 14868 13694
rect 14924 13020 14980 13076
rect 15148 12908 15204 12964
rect 14476 12012 14532 12068
rect 14364 11900 14420 11956
rect 14028 10050 14084 10052
rect 14028 9998 14030 10050
rect 14030 9998 14082 10050
rect 14082 9998 14084 10050
rect 14028 9996 14084 9998
rect 14140 11004 14196 11060
rect 15036 11900 15092 11956
rect 14700 11004 14756 11060
rect 15820 13132 15876 13188
rect 16940 13186 16996 13188
rect 16940 13134 16942 13186
rect 16942 13134 16994 13186
rect 16994 13134 16996 13186
rect 16940 13132 16996 13134
rect 16492 13020 16548 13076
rect 16380 12908 16436 12964
rect 15484 12796 15540 12852
rect 15260 11900 15316 11956
rect 15372 12066 15428 12068
rect 15372 12014 15374 12066
rect 15374 12014 15426 12066
rect 15426 12014 15428 12066
rect 15372 12012 15428 12014
rect 14924 10556 14980 10612
rect 14476 8930 14532 8932
rect 14476 8878 14478 8930
rect 14478 8878 14530 8930
rect 14530 8878 14532 8930
rect 14476 8876 14532 8878
rect 14252 8204 14308 8260
rect 15036 8258 15092 8260
rect 15036 8206 15038 8258
rect 15038 8206 15090 8258
rect 15090 8206 15092 8258
rect 15036 8204 15092 8206
rect 5852 6860 5908 6916
rect 15484 11788 15540 11844
rect 16380 11788 16436 11844
rect 15708 11340 15764 11396
rect 17276 12738 17332 12740
rect 17276 12686 17278 12738
rect 17278 12686 17330 12738
rect 17330 12686 17332 12738
rect 17276 12684 17332 12686
rect 17052 12236 17108 12292
rect 16828 11394 16884 11396
rect 16828 11342 16830 11394
rect 16830 11342 16882 11394
rect 16882 11342 16884 11394
rect 16828 11340 16884 11342
rect 18732 17052 18788 17108
rect 18732 16492 18788 16548
rect 18620 15986 18676 15988
rect 18620 15934 18622 15986
rect 18622 15934 18674 15986
rect 18674 15934 18676 15986
rect 18620 15932 18676 15934
rect 17612 13916 17668 13972
rect 17612 13356 17668 13412
rect 17836 13916 17892 13972
rect 19292 24050 19348 24052
rect 19292 23998 19294 24050
rect 19294 23998 19346 24050
rect 19346 23998 19348 24050
rect 19292 23996 19348 23998
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 21644 32172 21700 32228
rect 21980 34690 22036 34692
rect 21980 34638 21982 34690
rect 21982 34638 22034 34690
rect 22034 34638 22036 34690
rect 21980 34636 22036 34638
rect 22092 34524 22148 34580
rect 22204 35196 22260 35252
rect 21868 33628 21924 33684
rect 22428 36316 22484 36372
rect 22988 38050 23044 38052
rect 22988 37998 22990 38050
rect 22990 37998 23042 38050
rect 23042 37998 23044 38050
rect 22988 37996 23044 37998
rect 22764 36876 22820 36932
rect 22540 36204 22596 36260
rect 22652 34972 22708 35028
rect 22876 36204 22932 36260
rect 22876 35420 22932 35476
rect 22876 35196 22932 35252
rect 23772 38220 23828 38276
rect 25564 41356 25620 41412
rect 25452 40348 25508 40404
rect 24108 38668 24164 38724
rect 25452 38668 25508 38724
rect 24556 38220 24612 38276
rect 23436 37772 23492 37828
rect 22428 34242 22484 34244
rect 22428 34190 22430 34242
rect 22430 34190 22482 34242
rect 22482 34190 22484 34242
rect 22428 34188 22484 34190
rect 23212 34524 23268 34580
rect 23548 36988 23604 37044
rect 23548 35756 23604 35812
rect 23212 33852 23268 33908
rect 22652 33628 22708 33684
rect 21756 31778 21812 31780
rect 21756 31726 21758 31778
rect 21758 31726 21810 31778
rect 21810 31726 21812 31778
rect 21756 31724 21812 31726
rect 21644 31612 21700 31668
rect 22428 33346 22484 33348
rect 22428 33294 22430 33346
rect 22430 33294 22482 33346
rect 22482 33294 22484 33346
rect 22428 33292 22484 33294
rect 22204 33234 22260 33236
rect 22204 33182 22206 33234
rect 22206 33182 22258 33234
rect 22258 33182 22260 33234
rect 22204 33180 22260 33182
rect 22204 32674 22260 32676
rect 22204 32622 22206 32674
rect 22206 32622 22258 32674
rect 22258 32622 22260 32674
rect 22204 32620 22260 32622
rect 22204 32284 22260 32340
rect 22092 31836 22148 31892
rect 21756 29986 21812 29988
rect 21756 29934 21758 29986
rect 21758 29934 21810 29986
rect 21810 29934 21812 29986
rect 21756 29932 21812 29934
rect 21196 29708 21252 29764
rect 21308 28530 21364 28532
rect 21308 28478 21310 28530
rect 21310 28478 21362 28530
rect 21362 28478 21364 28530
rect 21308 28476 21364 28478
rect 21420 28418 21476 28420
rect 21420 28366 21422 28418
rect 21422 28366 21474 28418
rect 21474 28366 21476 28418
rect 21420 28364 21476 28366
rect 20972 26460 21028 26516
rect 20972 26012 21028 26068
rect 20188 25004 20244 25060
rect 19740 24892 19796 24948
rect 20412 24892 20468 24948
rect 19404 23884 19460 23940
rect 19292 23660 19348 23716
rect 19292 22092 19348 22148
rect 19516 21756 19572 21812
rect 20188 24834 20244 24836
rect 20188 24782 20190 24834
rect 20190 24782 20242 24834
rect 20242 24782 20244 24834
rect 20188 24780 20244 24782
rect 20188 23938 20244 23940
rect 20188 23886 20190 23938
rect 20190 23886 20242 23938
rect 20242 23886 20244 23938
rect 20188 23884 20244 23886
rect 19740 23660 19796 23716
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20300 23212 20356 23268
rect 19964 22370 20020 22372
rect 19964 22318 19966 22370
rect 19966 22318 20018 22370
rect 20018 22318 20020 22370
rect 19964 22316 20020 22318
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20524 22482 20580 22484
rect 20524 22430 20526 22482
rect 20526 22430 20578 22482
rect 20578 22430 20580 22482
rect 20524 22428 20580 22430
rect 21308 27804 21364 27860
rect 21980 30604 22036 30660
rect 22092 30210 22148 30212
rect 22092 30158 22094 30210
rect 22094 30158 22146 30210
rect 22146 30158 22148 30210
rect 22092 30156 22148 30158
rect 22764 33122 22820 33124
rect 22764 33070 22766 33122
rect 22766 33070 22818 33122
rect 22818 33070 22820 33122
rect 22764 33068 22820 33070
rect 22540 31164 22596 31220
rect 22428 30604 22484 30660
rect 22540 29932 22596 29988
rect 23100 29820 23156 29876
rect 23324 33068 23380 33124
rect 23436 31724 23492 31780
rect 22316 29260 22372 29316
rect 22652 29372 22708 29428
rect 21980 29036 22036 29092
rect 21644 27804 21700 27860
rect 21532 27356 21588 27412
rect 21308 26012 21364 26068
rect 21308 25340 21364 25396
rect 21308 24220 21364 24276
rect 20748 23378 20804 23380
rect 20748 23326 20750 23378
rect 20750 23326 20802 23378
rect 20802 23326 20804 23378
rect 20748 23324 20804 23326
rect 21756 27244 21812 27300
rect 22316 28588 22372 28644
rect 22092 28418 22148 28420
rect 22092 28366 22094 28418
rect 22094 28366 22146 28418
rect 22146 28366 22148 28418
rect 22092 28364 22148 28366
rect 21980 27804 22036 27860
rect 22204 27580 22260 27636
rect 22092 27132 22148 27188
rect 22428 27020 22484 27076
rect 21980 26796 22036 26852
rect 21980 26402 22036 26404
rect 21980 26350 21982 26402
rect 21982 26350 22034 26402
rect 22034 26350 22036 26402
rect 21980 26348 22036 26350
rect 21756 26290 21812 26292
rect 21756 26238 21758 26290
rect 21758 26238 21810 26290
rect 21810 26238 21812 26290
rect 21756 26236 21812 26238
rect 21644 25900 21700 25956
rect 21644 25452 21700 25508
rect 21420 23154 21476 23156
rect 21420 23102 21422 23154
rect 21422 23102 21474 23154
rect 21474 23102 21476 23154
rect 21420 23100 21476 23102
rect 21420 22652 21476 22708
rect 20636 22316 20692 22372
rect 20412 21810 20468 21812
rect 20412 21758 20414 21810
rect 20414 21758 20466 21810
rect 20466 21758 20468 21810
rect 20412 21756 20468 21758
rect 20636 21756 20692 21812
rect 20300 21084 20356 21140
rect 19628 20860 19684 20916
rect 20300 20914 20356 20916
rect 20300 20862 20302 20914
rect 20302 20862 20354 20914
rect 20354 20862 20356 20914
rect 20300 20860 20356 20862
rect 20972 21644 21028 21700
rect 20860 21196 20916 21252
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20076 20076 20132 20132
rect 19628 19516 19684 19572
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19740 18508 19796 18564
rect 19180 16716 19236 16772
rect 19292 18284 19348 18340
rect 19068 16492 19124 16548
rect 19404 17500 19460 17556
rect 21420 22370 21476 22372
rect 21420 22318 21422 22370
rect 21422 22318 21474 22370
rect 21474 22318 21476 22370
rect 21420 22316 21476 22318
rect 21084 20076 21140 20132
rect 21532 21756 21588 21812
rect 22428 26012 22484 26068
rect 22316 25506 22372 25508
rect 22316 25454 22318 25506
rect 22318 25454 22370 25506
rect 22370 25454 22372 25506
rect 22316 25452 22372 25454
rect 22988 29148 23044 29204
rect 23100 29260 23156 29316
rect 23436 29372 23492 29428
rect 23436 29148 23492 29204
rect 23324 28588 23380 28644
rect 23212 28028 23268 28084
rect 23436 28418 23492 28420
rect 23436 28366 23438 28418
rect 23438 28366 23490 28418
rect 23490 28366 23492 28418
rect 23436 28364 23492 28366
rect 23100 27074 23156 27076
rect 23100 27022 23102 27074
rect 23102 27022 23154 27074
rect 23154 27022 23156 27074
rect 23100 27020 23156 27022
rect 23996 37884 24052 37940
rect 23996 37266 24052 37268
rect 23996 37214 23998 37266
rect 23998 37214 24050 37266
rect 24050 37214 24052 37266
rect 23996 37212 24052 37214
rect 24220 37826 24276 37828
rect 24220 37774 24222 37826
rect 24222 37774 24274 37826
rect 24274 37774 24276 37826
rect 24220 37772 24276 37774
rect 24556 37826 24612 37828
rect 24556 37774 24558 37826
rect 24558 37774 24610 37826
rect 24610 37774 24612 37826
rect 24556 37772 24612 37774
rect 24444 37100 24500 37156
rect 24108 36652 24164 36708
rect 24556 36988 24612 37044
rect 25228 37826 25284 37828
rect 25228 37774 25230 37826
rect 25230 37774 25282 37826
rect 25282 37774 25284 37826
rect 25228 37772 25284 37774
rect 25452 37212 25508 37268
rect 24892 36428 24948 36484
rect 25340 37154 25396 37156
rect 25340 37102 25342 37154
rect 25342 37102 25394 37154
rect 25394 37102 25396 37154
rect 25340 37100 25396 37102
rect 26236 38220 26292 38276
rect 25900 37884 25956 37940
rect 25788 37490 25844 37492
rect 25788 37438 25790 37490
rect 25790 37438 25842 37490
rect 25842 37438 25844 37490
rect 25788 37436 25844 37438
rect 25676 36540 25732 36596
rect 24332 35420 24388 35476
rect 25564 35474 25620 35476
rect 25564 35422 25566 35474
rect 25566 35422 25618 35474
rect 25618 35422 25620 35474
rect 25564 35420 25620 35422
rect 23772 34636 23828 34692
rect 23660 34188 23716 34244
rect 26124 37660 26180 37716
rect 26908 42028 26964 42084
rect 28028 42476 28084 42532
rect 27244 41356 27300 41412
rect 27132 41132 27188 41188
rect 27132 40460 27188 40516
rect 27356 39676 27412 39732
rect 26572 37772 26628 37828
rect 26460 37266 26516 37268
rect 26460 37214 26462 37266
rect 26462 37214 26514 37266
rect 26514 37214 26516 37266
rect 26460 37212 26516 37214
rect 26348 36876 26404 36932
rect 26348 34972 26404 35028
rect 25228 34242 25284 34244
rect 25228 34190 25230 34242
rect 25230 34190 25282 34242
rect 25282 34190 25284 34242
rect 25228 34188 25284 34190
rect 27132 37100 27188 37156
rect 26684 36204 26740 36260
rect 27580 39564 27636 39620
rect 27692 39506 27748 39508
rect 27692 39454 27694 39506
rect 27694 39454 27746 39506
rect 27746 39454 27748 39506
rect 27692 39452 27748 39454
rect 29484 43538 29540 43540
rect 29484 43486 29486 43538
rect 29486 43486 29538 43538
rect 29538 43486 29540 43538
rect 29484 43484 29540 43486
rect 30492 43484 30548 43540
rect 28364 42700 28420 42756
rect 28252 40572 28308 40628
rect 28364 42476 28420 42532
rect 28028 39228 28084 39284
rect 27804 37884 27860 37940
rect 28700 41916 28756 41972
rect 28476 41020 28532 41076
rect 28476 40402 28532 40404
rect 28476 40350 28478 40402
rect 28478 40350 28530 40402
rect 28530 40350 28532 40402
rect 28476 40348 28532 40350
rect 29148 39394 29204 39396
rect 29148 39342 29150 39394
rect 29150 39342 29202 39394
rect 29202 39342 29204 39394
rect 29148 39340 29204 39342
rect 30492 42754 30548 42756
rect 30492 42702 30494 42754
rect 30494 42702 30546 42754
rect 30546 42702 30548 42754
rect 30492 42700 30548 42702
rect 30044 41970 30100 41972
rect 30044 41918 30046 41970
rect 30046 41918 30098 41970
rect 30098 41918 30100 41970
rect 30044 41916 30100 41918
rect 29484 41186 29540 41188
rect 29484 41134 29486 41186
rect 29486 41134 29538 41186
rect 29538 41134 29540 41186
rect 29484 41132 29540 41134
rect 29932 41186 29988 41188
rect 29932 41134 29934 41186
rect 29934 41134 29986 41186
rect 29986 41134 29988 41186
rect 29932 41132 29988 41134
rect 29708 40348 29764 40404
rect 30156 40962 30212 40964
rect 30156 40910 30158 40962
rect 30158 40910 30210 40962
rect 30210 40910 30212 40962
rect 30156 40908 30212 40910
rect 30604 41074 30660 41076
rect 30604 41022 30606 41074
rect 30606 41022 30658 41074
rect 30658 41022 30660 41074
rect 30604 41020 30660 41022
rect 30492 40460 30548 40516
rect 29708 39564 29764 39620
rect 30044 39618 30100 39620
rect 30044 39566 30046 39618
rect 30046 39566 30098 39618
rect 30098 39566 30100 39618
rect 30044 39564 30100 39566
rect 29372 39506 29428 39508
rect 29372 39454 29374 39506
rect 29374 39454 29426 39506
rect 29426 39454 29428 39506
rect 29372 39452 29428 39454
rect 30716 38892 30772 38948
rect 30044 38668 30100 38724
rect 27020 35420 27076 35476
rect 26572 35026 26628 35028
rect 26572 34974 26574 35026
rect 26574 34974 26626 35026
rect 26626 34974 26628 35026
rect 26572 34972 26628 34974
rect 26348 33852 26404 33908
rect 24444 33628 24500 33684
rect 25564 33516 25620 33572
rect 23996 33404 24052 33460
rect 25228 33346 25284 33348
rect 25228 33294 25230 33346
rect 25230 33294 25282 33346
rect 25282 33294 25284 33346
rect 25228 33292 25284 33294
rect 24556 33068 24612 33124
rect 25452 33122 25508 33124
rect 25452 33070 25454 33122
rect 25454 33070 25506 33122
rect 25506 33070 25508 33122
rect 25452 33068 25508 33070
rect 24444 32508 24500 32564
rect 23884 29708 23940 29764
rect 24108 31164 24164 31220
rect 24332 30828 24388 30884
rect 24332 29820 24388 29876
rect 23660 29484 23716 29540
rect 23884 28642 23940 28644
rect 23884 28590 23886 28642
rect 23886 28590 23938 28642
rect 23938 28590 23940 28642
rect 23884 28588 23940 28590
rect 23660 27858 23716 27860
rect 23660 27806 23662 27858
rect 23662 27806 23714 27858
rect 23714 27806 23716 27858
rect 23660 27804 23716 27806
rect 23548 26908 23604 26964
rect 22540 25900 22596 25956
rect 22652 25340 22708 25396
rect 22316 24610 22372 24612
rect 22316 24558 22318 24610
rect 22318 24558 22370 24610
rect 22370 24558 22372 24610
rect 22316 24556 22372 24558
rect 21756 23212 21812 23268
rect 22204 23100 22260 23156
rect 22764 25004 22820 25060
rect 22764 23660 22820 23716
rect 21868 22370 21924 22372
rect 21868 22318 21870 22370
rect 21870 22318 21922 22370
rect 21922 22318 21924 22370
rect 21868 22316 21924 22318
rect 22092 21810 22148 21812
rect 22092 21758 22094 21810
rect 22094 21758 22146 21810
rect 22146 21758 22148 21810
rect 22092 21756 22148 21758
rect 21196 18620 21252 18676
rect 21756 19346 21812 19348
rect 21756 19294 21758 19346
rect 21758 19294 21810 19346
rect 21810 19294 21812 19346
rect 21756 19292 21812 19294
rect 20524 18284 20580 18340
rect 20076 17554 20132 17556
rect 20076 17502 20078 17554
rect 20078 17502 20130 17554
rect 20130 17502 20132 17554
rect 20076 17500 20132 17502
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19516 16828 19572 16884
rect 19404 16268 19460 16324
rect 19516 16492 19572 16548
rect 20412 17836 20468 17892
rect 20300 17164 20356 17220
rect 19516 15932 19572 15988
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20300 15538 20356 15540
rect 20300 15486 20302 15538
rect 20302 15486 20354 15538
rect 20354 15486 20356 15538
rect 20300 15484 20356 15486
rect 19628 15148 19684 15204
rect 18732 13970 18788 13972
rect 18732 13918 18734 13970
rect 18734 13918 18786 13970
rect 18786 13918 18788 13970
rect 18732 13916 18788 13918
rect 18284 13356 18340 13412
rect 19964 14924 20020 14980
rect 19740 14252 19796 14308
rect 20188 14252 20244 14308
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 18172 12908 18228 12964
rect 17948 12684 18004 12740
rect 16716 10780 16772 10836
rect 16044 10610 16100 10612
rect 16044 10558 16046 10610
rect 16046 10558 16098 10610
rect 16098 10558 16100 10610
rect 16044 10556 16100 10558
rect 17388 10610 17444 10612
rect 17388 10558 17390 10610
rect 17390 10558 17442 10610
rect 17442 10558 17444 10610
rect 17388 10556 17444 10558
rect 16604 9996 16660 10052
rect 17276 9996 17332 10052
rect 16044 9660 16100 9716
rect 15484 8204 15540 8260
rect 16828 9548 16884 9604
rect 17724 11788 17780 11844
rect 17612 9660 17668 9716
rect 17948 12348 18004 12404
rect 17948 11788 18004 11844
rect 18172 12402 18228 12404
rect 18172 12350 18174 12402
rect 18174 12350 18226 12402
rect 18226 12350 18228 12402
rect 18172 12348 18228 12350
rect 18172 11900 18228 11956
rect 17500 9548 17556 9604
rect 16156 9100 16212 9156
rect 16380 8428 16436 8484
rect 16156 8316 16212 8372
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 18172 10498 18228 10500
rect 18172 10446 18174 10498
rect 18174 10446 18226 10498
rect 18226 10446 18228 10498
rect 18172 10444 18228 10446
rect 18396 11788 18452 11844
rect 19292 12290 19348 12292
rect 19292 12238 19294 12290
rect 19294 12238 19346 12290
rect 19346 12238 19348 12290
rect 19292 12236 19348 12238
rect 19516 12236 19572 12292
rect 18508 10498 18564 10500
rect 18508 10446 18510 10498
rect 18510 10446 18562 10498
rect 18562 10446 18564 10498
rect 18508 10444 18564 10446
rect 18172 9548 18228 9604
rect 18620 9154 18676 9156
rect 18620 9102 18622 9154
rect 18622 9102 18674 9154
rect 18674 9102 18676 9154
rect 18620 9100 18676 9102
rect 17836 8428 17892 8484
rect 19852 13916 19908 13972
rect 19852 12962 19908 12964
rect 19852 12910 19854 12962
rect 19854 12910 19906 12962
rect 19906 12910 19908 12962
rect 19852 12908 19908 12910
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19852 12348 19908 12404
rect 19740 12290 19796 12292
rect 19740 12238 19742 12290
rect 19742 12238 19794 12290
rect 19794 12238 19796 12290
rect 19740 12236 19796 12238
rect 19628 11564 19684 11620
rect 21532 17276 21588 17332
rect 21644 16716 21700 16772
rect 20524 16268 20580 16324
rect 20524 15874 20580 15876
rect 20524 15822 20526 15874
rect 20526 15822 20578 15874
rect 20578 15822 20580 15874
rect 20524 15820 20580 15822
rect 20748 15202 20804 15204
rect 20748 15150 20750 15202
rect 20750 15150 20802 15202
rect 20802 15150 20804 15202
rect 20748 15148 20804 15150
rect 21420 16380 21476 16436
rect 21644 16492 21700 16548
rect 22316 21810 22372 21812
rect 22316 21758 22318 21810
rect 22318 21758 22370 21810
rect 22370 21758 22372 21810
rect 22316 21756 22372 21758
rect 22092 21420 22148 21476
rect 23100 26236 23156 26292
rect 22988 23436 23044 23492
rect 22876 22876 22932 22932
rect 23548 26290 23604 26292
rect 23548 26238 23550 26290
rect 23550 26238 23602 26290
rect 23602 26238 23604 26290
rect 23548 26236 23604 26238
rect 23436 25394 23492 25396
rect 23436 25342 23438 25394
rect 23438 25342 23490 25394
rect 23490 25342 23492 25394
rect 23436 25340 23492 25342
rect 23772 25506 23828 25508
rect 23772 25454 23774 25506
rect 23774 25454 23826 25506
rect 23826 25454 23828 25506
rect 23772 25452 23828 25454
rect 23660 25116 23716 25172
rect 24220 28476 24276 28532
rect 23996 28082 24052 28084
rect 23996 28030 23998 28082
rect 23998 28030 24050 28082
rect 24050 28030 24052 28082
rect 23996 28028 24052 28030
rect 25340 32060 25396 32116
rect 25676 33404 25732 33460
rect 25564 32396 25620 32452
rect 25228 31778 25284 31780
rect 25228 31726 25230 31778
rect 25230 31726 25282 31778
rect 25282 31726 25284 31778
rect 25228 31724 25284 31726
rect 25228 30882 25284 30884
rect 25228 30830 25230 30882
rect 25230 30830 25282 30882
rect 25282 30830 25284 30882
rect 25228 30828 25284 30830
rect 26572 33180 26628 33236
rect 26348 33068 26404 33124
rect 25900 32562 25956 32564
rect 25900 32510 25902 32562
rect 25902 32510 25954 32562
rect 25954 32510 25956 32562
rect 25900 32508 25956 32510
rect 27132 35196 27188 35252
rect 27692 36652 27748 36708
rect 29260 38556 29316 38612
rect 27804 35980 27860 36036
rect 27580 35308 27636 35364
rect 28252 35308 28308 35364
rect 28476 36316 28532 36372
rect 28588 35980 28644 36036
rect 28028 33740 28084 33796
rect 28588 33404 28644 33460
rect 28252 33234 28308 33236
rect 28252 33182 28254 33234
rect 28254 33182 28306 33234
rect 28306 33182 28308 33234
rect 28252 33180 28308 33182
rect 28028 32562 28084 32564
rect 28028 32510 28030 32562
rect 28030 32510 28082 32562
rect 28082 32510 28084 32562
rect 28028 32508 28084 32510
rect 28700 33122 28756 33124
rect 28700 33070 28702 33122
rect 28702 33070 28754 33122
rect 28754 33070 28756 33122
rect 28700 33068 28756 33070
rect 27020 32396 27076 32452
rect 27020 31948 27076 32004
rect 25564 31554 25620 31556
rect 25564 31502 25566 31554
rect 25566 31502 25618 31554
rect 25618 31502 25620 31554
rect 25564 31500 25620 31502
rect 25564 31164 25620 31220
rect 24556 30156 24612 30212
rect 25340 30268 25396 30324
rect 24892 29484 24948 29540
rect 24556 29372 24612 29428
rect 25116 28476 25172 28532
rect 24892 28364 24948 28420
rect 24556 28028 24612 28084
rect 24220 27580 24276 27636
rect 24332 27356 24388 27412
rect 23996 27074 24052 27076
rect 23996 27022 23998 27074
rect 23998 27022 24050 27074
rect 24050 27022 24052 27074
rect 23996 27020 24052 27022
rect 24220 26852 24276 26908
rect 23996 26348 24052 26404
rect 24444 26572 24500 26628
rect 24668 27580 24724 27636
rect 25004 27580 25060 27636
rect 24780 26908 24836 26964
rect 24108 26012 24164 26068
rect 23996 25116 24052 25172
rect 23324 24668 23380 24724
rect 23324 23938 23380 23940
rect 23324 23886 23326 23938
rect 23326 23886 23378 23938
rect 23378 23886 23380 23938
rect 23324 23884 23380 23886
rect 23548 23772 23604 23828
rect 23436 23660 23492 23716
rect 23212 22764 23268 22820
rect 23436 22876 23492 22932
rect 23324 22428 23380 22484
rect 22652 21532 22708 21588
rect 22540 21308 22596 21364
rect 23548 22652 23604 22708
rect 23100 22092 23156 22148
rect 23324 21308 23380 21364
rect 22876 20860 22932 20916
rect 22092 20524 22148 20580
rect 22540 19852 22596 19908
rect 22540 18508 22596 18564
rect 22764 19292 22820 19348
rect 23100 18396 23156 18452
rect 22876 17724 22932 17780
rect 21980 17554 22036 17556
rect 21980 17502 21982 17554
rect 21982 17502 22034 17554
rect 22034 17502 22036 17554
rect 21980 17500 22036 17502
rect 21868 16604 21924 16660
rect 21868 16380 21924 16436
rect 21868 16044 21924 16100
rect 21308 14924 21364 14980
rect 20524 13020 20580 13076
rect 20412 12962 20468 12964
rect 20412 12910 20414 12962
rect 20414 12910 20466 12962
rect 20466 12910 20468 12962
rect 20412 12908 20468 12910
rect 21532 12796 21588 12852
rect 20076 11788 20132 11844
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19964 10610 20020 10612
rect 19964 10558 19966 10610
rect 19966 10558 20018 10610
rect 20018 10558 20020 10610
rect 19964 10556 20020 10558
rect 19628 10108 19684 10164
rect 20188 9826 20244 9828
rect 20188 9774 20190 9826
rect 20190 9774 20242 9826
rect 20242 9774 20244 9826
rect 20188 9772 20244 9774
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 17724 8316 17780 8372
rect 18732 8258 18788 8260
rect 18732 8206 18734 8258
rect 18734 8206 18786 8258
rect 18786 8206 18788 8258
rect 18732 8204 18788 8206
rect 18844 7980 18900 8036
rect 18284 6466 18340 6468
rect 18284 6414 18286 6466
rect 18286 6414 18338 6466
rect 18338 6414 18340 6466
rect 18284 6412 18340 6414
rect 18508 6076 18564 6132
rect 1708 4898 1764 4900
rect 1708 4846 1710 4898
rect 1710 4846 1762 4898
rect 1762 4846 1764 4898
rect 1708 4844 1764 4846
rect 16716 4508 16772 4564
rect 18956 6076 19012 6132
rect 18620 5906 18676 5908
rect 18620 5854 18622 5906
rect 18622 5854 18674 5906
rect 18674 5854 18676 5906
rect 18620 5852 18676 5854
rect 19628 8818 19684 8820
rect 19628 8766 19630 8818
rect 19630 8766 19682 8818
rect 19682 8766 19684 8818
rect 19628 8764 19684 8766
rect 19964 8988 20020 9044
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19180 6636 19236 6692
rect 19292 5852 19348 5908
rect 19068 5068 19124 5124
rect 19180 5628 19236 5684
rect 20748 11676 20804 11732
rect 21308 11564 21364 11620
rect 20636 10108 20692 10164
rect 21644 9884 21700 9940
rect 21308 9826 21364 9828
rect 21308 9774 21310 9826
rect 21310 9774 21362 9826
rect 21362 9774 21364 9826
rect 21308 9772 21364 9774
rect 20636 9602 20692 9604
rect 20636 9550 20638 9602
rect 20638 9550 20690 9602
rect 20690 9550 20692 9602
rect 20636 9548 20692 9550
rect 20636 9042 20692 9044
rect 20636 8990 20638 9042
rect 20638 8990 20690 9042
rect 20690 8990 20692 9042
rect 20636 8988 20692 8990
rect 24220 24722 24276 24724
rect 24220 24670 24222 24722
rect 24222 24670 24274 24722
rect 24274 24670 24276 24722
rect 24220 24668 24276 24670
rect 24444 23996 24500 24052
rect 24780 26514 24836 26516
rect 24780 26462 24782 26514
rect 24782 26462 24834 26514
rect 24834 26462 24836 26514
rect 24780 26460 24836 26462
rect 25564 29314 25620 29316
rect 25564 29262 25566 29314
rect 25566 29262 25618 29314
rect 25618 29262 25620 29314
rect 25564 29260 25620 29262
rect 26124 31500 26180 31556
rect 25788 30210 25844 30212
rect 25788 30158 25790 30210
rect 25790 30158 25842 30210
rect 25842 30158 25844 30210
rect 25788 30156 25844 30158
rect 25788 29820 25844 29876
rect 25788 29484 25844 29540
rect 25340 28082 25396 28084
rect 25340 28030 25342 28082
rect 25342 28030 25394 28082
rect 25394 28030 25396 28082
rect 25340 28028 25396 28030
rect 26124 27970 26180 27972
rect 26124 27918 26126 27970
rect 26126 27918 26178 27970
rect 26178 27918 26180 27970
rect 26124 27916 26180 27918
rect 25116 27132 25172 27188
rect 25340 27074 25396 27076
rect 25340 27022 25342 27074
rect 25342 27022 25394 27074
rect 25394 27022 25396 27074
rect 25340 27020 25396 27022
rect 25452 26908 25508 26964
rect 25116 26572 25172 26628
rect 23772 22652 23828 22708
rect 24220 23884 24276 23940
rect 25004 25618 25060 25620
rect 25004 25566 25006 25618
rect 25006 25566 25058 25618
rect 25058 25566 25060 25618
rect 25004 25564 25060 25566
rect 25788 26460 25844 26516
rect 25564 25506 25620 25508
rect 25564 25454 25566 25506
rect 25566 25454 25618 25506
rect 25618 25454 25620 25506
rect 25564 25452 25620 25454
rect 24332 22258 24388 22260
rect 24332 22206 24334 22258
rect 24334 22206 24386 22258
rect 24386 22206 24388 22258
rect 24332 22204 24388 22206
rect 24556 23324 24612 23380
rect 24444 21980 24500 22036
rect 24668 22652 24724 22708
rect 25676 25228 25732 25284
rect 25228 23772 25284 23828
rect 25676 23660 25732 23716
rect 26124 26178 26180 26180
rect 26124 26126 26126 26178
rect 26126 26126 26178 26178
rect 26178 26126 26180 26178
rect 26124 26124 26180 26126
rect 26796 31388 26852 31444
rect 26572 30604 26628 30660
rect 26684 31164 26740 31220
rect 26348 30268 26404 30324
rect 26796 30268 26852 30324
rect 26908 27020 26964 27076
rect 26348 26908 26404 26964
rect 26572 26908 26628 26964
rect 26236 26012 26292 26068
rect 26796 26796 26852 26852
rect 26348 25564 26404 25620
rect 26236 25228 26292 25284
rect 27244 31948 27300 32004
rect 27132 30210 27188 30212
rect 27132 30158 27134 30210
rect 27134 30158 27186 30210
rect 27186 30158 27188 30210
rect 27132 30156 27188 30158
rect 27132 27970 27188 27972
rect 27132 27918 27134 27970
rect 27134 27918 27186 27970
rect 27186 27918 27188 27970
rect 27132 27916 27188 27918
rect 28700 31948 28756 32004
rect 27804 31890 27860 31892
rect 27804 31838 27806 31890
rect 27806 31838 27858 31890
rect 27858 31838 27860 31890
rect 27804 31836 27860 31838
rect 28364 31778 28420 31780
rect 28364 31726 28366 31778
rect 28366 31726 28418 31778
rect 28418 31726 28420 31778
rect 28364 31724 28420 31726
rect 27580 31500 27636 31556
rect 28028 31052 28084 31108
rect 27692 30156 27748 30212
rect 28812 31106 28868 31108
rect 28812 31054 28814 31106
rect 28814 31054 28866 31106
rect 28866 31054 28868 31106
rect 28812 31052 28868 31054
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 31724 42028 31780 42084
rect 46172 42364 46228 42420
rect 33516 42082 33572 42084
rect 33516 42030 33518 42082
rect 33518 42030 33570 42082
rect 33570 42030 33572 42082
rect 33516 42028 33572 42030
rect 32508 41970 32564 41972
rect 32508 41918 32510 41970
rect 32510 41918 32562 41970
rect 32562 41918 32564 41970
rect 32508 41916 32564 41918
rect 33628 41916 33684 41972
rect 31724 41132 31780 41188
rect 31724 40572 31780 40628
rect 31276 40402 31332 40404
rect 31276 40350 31278 40402
rect 31278 40350 31330 40402
rect 31330 40350 31332 40402
rect 31276 40348 31332 40350
rect 30828 38556 30884 38612
rect 32284 39788 32340 39844
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35084 40572 35140 40628
rect 35532 40402 35588 40404
rect 35532 40350 35534 40402
rect 35534 40350 35586 40402
rect 35586 40350 35588 40402
rect 35532 40348 35588 40350
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 34188 39842 34244 39844
rect 34188 39790 34190 39842
rect 34190 39790 34242 39842
rect 34242 39790 34244 39842
rect 34188 39788 34244 39790
rect 33180 39340 33236 39396
rect 33068 39228 33124 39284
rect 32284 38556 32340 38612
rect 31276 37324 31332 37380
rect 29372 36876 29428 36932
rect 29148 36370 29204 36372
rect 29148 36318 29150 36370
rect 29150 36318 29202 36370
rect 29202 36318 29204 36370
rect 29148 36316 29204 36318
rect 29148 35196 29204 35252
rect 30156 36258 30212 36260
rect 30156 36206 30158 36258
rect 30158 36206 30210 36258
rect 30210 36206 30212 36258
rect 30156 36204 30212 36206
rect 30156 35196 30212 35252
rect 29484 33740 29540 33796
rect 29260 33458 29316 33460
rect 29260 33406 29262 33458
rect 29262 33406 29314 33458
rect 29314 33406 29316 33458
rect 29260 33404 29316 33406
rect 29036 33180 29092 33236
rect 29708 33292 29764 33348
rect 29372 33122 29428 33124
rect 29372 33070 29374 33122
rect 29374 33070 29426 33122
rect 29426 33070 29428 33122
rect 29372 33068 29428 33070
rect 29260 31836 29316 31892
rect 29596 31724 29652 31780
rect 30268 31724 30324 31780
rect 29484 31500 29540 31556
rect 29372 31388 29428 31444
rect 28364 30156 28420 30212
rect 29148 30210 29204 30212
rect 29148 30158 29150 30210
rect 29150 30158 29202 30210
rect 29202 30158 29204 30210
rect 29148 30156 29204 30158
rect 28252 29932 28308 29988
rect 27804 29538 27860 29540
rect 27804 29486 27806 29538
rect 27806 29486 27858 29538
rect 27858 29486 27860 29538
rect 27804 29484 27860 29486
rect 28140 28924 28196 28980
rect 27692 28642 27748 28644
rect 27692 28590 27694 28642
rect 27694 28590 27746 28642
rect 27746 28590 27748 28642
rect 27692 28588 27748 28590
rect 28476 29484 28532 29540
rect 28364 28754 28420 28756
rect 28364 28702 28366 28754
rect 28366 28702 28418 28754
rect 28418 28702 28420 28754
rect 28364 28700 28420 28702
rect 29260 29426 29316 29428
rect 29260 29374 29262 29426
rect 29262 29374 29314 29426
rect 29314 29374 29316 29426
rect 29260 29372 29316 29374
rect 28924 28924 28980 28980
rect 27468 26236 27524 26292
rect 28588 27916 28644 27972
rect 28364 26684 28420 26740
rect 28028 26514 28084 26516
rect 28028 26462 28030 26514
rect 28030 26462 28082 26514
rect 28082 26462 28084 26514
rect 28028 26460 28084 26462
rect 28700 27692 28756 27748
rect 28588 27074 28644 27076
rect 28588 27022 28590 27074
rect 28590 27022 28642 27074
rect 28642 27022 28644 27074
rect 28588 27020 28644 27022
rect 28476 26460 28532 26516
rect 28700 26348 28756 26404
rect 28252 26236 28308 26292
rect 27916 25564 27972 25620
rect 27020 25340 27076 25396
rect 26124 24722 26180 24724
rect 26124 24670 26126 24722
rect 26126 24670 26178 24722
rect 26178 24670 26180 24722
rect 26124 24668 26180 24670
rect 26908 25282 26964 25284
rect 26908 25230 26910 25282
rect 26910 25230 26962 25282
rect 26962 25230 26964 25282
rect 26908 25228 26964 25230
rect 27132 25116 27188 25172
rect 26796 24556 26852 24612
rect 26460 24220 26516 24276
rect 26684 23996 26740 24052
rect 26460 23938 26516 23940
rect 26460 23886 26462 23938
rect 26462 23886 26514 23938
rect 26514 23886 26516 23938
rect 26460 23884 26516 23886
rect 26348 23826 26404 23828
rect 26348 23774 26350 23826
rect 26350 23774 26402 23826
rect 26402 23774 26404 23826
rect 26348 23772 26404 23774
rect 27580 25282 27636 25284
rect 27580 25230 27582 25282
rect 27582 25230 27634 25282
rect 27634 25230 27636 25282
rect 27580 25228 27636 25230
rect 27468 25116 27524 25172
rect 27356 24108 27412 24164
rect 28364 26124 28420 26180
rect 29260 28642 29316 28644
rect 29260 28590 29262 28642
rect 29262 28590 29314 28642
rect 29314 28590 29316 28642
rect 29260 28588 29316 28590
rect 30940 37100 30996 37156
rect 30604 36482 30660 36484
rect 30604 36430 30606 36482
rect 30606 36430 30658 36482
rect 30658 36430 30660 36482
rect 30604 36428 30660 36430
rect 31612 37154 31668 37156
rect 31612 37102 31614 37154
rect 31614 37102 31666 37154
rect 31666 37102 31668 37154
rect 31612 37100 31668 37102
rect 32060 33346 32116 33348
rect 32060 33294 32062 33346
rect 32062 33294 32114 33346
rect 32114 33294 32116 33346
rect 32060 33292 32116 33294
rect 30828 31388 30884 31444
rect 30604 29986 30660 29988
rect 30604 29934 30606 29986
rect 30606 29934 30658 29986
rect 30658 29934 30660 29986
rect 30604 29932 30660 29934
rect 30380 29484 30436 29540
rect 29932 29372 29988 29428
rect 29372 27804 29428 27860
rect 29148 27580 29204 27636
rect 29148 27020 29204 27076
rect 29820 27916 29876 27972
rect 28364 25564 28420 25620
rect 28364 25228 28420 25284
rect 27804 24050 27860 24052
rect 27804 23998 27806 24050
rect 27806 23998 27858 24050
rect 27858 23998 27860 24050
rect 27804 23996 27860 23998
rect 28588 25282 28644 25284
rect 28588 25230 28590 25282
rect 28590 25230 28642 25282
rect 28642 25230 28644 25282
rect 28588 25228 28644 25230
rect 29596 24668 29652 24724
rect 29036 23884 29092 23940
rect 25788 23212 25844 23268
rect 25452 22988 25508 23044
rect 25340 22876 25396 22932
rect 25004 21980 25060 22036
rect 24892 21420 24948 21476
rect 23772 20130 23828 20132
rect 23772 20078 23774 20130
rect 23774 20078 23826 20130
rect 23826 20078 23828 20130
rect 23772 20076 23828 20078
rect 23548 18620 23604 18676
rect 23212 17666 23268 17668
rect 23212 17614 23214 17666
rect 23214 17614 23266 17666
rect 23266 17614 23268 17666
rect 23212 17612 23268 17614
rect 22540 17276 22596 17332
rect 22652 16828 22708 16884
rect 22428 16268 22484 16324
rect 23436 17500 23492 17556
rect 23100 16044 23156 16100
rect 22764 15484 22820 15540
rect 22540 14924 22596 14980
rect 22204 13356 22260 13412
rect 22204 12402 22260 12404
rect 22204 12350 22206 12402
rect 22206 12350 22258 12402
rect 22258 12350 22260 12402
rect 22204 12348 22260 12350
rect 22428 12796 22484 12852
rect 22092 8876 22148 8932
rect 22204 11004 22260 11060
rect 22204 10556 22260 10612
rect 21980 8428 22036 8484
rect 20636 8034 20692 8036
rect 20636 7982 20638 8034
rect 20638 7982 20690 8034
rect 20690 7982 20692 8034
rect 20636 7980 20692 7982
rect 20412 7756 20468 7812
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20188 6076 20244 6132
rect 19852 6018 19908 6020
rect 19852 5966 19854 6018
rect 19854 5966 19906 6018
rect 19906 5966 19908 6018
rect 19852 5964 19908 5966
rect 20300 5180 20356 5236
rect 21308 7756 21364 7812
rect 21308 7308 21364 7364
rect 21420 7420 21476 7476
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20524 6412 20580 6468
rect 19740 4508 19796 4564
rect 18620 4060 18676 4116
rect 19516 4060 19572 4116
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 21532 7308 21588 7364
rect 20972 6076 21028 6132
rect 20860 5740 20916 5796
rect 21308 5964 21364 6020
rect 21644 6690 21700 6692
rect 21644 6638 21646 6690
rect 21646 6638 21698 6690
rect 21698 6638 21700 6690
rect 21644 6636 21700 6638
rect 21196 5906 21252 5908
rect 21196 5854 21198 5906
rect 21198 5854 21250 5906
rect 21250 5854 21252 5906
rect 21196 5852 21252 5854
rect 23100 11394 23156 11396
rect 23100 11342 23102 11394
rect 23102 11342 23154 11394
rect 23154 11342 23156 11394
rect 23100 11340 23156 11342
rect 22652 11116 22708 11172
rect 21420 5234 21476 5236
rect 21420 5182 21422 5234
rect 21422 5182 21474 5234
rect 21474 5182 21476 5234
rect 21420 5180 21476 5182
rect 21532 5122 21588 5124
rect 21532 5070 21534 5122
rect 21534 5070 21586 5122
rect 21586 5070 21588 5122
rect 21532 5068 21588 5070
rect 21756 5740 21812 5796
rect 22204 5906 22260 5908
rect 22204 5854 22206 5906
rect 22206 5854 22258 5906
rect 22258 5854 22260 5906
rect 22204 5852 22260 5854
rect 22092 5628 22148 5684
rect 23212 11004 23268 11060
rect 23324 12236 23380 12292
rect 23436 12684 23492 12740
rect 24556 19906 24612 19908
rect 24556 19854 24558 19906
rect 24558 19854 24610 19906
rect 24610 19854 24612 19906
rect 24556 19852 24612 19854
rect 24780 19292 24836 19348
rect 24108 18508 24164 18564
rect 23884 18396 23940 18452
rect 23884 16828 23940 16884
rect 23772 16770 23828 16772
rect 23772 16718 23774 16770
rect 23774 16718 23826 16770
rect 23826 16718 23828 16770
rect 23772 16716 23828 16718
rect 23660 15596 23716 15652
rect 24220 18450 24276 18452
rect 24220 18398 24222 18450
rect 24222 18398 24274 18450
rect 24274 18398 24276 18450
rect 24220 18396 24276 18398
rect 24668 18060 24724 18116
rect 24668 17106 24724 17108
rect 24668 17054 24670 17106
rect 24670 17054 24722 17106
rect 24722 17054 24724 17106
rect 24668 17052 24724 17054
rect 24332 15874 24388 15876
rect 24332 15822 24334 15874
rect 24334 15822 24386 15874
rect 24386 15822 24388 15874
rect 24332 15820 24388 15822
rect 24332 15372 24388 15428
rect 24220 14812 24276 14868
rect 24108 14642 24164 14644
rect 24108 14590 24110 14642
rect 24110 14590 24162 14642
rect 24162 14590 24164 14642
rect 24108 14588 24164 14590
rect 26124 22988 26180 23044
rect 26012 22876 26068 22932
rect 26124 21980 26180 22036
rect 25788 21644 25844 21700
rect 26124 20748 26180 20804
rect 25452 19964 25508 20020
rect 26124 19852 26180 19908
rect 25340 18338 25396 18340
rect 25340 18286 25342 18338
rect 25342 18286 25394 18338
rect 25394 18286 25396 18338
rect 25340 18284 25396 18286
rect 25004 17612 25060 17668
rect 26236 18284 26292 18340
rect 25676 16658 25732 16660
rect 25676 16606 25678 16658
rect 25678 16606 25730 16658
rect 25730 16606 25732 16658
rect 25676 16604 25732 16606
rect 26012 16604 26068 16660
rect 24892 14812 24948 14868
rect 25116 15596 25172 15652
rect 25004 14642 25060 14644
rect 25004 14590 25006 14642
rect 25006 14590 25058 14642
rect 25058 14590 25060 14642
rect 25004 14588 25060 14590
rect 24780 14476 24836 14532
rect 25228 15314 25284 15316
rect 25228 15262 25230 15314
rect 25230 15262 25282 15314
rect 25282 15262 25284 15314
rect 25228 15260 25284 15262
rect 26012 15426 26068 15428
rect 26012 15374 26014 15426
rect 26014 15374 26066 15426
rect 26066 15374 26068 15426
rect 26012 15372 26068 15374
rect 25452 14700 25508 14756
rect 25900 14588 25956 14644
rect 26012 15148 26068 15204
rect 25788 14530 25844 14532
rect 25788 14478 25790 14530
rect 25790 14478 25842 14530
rect 25842 14478 25844 14530
rect 25788 14476 25844 14478
rect 23996 12908 24052 12964
rect 24332 12178 24388 12180
rect 24332 12126 24334 12178
rect 24334 12126 24386 12178
rect 24386 12126 24388 12178
rect 24332 12124 24388 12126
rect 24556 12012 24612 12068
rect 24220 11394 24276 11396
rect 24220 11342 24222 11394
rect 24222 11342 24274 11394
rect 24274 11342 24276 11394
rect 24220 11340 24276 11342
rect 24668 11452 24724 11508
rect 23212 10050 23268 10052
rect 23212 9998 23214 10050
rect 23214 9998 23266 10050
rect 23266 9998 23268 10050
rect 23212 9996 23268 9998
rect 23996 9884 24052 9940
rect 24108 10108 24164 10164
rect 23324 9660 23380 9716
rect 23324 8876 23380 8932
rect 22988 7644 23044 7700
rect 24668 9996 24724 10052
rect 25228 12738 25284 12740
rect 25228 12686 25230 12738
rect 25230 12686 25282 12738
rect 25282 12686 25284 12738
rect 25228 12684 25284 12686
rect 26348 15260 26404 15316
rect 26684 22988 26740 23044
rect 26796 22876 26852 22932
rect 27244 23324 27300 23380
rect 27692 23714 27748 23716
rect 27692 23662 27694 23714
rect 27694 23662 27746 23714
rect 27746 23662 27748 23714
rect 27692 23660 27748 23662
rect 29372 23714 29428 23716
rect 29372 23662 29374 23714
rect 29374 23662 29426 23714
rect 29426 23662 29428 23714
rect 29372 23660 29428 23662
rect 27244 22764 27300 22820
rect 27916 23378 27972 23380
rect 27916 23326 27918 23378
rect 27918 23326 27970 23378
rect 27970 23326 27972 23378
rect 27916 23324 27972 23326
rect 29372 23324 29428 23380
rect 28364 22540 28420 22596
rect 26572 21196 26628 21252
rect 26684 21980 26740 22036
rect 26572 16156 26628 16212
rect 26572 15820 26628 15876
rect 26908 22316 26964 22372
rect 27132 21756 27188 21812
rect 27580 22370 27636 22372
rect 27580 22318 27582 22370
rect 27582 22318 27634 22370
rect 27634 22318 27636 22370
rect 27580 22316 27636 22318
rect 27244 21586 27300 21588
rect 27244 21534 27246 21586
rect 27246 21534 27298 21586
rect 27298 21534 27300 21586
rect 27244 21532 27300 21534
rect 27020 21420 27076 21476
rect 27244 21084 27300 21140
rect 26796 20748 26852 20804
rect 27132 20802 27188 20804
rect 27132 20750 27134 20802
rect 27134 20750 27186 20802
rect 27186 20750 27188 20802
rect 27132 20748 27188 20750
rect 27916 22258 27972 22260
rect 27916 22206 27918 22258
rect 27918 22206 27970 22258
rect 27970 22206 27972 22258
rect 27916 22204 27972 22206
rect 28028 21698 28084 21700
rect 28028 21646 28030 21698
rect 28030 21646 28082 21698
rect 28082 21646 28084 21698
rect 28028 21644 28084 21646
rect 27804 21532 27860 21588
rect 29036 22316 29092 22372
rect 29260 22370 29316 22372
rect 29260 22318 29262 22370
rect 29262 22318 29314 22370
rect 29314 22318 29316 22370
rect 29260 22316 29316 22318
rect 29036 21980 29092 22036
rect 29148 22204 29204 22260
rect 28588 21868 28644 21924
rect 28588 21532 28644 21588
rect 28364 21474 28420 21476
rect 28364 21422 28366 21474
rect 28366 21422 28418 21474
rect 28418 21422 28420 21474
rect 28364 21420 28420 21422
rect 28364 21196 28420 21252
rect 27804 20802 27860 20804
rect 27804 20750 27806 20802
rect 27806 20750 27858 20802
rect 27858 20750 27860 20802
rect 27804 20748 27860 20750
rect 26796 17052 26852 17108
rect 26908 16380 26964 16436
rect 27468 20188 27524 20244
rect 27244 16380 27300 16436
rect 27468 16716 27524 16772
rect 27356 15372 27412 15428
rect 26012 13692 26068 13748
rect 26348 13858 26404 13860
rect 26348 13806 26350 13858
rect 26350 13806 26402 13858
rect 26402 13806 26404 13858
rect 26348 13804 26404 13806
rect 26796 13804 26852 13860
rect 26684 13746 26740 13748
rect 26684 13694 26686 13746
rect 26686 13694 26738 13746
rect 26738 13694 26740 13746
rect 26684 13692 26740 13694
rect 26124 13132 26180 13188
rect 26012 12684 26068 12740
rect 26348 13132 26404 13188
rect 26460 12962 26516 12964
rect 26460 12910 26462 12962
rect 26462 12910 26514 12962
rect 26514 12910 26516 12962
rect 26460 12908 26516 12910
rect 26348 12348 26404 12404
rect 25228 12066 25284 12068
rect 25228 12014 25230 12066
rect 25230 12014 25282 12066
rect 25282 12014 25284 12066
rect 25228 12012 25284 12014
rect 25004 9714 25060 9716
rect 25004 9662 25006 9714
rect 25006 9662 25058 9714
rect 25058 9662 25060 9714
rect 25004 9660 25060 9662
rect 25228 9042 25284 9044
rect 25228 8990 25230 9042
rect 25230 8990 25282 9042
rect 25282 8990 25284 9042
rect 25228 8988 25284 8990
rect 25004 8876 25060 8932
rect 24556 8540 24612 8596
rect 24220 8316 24276 8372
rect 23884 8034 23940 8036
rect 23884 7982 23886 8034
rect 23886 7982 23938 8034
rect 23938 7982 23940 8034
rect 23884 7980 23940 7982
rect 22876 7474 22932 7476
rect 22876 7422 22878 7474
rect 22878 7422 22930 7474
rect 22930 7422 22932 7474
rect 22876 7420 22932 7422
rect 24892 8316 24948 8372
rect 23436 7362 23492 7364
rect 23436 7310 23438 7362
rect 23438 7310 23490 7362
rect 23490 7310 23492 7362
rect 23436 7308 23492 7310
rect 22876 5628 22932 5684
rect 23436 5740 23492 5796
rect 21644 4732 21700 4788
rect 22316 4956 22372 5012
rect 23100 4956 23156 5012
rect 24668 7756 24724 7812
rect 26012 11452 26068 11508
rect 26908 12962 26964 12964
rect 26908 12910 26910 12962
rect 26910 12910 26962 12962
rect 26962 12910 26964 12962
rect 26908 12908 26964 12910
rect 28028 16268 28084 16324
rect 27580 16156 27636 16212
rect 28700 21362 28756 21364
rect 28700 21310 28702 21362
rect 28702 21310 28754 21362
rect 28754 21310 28756 21362
rect 28700 21308 28756 21310
rect 28588 20748 28644 20804
rect 28700 20300 28756 20356
rect 28252 17554 28308 17556
rect 28252 17502 28254 17554
rect 28254 17502 28306 17554
rect 28306 17502 28308 17554
rect 28252 17500 28308 17502
rect 29596 21868 29652 21924
rect 29260 20802 29316 20804
rect 29260 20750 29262 20802
rect 29262 20750 29314 20802
rect 29314 20750 29316 20802
rect 29260 20748 29316 20750
rect 29260 20300 29316 20356
rect 29820 27020 29876 27076
rect 30492 28588 30548 28644
rect 29932 26572 29988 26628
rect 30044 27692 30100 27748
rect 30268 27132 30324 27188
rect 32060 29484 32116 29540
rect 31164 28924 31220 28980
rect 31836 28588 31892 28644
rect 32508 38780 32564 38836
rect 33516 38834 33572 38836
rect 33516 38782 33518 38834
rect 33518 38782 33570 38834
rect 33570 38782 33572 38834
rect 33516 38780 33572 38782
rect 34748 39394 34804 39396
rect 34748 39342 34750 39394
rect 34750 39342 34802 39394
rect 34802 39342 34804 39394
rect 34748 39340 34804 39342
rect 32396 37378 32452 37380
rect 32396 37326 32398 37378
rect 32398 37326 32450 37378
rect 32450 37326 32452 37378
rect 32396 37324 32452 37326
rect 33516 37324 33572 37380
rect 33964 36988 34020 37044
rect 34188 36428 34244 36484
rect 34300 35308 34356 35364
rect 33628 35084 33684 35140
rect 32396 32508 32452 32564
rect 32956 33292 33012 33348
rect 33516 32562 33572 32564
rect 33516 32510 33518 32562
rect 33518 32510 33570 32562
rect 33570 32510 33572 32562
rect 33516 32508 33572 32510
rect 32620 32396 32676 32452
rect 32284 28700 32340 28756
rect 31500 27746 31556 27748
rect 31500 27694 31502 27746
rect 31502 27694 31554 27746
rect 31554 27694 31556 27746
rect 31500 27692 31556 27694
rect 30716 27186 30772 27188
rect 30716 27134 30718 27186
rect 30718 27134 30770 27186
rect 30770 27134 30772 27186
rect 30716 27132 30772 27134
rect 30380 27020 30436 27076
rect 31164 27074 31220 27076
rect 31164 27022 31166 27074
rect 31166 27022 31218 27074
rect 31218 27022 31220 27074
rect 31164 27020 31220 27022
rect 31836 27020 31892 27076
rect 31724 26962 31780 26964
rect 31724 26910 31726 26962
rect 31726 26910 31778 26962
rect 31778 26910 31780 26962
rect 31724 26908 31780 26910
rect 31724 26572 31780 26628
rect 30044 24722 30100 24724
rect 30044 24670 30046 24722
rect 30046 24670 30098 24722
rect 30098 24670 30100 24722
rect 30044 24668 30100 24670
rect 30940 26290 30996 26292
rect 30940 26238 30942 26290
rect 30942 26238 30994 26290
rect 30994 26238 30996 26290
rect 30940 26236 30996 26238
rect 29932 23938 29988 23940
rect 29932 23886 29934 23938
rect 29934 23886 29986 23938
rect 29986 23886 29988 23938
rect 29932 23884 29988 23886
rect 30380 23938 30436 23940
rect 30380 23886 30382 23938
rect 30382 23886 30434 23938
rect 30434 23886 30436 23938
rect 30380 23884 30436 23886
rect 30604 23436 30660 23492
rect 30156 22428 30212 22484
rect 29820 22316 29876 22372
rect 30268 21698 30324 21700
rect 30268 21646 30270 21698
rect 30270 21646 30322 21698
rect 30322 21646 30324 21698
rect 30268 21644 30324 21646
rect 30604 22482 30660 22484
rect 30604 22430 30606 22482
rect 30606 22430 30658 22482
rect 30658 22430 30660 22482
rect 30604 22428 30660 22430
rect 30716 21980 30772 22036
rect 30604 21644 30660 21700
rect 29708 20914 29764 20916
rect 29708 20862 29710 20914
rect 29710 20862 29762 20914
rect 29762 20862 29764 20914
rect 29708 20860 29764 20862
rect 29372 18956 29428 19012
rect 30492 20860 30548 20916
rect 30380 20300 30436 20356
rect 29372 17948 29428 18004
rect 29596 17948 29652 18004
rect 29708 17500 29764 17556
rect 28588 17276 28644 17332
rect 28364 17052 28420 17108
rect 28364 16268 28420 16324
rect 29596 16716 29652 16772
rect 28476 16156 28532 16212
rect 29260 16268 29316 16324
rect 30044 17276 30100 17332
rect 30044 16210 30100 16212
rect 30044 16158 30046 16210
rect 30046 16158 30098 16210
rect 30098 16158 30100 16210
rect 30044 16156 30100 16158
rect 28588 15484 28644 15540
rect 29932 15484 29988 15540
rect 29260 15372 29316 15428
rect 27804 14140 27860 14196
rect 28140 13746 28196 13748
rect 28140 13694 28142 13746
rect 28142 13694 28194 13746
rect 28194 13694 28196 13746
rect 28140 13692 28196 13694
rect 26236 10722 26292 10724
rect 26236 10670 26238 10722
rect 26238 10670 26290 10722
rect 26290 10670 26292 10722
rect 26236 10668 26292 10670
rect 25676 10108 25732 10164
rect 25676 8930 25732 8932
rect 25676 8878 25678 8930
rect 25678 8878 25730 8930
rect 25730 8878 25732 8930
rect 25676 8876 25732 8878
rect 25564 8540 25620 8596
rect 26124 8540 26180 8596
rect 25452 8204 25508 8260
rect 24444 6690 24500 6692
rect 24444 6638 24446 6690
rect 24446 6638 24498 6690
rect 24498 6638 24500 6690
rect 24444 6636 24500 6638
rect 24108 5628 24164 5684
rect 23884 5010 23940 5012
rect 23884 4958 23886 5010
rect 23886 4958 23938 5010
rect 23938 4958 23940 5010
rect 23884 4956 23940 4958
rect 24780 5852 24836 5908
rect 25116 8146 25172 8148
rect 25116 8094 25118 8146
rect 25118 8094 25170 8146
rect 25170 8094 25172 8146
rect 25116 8092 25172 8094
rect 27020 12124 27076 12180
rect 27580 11452 27636 11508
rect 29148 14588 29204 14644
rect 28476 14530 28532 14532
rect 28476 14478 28478 14530
rect 28478 14478 28530 14530
rect 28530 14478 28532 14530
rect 28476 14476 28532 14478
rect 29484 14530 29540 14532
rect 29484 14478 29486 14530
rect 29486 14478 29538 14530
rect 29538 14478 29540 14530
rect 29484 14476 29540 14478
rect 30044 15314 30100 15316
rect 30044 15262 30046 15314
rect 30046 15262 30098 15314
rect 30098 15262 30100 15314
rect 30044 15260 30100 15262
rect 30380 17724 30436 17780
rect 30604 16940 30660 16996
rect 30268 15932 30324 15988
rect 30492 15314 30548 15316
rect 30492 15262 30494 15314
rect 30494 15262 30546 15314
rect 30546 15262 30548 15314
rect 30492 15260 30548 15262
rect 31500 24332 31556 24388
rect 31052 23938 31108 23940
rect 31052 23886 31054 23938
rect 31054 23886 31106 23938
rect 31106 23886 31108 23938
rect 31052 23884 31108 23886
rect 31388 23714 31444 23716
rect 31388 23662 31390 23714
rect 31390 23662 31442 23714
rect 31442 23662 31444 23714
rect 31388 23660 31444 23662
rect 32172 27804 32228 27860
rect 32172 27356 32228 27412
rect 31836 24108 31892 24164
rect 32396 27468 32452 27524
rect 32396 26012 32452 26068
rect 32284 25228 32340 25284
rect 34300 32284 34356 32340
rect 33180 29932 33236 29988
rect 33068 29596 33124 29652
rect 32956 28754 33012 28756
rect 32956 28702 32958 28754
rect 32958 28702 33010 28754
rect 33010 28702 33012 28754
rect 32956 28700 33012 28702
rect 32844 28642 32900 28644
rect 32844 28590 32846 28642
rect 32846 28590 32898 28642
rect 32898 28590 32900 28642
rect 32844 28588 32900 28590
rect 32956 28476 33012 28532
rect 33404 29148 33460 29204
rect 33516 29538 33572 29540
rect 33516 29486 33518 29538
rect 33518 29486 33570 29538
rect 33570 29486 33572 29538
rect 33516 29484 33572 29486
rect 33964 29036 34020 29092
rect 36316 38892 36372 38948
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35420 37100 35476 37156
rect 34860 36988 34916 37044
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34748 34860 34804 34916
rect 35868 36988 35924 37044
rect 36092 37938 36148 37940
rect 36092 37886 36094 37938
rect 36094 37886 36146 37938
rect 36146 37886 36148 37938
rect 36092 37884 36148 37886
rect 35980 37100 36036 37156
rect 36092 37324 36148 37380
rect 36988 37938 37044 37940
rect 36988 37886 36990 37938
rect 36990 37886 37042 37938
rect 37042 37886 37044 37938
rect 36988 37884 37044 37886
rect 36204 36482 36260 36484
rect 36204 36430 36206 36482
rect 36206 36430 36258 36482
rect 36258 36430 36260 36482
rect 36204 36428 36260 36430
rect 37660 38780 37716 38836
rect 37772 39004 37828 39060
rect 38556 38834 38612 38836
rect 38556 38782 38558 38834
rect 38558 38782 38610 38834
rect 38610 38782 38612 38834
rect 38556 38780 38612 38782
rect 37100 37212 37156 37268
rect 37436 37660 37492 37716
rect 36652 36988 36708 37044
rect 37100 36988 37156 37044
rect 35756 34412 35812 34468
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 33516 28588 33572 28644
rect 33628 28924 33684 28980
rect 33404 28082 33460 28084
rect 33404 28030 33406 28082
rect 33406 28030 33458 28082
rect 33458 28030 33460 28082
rect 33404 28028 33460 28030
rect 33964 28028 34020 28084
rect 33068 27804 33124 27860
rect 33852 27468 33908 27524
rect 33068 26684 33124 26740
rect 33292 26348 33348 26404
rect 32844 26012 32900 26068
rect 34300 28028 34356 28084
rect 35756 31836 35812 31892
rect 34636 31106 34692 31108
rect 34636 31054 34638 31106
rect 34638 31054 34690 31106
rect 34690 31054 34692 31106
rect 34636 31052 34692 31054
rect 34748 30098 34804 30100
rect 34748 30046 34750 30098
rect 34750 30046 34802 30098
rect 34802 30046 34804 30098
rect 34748 30044 34804 30046
rect 34188 27916 34244 27972
rect 34300 27858 34356 27860
rect 34300 27806 34302 27858
rect 34302 27806 34354 27858
rect 34354 27806 34356 27858
rect 34300 27804 34356 27806
rect 34076 27020 34132 27076
rect 34300 26236 34356 26292
rect 33852 25676 33908 25732
rect 33740 25340 33796 25396
rect 34748 29596 34804 29652
rect 34748 29372 34804 29428
rect 35532 30882 35588 30884
rect 35532 30830 35534 30882
rect 35534 30830 35586 30882
rect 35586 30830 35588 30882
rect 35532 30828 35588 30830
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34860 29036 34916 29092
rect 34524 28642 34580 28644
rect 34524 28590 34526 28642
rect 34526 28590 34578 28642
rect 34578 28590 34580 28642
rect 34524 28588 34580 28590
rect 34748 28028 34804 28084
rect 34524 27074 34580 27076
rect 34524 27022 34526 27074
rect 34526 27022 34578 27074
rect 34578 27022 34580 27074
rect 34524 27020 34580 27022
rect 34524 26460 34580 26516
rect 34412 26124 34468 26180
rect 34972 28476 35028 28532
rect 35532 29596 35588 29652
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 36428 32396 36484 32452
rect 36428 32060 36484 32116
rect 37548 37324 37604 37380
rect 37436 37154 37492 37156
rect 37436 37102 37438 37154
rect 37438 37102 37490 37154
rect 37490 37102 37492 37154
rect 37436 37100 37492 37102
rect 37660 36316 37716 36372
rect 37548 36258 37604 36260
rect 37548 36206 37550 36258
rect 37550 36206 37602 36258
rect 37602 36206 37604 36258
rect 37548 36204 37604 36206
rect 37660 34802 37716 34804
rect 37660 34750 37662 34802
rect 37662 34750 37714 34802
rect 37714 34750 37716 34802
rect 37660 34748 37716 34750
rect 37100 34690 37156 34692
rect 37100 34638 37102 34690
rect 37102 34638 37154 34690
rect 37154 34638 37156 34690
rect 37100 34636 37156 34638
rect 37212 34412 37268 34468
rect 36988 34018 37044 34020
rect 36988 33966 36990 34018
rect 36990 33966 37042 34018
rect 37042 33966 37044 34018
rect 36988 33964 37044 33966
rect 37212 33628 37268 33684
rect 36540 31836 36596 31892
rect 36764 32508 36820 32564
rect 36540 31276 36596 31332
rect 36092 30828 36148 30884
rect 35756 30098 35812 30100
rect 35756 30046 35758 30098
rect 35758 30046 35810 30098
rect 35810 30046 35812 30098
rect 35756 30044 35812 30046
rect 36988 32396 37044 32452
rect 38108 37154 38164 37156
rect 38108 37102 38110 37154
rect 38110 37102 38162 37154
rect 38162 37102 38164 37154
rect 38108 37100 38164 37102
rect 37996 36988 38052 37044
rect 38556 38556 38612 38612
rect 38220 36428 38276 36484
rect 38444 37660 38500 37716
rect 38108 36370 38164 36372
rect 38108 36318 38110 36370
rect 38110 36318 38162 36370
rect 38162 36318 38164 36370
rect 38108 36316 38164 36318
rect 37436 34130 37492 34132
rect 37436 34078 37438 34130
rect 37438 34078 37490 34130
rect 37490 34078 37492 34130
rect 37436 34076 37492 34078
rect 37660 33122 37716 33124
rect 37660 33070 37662 33122
rect 37662 33070 37714 33122
rect 37714 33070 37716 33122
rect 37660 33068 37716 33070
rect 37548 31890 37604 31892
rect 37548 31838 37550 31890
rect 37550 31838 37602 31890
rect 37602 31838 37604 31890
rect 37548 31836 37604 31838
rect 37324 31276 37380 31332
rect 37548 31052 37604 31108
rect 36876 30828 36932 30884
rect 37324 30828 37380 30884
rect 36316 29484 36372 29540
rect 35868 28812 35924 28868
rect 35196 27132 35252 27188
rect 35084 26850 35140 26852
rect 35084 26798 35086 26850
rect 35086 26798 35138 26850
rect 35138 26798 35140 26850
rect 35084 26796 35140 26798
rect 36764 30380 36820 30436
rect 36428 29036 36484 29092
rect 36540 28812 36596 28868
rect 36316 28476 36372 28532
rect 36092 27074 36148 27076
rect 36092 27022 36094 27074
rect 36094 27022 36146 27074
rect 36146 27022 36148 27074
rect 36092 27020 36148 27022
rect 35756 26572 35812 26628
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34300 25340 34356 25396
rect 35196 25676 35252 25732
rect 36428 25506 36484 25508
rect 36428 25454 36430 25506
rect 36430 25454 36482 25506
rect 36482 25454 36484 25506
rect 36428 25452 36484 25454
rect 36764 25452 36820 25508
rect 35644 25340 35700 25396
rect 32620 23884 32676 23940
rect 32732 23772 32788 23828
rect 31500 23324 31556 23380
rect 32284 23378 32340 23380
rect 32284 23326 32286 23378
rect 32286 23326 32338 23378
rect 32338 23326 32340 23378
rect 32284 23324 32340 23326
rect 32620 23100 32676 23156
rect 32284 22204 32340 22260
rect 31164 21868 31220 21924
rect 31276 21644 31332 21700
rect 32284 21980 32340 22036
rect 31500 21586 31556 21588
rect 31500 21534 31502 21586
rect 31502 21534 31554 21586
rect 31554 21534 31556 21586
rect 31500 21532 31556 21534
rect 31164 21308 31220 21364
rect 32060 20972 32116 21028
rect 31724 20018 31780 20020
rect 31724 19966 31726 20018
rect 31726 19966 31778 20018
rect 31778 19966 31780 20018
rect 31724 19964 31780 19966
rect 32172 19628 32228 19684
rect 31724 18338 31780 18340
rect 31724 18286 31726 18338
rect 31726 18286 31778 18338
rect 31778 18286 31780 18338
rect 31724 18284 31780 18286
rect 31388 17724 31444 17780
rect 30828 16940 30884 16996
rect 30940 16716 30996 16772
rect 31724 17666 31780 17668
rect 31724 17614 31726 17666
rect 31726 17614 31778 17666
rect 31778 17614 31780 17666
rect 31724 17612 31780 17614
rect 31052 15538 31108 15540
rect 31052 15486 31054 15538
rect 31054 15486 31106 15538
rect 31106 15486 31108 15538
rect 31052 15484 31108 15486
rect 32508 19740 32564 19796
rect 32396 19068 32452 19124
rect 31948 18562 32004 18564
rect 31948 18510 31950 18562
rect 31950 18510 32002 18562
rect 32002 18510 32004 18562
rect 31948 18508 32004 18510
rect 30268 14476 30324 14532
rect 29484 14140 29540 14196
rect 28252 12348 28308 12404
rect 29260 13244 29316 13300
rect 28476 12236 28532 12292
rect 27804 11452 27860 11508
rect 27804 10668 27860 10724
rect 29148 11170 29204 11172
rect 29148 11118 29150 11170
rect 29150 11118 29202 11170
rect 29202 11118 29204 11170
rect 29148 11116 29204 11118
rect 29260 10444 29316 10500
rect 29708 13916 29764 13972
rect 29596 11900 29652 11956
rect 29596 11506 29652 11508
rect 29596 11454 29598 11506
rect 29598 11454 29650 11506
rect 29650 11454 29652 11506
rect 29596 11452 29652 11454
rect 29596 10498 29652 10500
rect 29596 10446 29598 10498
rect 29598 10446 29650 10498
rect 29650 10446 29652 10498
rect 29596 10444 29652 10446
rect 31164 14306 31220 14308
rect 31164 14254 31166 14306
rect 31166 14254 31218 14306
rect 31218 14254 31220 14306
rect 31164 14252 31220 14254
rect 30492 13916 30548 13972
rect 29820 13356 29876 13412
rect 29932 12796 29988 12852
rect 30380 12796 30436 12852
rect 30268 12572 30324 12628
rect 30268 12402 30324 12404
rect 30268 12350 30270 12402
rect 30270 12350 30322 12402
rect 30322 12350 30324 12402
rect 30268 12348 30324 12350
rect 30156 12012 30212 12068
rect 30268 11788 30324 11844
rect 26908 8764 26964 8820
rect 29596 8428 29652 8484
rect 26796 8204 26852 8260
rect 27244 8204 27300 8260
rect 27020 8146 27076 8148
rect 27020 8094 27022 8146
rect 27022 8094 27074 8146
rect 27074 8094 27076 8146
rect 27020 8092 27076 8094
rect 26908 7980 26964 8036
rect 26796 7698 26852 7700
rect 26796 7646 26798 7698
rect 26798 7646 26850 7698
rect 26850 7646 26852 7698
rect 26796 7644 26852 7646
rect 29484 8204 29540 8260
rect 27580 8146 27636 8148
rect 27580 8094 27582 8146
rect 27582 8094 27634 8146
rect 27634 8094 27636 8146
rect 27580 8092 27636 8094
rect 25340 6636 25396 6692
rect 28364 7420 28420 7476
rect 27580 6748 27636 6804
rect 25676 5906 25732 5908
rect 25676 5854 25678 5906
rect 25678 5854 25730 5906
rect 25730 5854 25732 5906
rect 25676 5852 25732 5854
rect 28364 6748 28420 6804
rect 28588 6636 28644 6692
rect 25228 5740 25284 5796
rect 25452 5682 25508 5684
rect 25452 5630 25454 5682
rect 25454 5630 25506 5682
rect 25506 5630 25508 5682
rect 25452 5628 25508 5630
rect 29484 7474 29540 7476
rect 29484 7422 29486 7474
rect 29486 7422 29538 7474
rect 29538 7422 29540 7474
rect 29484 7420 29540 7422
rect 29148 6636 29204 6692
rect 31724 14812 31780 14868
rect 32732 18396 32788 18452
rect 32508 18060 32564 18116
rect 32284 16828 32340 16884
rect 32172 16098 32228 16100
rect 32172 16046 32174 16098
rect 32174 16046 32226 16098
rect 32226 16046 32228 16098
rect 32172 16044 32228 16046
rect 33180 23436 33236 23492
rect 33180 23100 33236 23156
rect 33516 22876 33572 22932
rect 33628 22988 33684 23044
rect 33852 23154 33908 23156
rect 33852 23102 33854 23154
rect 33854 23102 33906 23154
rect 33906 23102 33908 23154
rect 33852 23100 33908 23102
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34076 23100 34132 23156
rect 33516 22370 33572 22372
rect 33516 22318 33518 22370
rect 33518 22318 33570 22370
rect 33570 22318 33572 22370
rect 33516 22316 33572 22318
rect 33292 21868 33348 21924
rect 32956 21586 33012 21588
rect 32956 21534 32958 21586
rect 32958 21534 33010 21586
rect 33010 21534 33012 21586
rect 32956 21532 33012 21534
rect 33292 20802 33348 20804
rect 33292 20750 33294 20802
rect 33294 20750 33346 20802
rect 33346 20750 33348 20802
rect 33292 20748 33348 20750
rect 33740 21644 33796 21700
rect 33740 21026 33796 21028
rect 33740 20974 33742 21026
rect 33742 20974 33794 21026
rect 33794 20974 33796 21026
rect 33740 20972 33796 20974
rect 33964 21532 34020 21588
rect 33516 20188 33572 20244
rect 33180 20018 33236 20020
rect 33180 19966 33182 20018
rect 33182 19966 33234 20018
rect 33234 19966 33236 20018
rect 33180 19964 33236 19966
rect 33516 19346 33572 19348
rect 33516 19294 33518 19346
rect 33518 19294 33570 19346
rect 33570 19294 33572 19346
rect 33516 19292 33572 19294
rect 32844 16604 32900 16660
rect 33068 18508 33124 18564
rect 33180 18284 33236 18340
rect 33068 16604 33124 16660
rect 32284 15596 32340 15652
rect 33180 15596 33236 15652
rect 32060 14700 32116 14756
rect 32620 14642 32676 14644
rect 32620 14590 32622 14642
rect 32622 14590 32674 14642
rect 32674 14590 32676 14642
rect 32620 14588 32676 14590
rect 32396 14364 32452 14420
rect 32284 14252 32340 14308
rect 31164 13356 31220 13412
rect 31052 12962 31108 12964
rect 31052 12910 31054 12962
rect 31054 12910 31106 12962
rect 31106 12910 31108 12962
rect 31052 12908 31108 12910
rect 30492 11340 30548 11396
rect 30604 12572 30660 12628
rect 30940 12236 30996 12292
rect 31388 13132 31444 13188
rect 31500 12684 31556 12740
rect 31164 11788 31220 11844
rect 31164 9884 31220 9940
rect 31388 9772 31444 9828
rect 30940 9266 30996 9268
rect 30940 9214 30942 9266
rect 30942 9214 30994 9266
rect 30994 9214 30996 9266
rect 30940 9212 30996 9214
rect 31836 12908 31892 12964
rect 31836 11788 31892 11844
rect 31724 11394 31780 11396
rect 31724 11342 31726 11394
rect 31726 11342 31778 11394
rect 31778 11342 31780 11394
rect 31724 11340 31780 11342
rect 32284 13186 32340 13188
rect 32284 13134 32286 13186
rect 32286 13134 32338 13186
rect 32338 13134 32340 13186
rect 32284 13132 32340 13134
rect 32060 12850 32116 12852
rect 32060 12798 32062 12850
rect 32062 12798 32114 12850
rect 32114 12798 32116 12850
rect 32060 12796 32116 12798
rect 32172 12738 32228 12740
rect 32172 12686 32174 12738
rect 32174 12686 32226 12738
rect 32226 12686 32228 12738
rect 32172 12684 32228 12686
rect 33628 18060 33684 18116
rect 35420 23772 35476 23828
rect 36204 23660 36260 23716
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34972 22204 35028 22260
rect 34524 21644 34580 21700
rect 34524 20802 34580 20804
rect 34524 20750 34526 20802
rect 34526 20750 34578 20802
rect 34578 20750 34580 20802
rect 34524 20748 34580 20750
rect 34412 20636 34468 20692
rect 35196 22428 35252 22484
rect 36204 23154 36260 23156
rect 36204 23102 36206 23154
rect 36206 23102 36258 23154
rect 36258 23102 36260 23154
rect 36204 23100 36260 23102
rect 35532 22316 35588 22372
rect 35868 22876 35924 22932
rect 35084 21586 35140 21588
rect 35084 21534 35086 21586
rect 35086 21534 35138 21586
rect 35138 21534 35140 21586
rect 35084 21532 35140 21534
rect 35868 22204 35924 22260
rect 37884 31724 37940 31780
rect 37996 33964 38052 34020
rect 37324 30156 37380 30212
rect 37100 28924 37156 28980
rect 37212 29426 37268 29428
rect 37212 29374 37214 29426
rect 37214 29374 37266 29426
rect 37266 29374 37268 29426
rect 37212 29372 37268 29374
rect 37436 27298 37492 27300
rect 37436 27246 37438 27298
rect 37438 27246 37490 27298
rect 37490 27246 37492 27298
rect 37436 27244 37492 27246
rect 37324 27020 37380 27076
rect 37100 26460 37156 26516
rect 36988 23826 37044 23828
rect 36988 23774 36990 23826
rect 36990 23774 37042 23826
rect 37042 23774 37044 23826
rect 36988 23772 37044 23774
rect 37436 25116 37492 25172
rect 37436 24444 37492 24500
rect 37212 23714 37268 23716
rect 37212 23662 37214 23714
rect 37214 23662 37266 23714
rect 37266 23662 37268 23714
rect 37212 23660 37268 23662
rect 37100 23212 37156 23268
rect 37884 30210 37940 30212
rect 37884 30158 37886 30210
rect 37886 30158 37938 30210
rect 37938 30158 37940 30210
rect 37884 30156 37940 30158
rect 38556 36988 38612 37044
rect 38892 38780 38948 38836
rect 39452 39058 39508 39060
rect 39452 39006 39454 39058
rect 39454 39006 39506 39058
rect 39506 39006 39508 39058
rect 39452 39004 39508 39006
rect 39228 38556 39284 38612
rect 38892 37100 38948 37156
rect 38668 35196 38724 35252
rect 38668 34914 38724 34916
rect 38668 34862 38670 34914
rect 38670 34862 38722 34914
rect 38722 34862 38724 34914
rect 38668 34860 38724 34862
rect 39228 37100 39284 37156
rect 39676 38834 39732 38836
rect 39676 38782 39678 38834
rect 39678 38782 39730 38834
rect 39730 38782 39732 38834
rect 39676 38780 39732 38782
rect 39340 36540 39396 36596
rect 39452 37996 39508 38052
rect 40908 38610 40964 38612
rect 40908 38558 40910 38610
rect 40910 38558 40962 38610
rect 40962 38558 40964 38610
rect 40908 38556 40964 38558
rect 40908 38050 40964 38052
rect 40908 37998 40910 38050
rect 40910 37998 40962 38050
rect 40962 37998 40964 38050
rect 40908 37996 40964 37998
rect 40012 37266 40068 37268
rect 40012 37214 40014 37266
rect 40014 37214 40066 37266
rect 40066 37214 40068 37266
rect 40012 37212 40068 37214
rect 40348 37100 40404 37156
rect 39564 36988 39620 37044
rect 40460 36988 40516 37044
rect 39452 35084 39508 35140
rect 38108 33852 38164 33908
rect 38108 33628 38164 33684
rect 38332 33852 38388 33908
rect 39788 36482 39844 36484
rect 39788 36430 39790 36482
rect 39790 36430 39842 36482
rect 39842 36430 39844 36482
rect 39788 36428 39844 36430
rect 40124 36258 40180 36260
rect 40124 36206 40126 36258
rect 40126 36206 40178 36258
rect 40178 36206 40180 36258
rect 40124 36204 40180 36206
rect 39900 35980 39956 36036
rect 39676 34748 39732 34804
rect 39116 34188 39172 34244
rect 39340 34636 39396 34692
rect 39004 34076 39060 34132
rect 38892 34018 38948 34020
rect 38892 33966 38894 34018
rect 38894 33966 38946 34018
rect 38946 33966 38948 34018
rect 38892 33964 38948 33966
rect 38668 33292 38724 33348
rect 38220 33068 38276 33124
rect 38332 32562 38388 32564
rect 38332 32510 38334 32562
rect 38334 32510 38386 32562
rect 38386 32510 38388 32562
rect 38332 32508 38388 32510
rect 38780 32284 38836 32340
rect 38892 32396 38948 32452
rect 39116 33292 39172 33348
rect 38108 30380 38164 30436
rect 38220 30940 38276 30996
rect 38220 29538 38276 29540
rect 38220 29486 38222 29538
rect 38222 29486 38274 29538
rect 38274 29486 38276 29538
rect 38220 29484 38276 29486
rect 37772 29036 37828 29092
rect 37772 27244 37828 27300
rect 37884 27804 37940 27860
rect 38220 27074 38276 27076
rect 38220 27022 38222 27074
rect 38222 27022 38274 27074
rect 38274 27022 38276 27074
rect 38220 27020 38276 27022
rect 39004 31612 39060 31668
rect 38892 30044 38948 30100
rect 39452 34354 39508 34356
rect 39452 34302 39454 34354
rect 39454 34302 39506 34354
rect 39506 34302 39508 34354
rect 39452 34300 39508 34302
rect 39788 35196 39844 35252
rect 40012 34748 40068 34804
rect 40684 37100 40740 37156
rect 41244 37324 41300 37380
rect 41356 37212 41412 37268
rect 41356 36988 41412 37044
rect 41356 36204 41412 36260
rect 40460 34300 40516 34356
rect 41132 34636 41188 34692
rect 39788 34130 39844 34132
rect 39788 34078 39790 34130
rect 39790 34078 39842 34130
rect 39842 34078 39844 34130
rect 39788 34076 39844 34078
rect 40908 34130 40964 34132
rect 40908 34078 40910 34130
rect 40910 34078 40962 34130
rect 40962 34078 40964 34130
rect 40908 34076 40964 34078
rect 41468 35420 41524 35476
rect 42028 37154 42084 37156
rect 42028 37102 42030 37154
rect 42030 37102 42082 37154
rect 42082 37102 42084 37154
rect 42028 37100 42084 37102
rect 41916 35868 41972 35924
rect 42364 36876 42420 36932
rect 42476 36540 42532 36596
rect 42700 36428 42756 36484
rect 41580 34748 41636 34804
rect 39564 32562 39620 32564
rect 39564 32510 39566 32562
rect 39566 32510 39618 32562
rect 39618 32510 39620 32562
rect 39564 32508 39620 32510
rect 39452 31724 39508 31780
rect 39564 31500 39620 31556
rect 40236 31554 40292 31556
rect 40236 31502 40238 31554
rect 40238 31502 40290 31554
rect 40290 31502 40292 31554
rect 40236 31500 40292 31502
rect 38780 28028 38836 28084
rect 38892 29596 38948 29652
rect 38668 27580 38724 27636
rect 39900 29596 39956 29652
rect 39340 29372 39396 29428
rect 39004 28924 39060 28980
rect 38108 26962 38164 26964
rect 38108 26910 38110 26962
rect 38110 26910 38162 26962
rect 38162 26910 38164 26962
rect 38108 26908 38164 26910
rect 40012 27804 40068 27860
rect 39564 27746 39620 27748
rect 39564 27694 39566 27746
rect 39566 27694 39618 27746
rect 39618 27694 39620 27746
rect 39564 27692 39620 27694
rect 39340 27356 39396 27412
rect 39004 26908 39060 26964
rect 38780 26460 38836 26516
rect 39228 27020 39284 27076
rect 37772 25564 37828 25620
rect 37660 25116 37716 25172
rect 37660 24108 37716 24164
rect 37772 23938 37828 23940
rect 37772 23886 37774 23938
rect 37774 23886 37826 23938
rect 37826 23886 37828 23938
rect 37772 23884 37828 23886
rect 37884 23772 37940 23828
rect 38332 24722 38388 24724
rect 38332 24670 38334 24722
rect 38334 24670 38386 24722
rect 38386 24670 38388 24722
rect 38332 24668 38388 24670
rect 38108 24444 38164 24500
rect 38444 24444 38500 24500
rect 38780 24220 38836 24276
rect 38444 24162 38500 24164
rect 38444 24110 38446 24162
rect 38446 24110 38498 24162
rect 38498 24110 38500 24162
rect 38444 24108 38500 24110
rect 38556 23660 38612 23716
rect 35980 21698 36036 21700
rect 35980 21646 35982 21698
rect 35982 21646 36034 21698
rect 36034 21646 36036 21698
rect 35980 21644 36036 21646
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 36204 21308 36260 21364
rect 34860 20188 34916 20244
rect 34076 19628 34132 19684
rect 33740 17612 33796 17668
rect 33740 16716 33796 16772
rect 35980 20690 36036 20692
rect 35980 20638 35982 20690
rect 35982 20638 36034 20690
rect 36034 20638 36036 20690
rect 35980 20636 36036 20638
rect 35756 20300 35812 20356
rect 34412 19068 34468 19124
rect 34748 19068 34804 19124
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34748 18396 34804 18452
rect 34524 18284 34580 18340
rect 34972 18396 35028 18452
rect 34972 18060 35028 18116
rect 35308 18396 35364 18452
rect 35420 19068 35476 19124
rect 35532 18956 35588 19012
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35084 17836 35140 17892
rect 34972 17612 35028 17668
rect 36092 20130 36148 20132
rect 36092 20078 36094 20130
rect 36094 20078 36146 20130
rect 36146 20078 36148 20130
rect 36092 20076 36148 20078
rect 35756 18956 35812 19012
rect 35868 19068 35924 19124
rect 35644 18620 35700 18676
rect 35308 17500 35364 17556
rect 34188 16716 34244 16772
rect 33852 15484 33908 15540
rect 33292 14588 33348 14644
rect 33180 14530 33236 14532
rect 33180 14478 33182 14530
rect 33182 14478 33234 14530
rect 33234 14478 33236 14530
rect 33180 14476 33236 14478
rect 32956 14418 33012 14420
rect 32956 14366 32958 14418
rect 32958 14366 33010 14418
rect 33010 14366 33012 14418
rect 32956 14364 33012 14366
rect 33628 13746 33684 13748
rect 33628 13694 33630 13746
rect 33630 13694 33682 13746
rect 33682 13694 33684 13746
rect 33628 13692 33684 13694
rect 32508 12572 32564 12628
rect 32172 12124 32228 12180
rect 32172 11506 32228 11508
rect 32172 11454 32174 11506
rect 32174 11454 32226 11506
rect 32226 11454 32228 11506
rect 32172 11452 32228 11454
rect 32508 12348 32564 12404
rect 33852 14754 33908 14756
rect 33852 14702 33854 14754
rect 33854 14702 33906 14754
rect 33906 14702 33908 14754
rect 33852 14700 33908 14702
rect 33964 13858 34020 13860
rect 33964 13806 33966 13858
rect 33966 13806 34018 13858
rect 34018 13806 34020 13858
rect 33964 13804 34020 13806
rect 32732 12962 32788 12964
rect 32732 12910 32734 12962
rect 32734 12910 32786 12962
rect 32786 12910 32788 12962
rect 32732 12908 32788 12910
rect 33180 12684 33236 12740
rect 32844 12124 32900 12180
rect 33180 12124 33236 12180
rect 33068 11900 33124 11956
rect 32956 11116 33012 11172
rect 31948 9884 32004 9940
rect 31724 9266 31780 9268
rect 31724 9214 31726 9266
rect 31726 9214 31778 9266
rect 31778 9214 31780 9266
rect 31724 9212 31780 9214
rect 30716 8428 30772 8484
rect 30604 8316 30660 8372
rect 31836 8316 31892 8372
rect 30044 8092 30100 8148
rect 30156 7308 30212 7364
rect 30156 6690 30212 6692
rect 30156 6638 30158 6690
rect 30158 6638 30210 6690
rect 30210 6638 30212 6690
rect 30156 6636 30212 6638
rect 31276 8258 31332 8260
rect 31276 8206 31278 8258
rect 31278 8206 31330 8258
rect 31330 8206 31332 8258
rect 31276 8204 31332 8206
rect 30828 8092 30884 8148
rect 32060 9826 32116 9828
rect 32060 9774 32062 9826
rect 32062 9774 32114 9826
rect 32114 9774 32116 9826
rect 32060 9772 32116 9774
rect 32060 9266 32116 9268
rect 32060 9214 32062 9266
rect 32062 9214 32114 9266
rect 32114 9214 32116 9266
rect 32060 9212 32116 9214
rect 33740 12908 33796 12964
rect 33628 12572 33684 12628
rect 33404 11900 33460 11956
rect 33852 12124 33908 12180
rect 33180 11452 33236 11508
rect 33292 11676 33348 11732
rect 33740 11676 33796 11732
rect 33516 11116 33572 11172
rect 33404 10556 33460 10612
rect 31948 8092 32004 8148
rect 34300 16492 34356 16548
rect 34412 16268 34468 16324
rect 34076 12348 34132 12404
rect 34412 12012 34468 12068
rect 33628 9772 33684 9828
rect 33628 8428 33684 8484
rect 32844 8092 32900 8148
rect 35532 16604 35588 16660
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 34972 15820 35028 15876
rect 34860 14588 34916 14644
rect 34972 13970 35028 13972
rect 34972 13918 34974 13970
rect 34974 13918 35026 13970
rect 35026 13918 35028 13970
rect 34972 13916 35028 13918
rect 36092 19234 36148 19236
rect 36092 19182 36094 19234
rect 36094 19182 36146 19234
rect 36146 19182 36148 19234
rect 36092 19180 36148 19182
rect 35868 18172 35924 18228
rect 36764 20188 36820 20244
rect 37660 20300 37716 20356
rect 36988 19068 37044 19124
rect 36540 19010 36596 19012
rect 36540 18958 36542 19010
rect 36542 18958 36594 19010
rect 36594 18958 36596 19010
rect 36540 18956 36596 18958
rect 37436 19740 37492 19796
rect 37548 19628 37604 19684
rect 37100 18956 37156 19012
rect 36652 18450 36708 18452
rect 36652 18398 36654 18450
rect 36654 18398 36706 18450
rect 36706 18398 36708 18450
rect 36652 18396 36708 18398
rect 37436 18338 37492 18340
rect 37436 18286 37438 18338
rect 37438 18286 37490 18338
rect 37490 18286 37492 18338
rect 37436 18284 37492 18286
rect 36428 17724 36484 17780
rect 36428 17554 36484 17556
rect 36428 17502 36430 17554
rect 36430 17502 36482 17554
rect 36482 17502 36484 17554
rect 36428 17500 36484 17502
rect 37436 17778 37492 17780
rect 37436 17726 37438 17778
rect 37438 17726 37490 17778
rect 37490 17726 37492 17778
rect 37436 17724 37492 17726
rect 36988 17554 37044 17556
rect 36988 17502 36990 17554
rect 36990 17502 37042 17554
rect 37042 17502 37044 17554
rect 36988 17500 37044 17502
rect 36540 16940 36596 16996
rect 36316 16716 36372 16772
rect 35756 16044 35812 16100
rect 37324 15538 37380 15540
rect 37324 15486 37326 15538
rect 37326 15486 37378 15538
rect 37378 15486 37380 15538
rect 37324 15484 37380 15486
rect 35532 15314 35588 15316
rect 35532 15262 35534 15314
rect 35534 15262 35586 15314
rect 35586 15262 35588 15314
rect 35532 15260 35588 15262
rect 37884 22204 37940 22260
rect 37996 21810 38052 21812
rect 37996 21758 37998 21810
rect 37998 21758 38050 21810
rect 38050 21758 38052 21810
rect 37996 21756 38052 21758
rect 38108 21644 38164 21700
rect 37884 19628 37940 19684
rect 38444 21756 38500 21812
rect 38668 22428 38724 22484
rect 38220 20076 38276 20132
rect 39676 27020 39732 27076
rect 40012 27132 40068 27188
rect 40796 29036 40852 29092
rect 40684 27692 40740 27748
rect 40124 26908 40180 26964
rect 40124 26572 40180 26628
rect 39676 26514 39732 26516
rect 39676 26462 39678 26514
rect 39678 26462 39730 26514
rect 39730 26462 39732 26514
rect 39676 26460 39732 26462
rect 40124 25618 40180 25620
rect 40124 25566 40126 25618
rect 40126 25566 40178 25618
rect 40178 25566 40180 25618
rect 40124 25564 40180 25566
rect 39116 24610 39172 24612
rect 39116 24558 39118 24610
rect 39118 24558 39170 24610
rect 39170 24558 39172 24610
rect 39116 24556 39172 24558
rect 39116 24220 39172 24276
rect 39116 23884 39172 23940
rect 39004 23826 39060 23828
rect 39004 23774 39006 23826
rect 39006 23774 39058 23826
rect 39058 23774 39060 23826
rect 39004 23772 39060 23774
rect 38892 22428 38948 22484
rect 39228 20018 39284 20020
rect 39228 19966 39230 20018
rect 39230 19966 39282 20018
rect 39282 19966 39284 20018
rect 39228 19964 39284 19966
rect 38668 19740 38724 19796
rect 38220 19180 38276 19236
rect 37884 18620 37940 18676
rect 38892 19234 38948 19236
rect 38892 19182 38894 19234
rect 38894 19182 38946 19234
rect 38946 19182 38948 19234
rect 38892 19180 38948 19182
rect 38332 18284 38388 18340
rect 38332 18060 38388 18116
rect 38444 19068 38500 19124
rect 37772 17052 37828 17108
rect 37660 15538 37716 15540
rect 37660 15486 37662 15538
rect 37662 15486 37714 15538
rect 37714 15486 37716 15538
rect 37660 15484 37716 15486
rect 38556 18508 38612 18564
rect 38780 18284 38836 18340
rect 39564 19740 39620 19796
rect 39004 18396 39060 18452
rect 38892 18172 38948 18228
rect 39452 18450 39508 18452
rect 39452 18398 39454 18450
rect 39454 18398 39506 18450
rect 39506 18398 39508 18450
rect 39452 18396 39508 18398
rect 39116 18172 39172 18228
rect 39228 18060 39284 18116
rect 38220 17276 38276 17332
rect 38108 15426 38164 15428
rect 38108 15374 38110 15426
rect 38110 15374 38162 15426
rect 38162 15374 38164 15426
rect 38108 15372 38164 15374
rect 38556 17106 38612 17108
rect 38556 17054 38558 17106
rect 38558 17054 38610 17106
rect 38610 17054 38612 17106
rect 38556 17052 38612 17054
rect 38892 16994 38948 16996
rect 38892 16942 38894 16994
rect 38894 16942 38946 16994
rect 38946 16942 38948 16994
rect 38892 16940 38948 16942
rect 38892 15484 38948 15540
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35532 14530 35588 14532
rect 35532 14478 35534 14530
rect 35534 14478 35586 14530
rect 35586 14478 35588 14530
rect 35532 14476 35588 14478
rect 36988 14140 37044 14196
rect 35420 13858 35476 13860
rect 35420 13806 35422 13858
rect 35422 13806 35474 13858
rect 35474 13806 35476 13858
rect 35420 13804 35476 13806
rect 35308 13746 35364 13748
rect 35308 13694 35310 13746
rect 35310 13694 35362 13746
rect 35362 13694 35364 13746
rect 35308 13692 35364 13694
rect 34860 13132 34916 13188
rect 34860 12236 34916 12292
rect 34524 10556 34580 10612
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 13132 35252 13188
rect 35532 12178 35588 12180
rect 35532 12126 35534 12178
rect 35534 12126 35586 12178
rect 35586 12126 35588 12178
rect 35532 12124 35588 12126
rect 36540 12124 36596 12180
rect 36652 12236 36708 12292
rect 36988 12236 37044 12292
rect 34972 11788 35028 11844
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 37324 13804 37380 13860
rect 37212 12012 37268 12068
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 34636 9826 34692 9828
rect 34636 9774 34638 9826
rect 34638 9774 34690 9826
rect 34690 9774 34692 9826
rect 34636 9772 34692 9774
rect 34076 8146 34132 8148
rect 34076 8094 34078 8146
rect 34078 8094 34130 8146
rect 34130 8094 34132 8146
rect 34076 8092 34132 8094
rect 33964 7474 34020 7476
rect 33964 7422 33966 7474
rect 33966 7422 34018 7474
rect 34018 7422 34020 7474
rect 33964 7420 34020 7422
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35532 8316 35588 8372
rect 35756 8258 35812 8260
rect 35756 8206 35758 8258
rect 35758 8206 35810 8258
rect 35810 8206 35812 8258
rect 35756 8204 35812 8206
rect 37996 15036 38052 15092
rect 37772 14252 37828 14308
rect 38220 14028 38276 14084
rect 37436 9212 37492 9268
rect 37884 12908 37940 12964
rect 37884 12348 37940 12404
rect 37660 12290 37716 12292
rect 37660 12238 37662 12290
rect 37662 12238 37714 12290
rect 37714 12238 37716 12290
rect 37660 12236 37716 12238
rect 37996 12796 38052 12852
rect 38668 15036 38724 15092
rect 38444 13692 38500 13748
rect 38332 12908 38388 12964
rect 38780 13970 38836 13972
rect 38780 13918 38782 13970
rect 38782 13918 38834 13970
rect 38834 13918 38836 13970
rect 38780 13916 38836 13918
rect 40236 25228 40292 25284
rect 40012 24668 40068 24724
rect 39788 24332 39844 24388
rect 39788 23772 39844 23828
rect 40012 21756 40068 21812
rect 39676 18060 39732 18116
rect 39788 19964 39844 20020
rect 39564 17164 39620 17220
rect 39452 16882 39508 16884
rect 39452 16830 39454 16882
rect 39454 16830 39506 16882
rect 39506 16830 39508 16882
rect 39452 16828 39508 16830
rect 39676 17836 39732 17892
rect 39900 19852 39956 19908
rect 39900 19068 39956 19124
rect 40012 18396 40068 18452
rect 40236 23884 40292 23940
rect 40684 25340 40740 25396
rect 41580 31836 41636 31892
rect 41020 30044 41076 30100
rect 41468 30156 41524 30212
rect 41020 29426 41076 29428
rect 41020 29374 41022 29426
rect 41022 29374 41074 29426
rect 41074 29374 41076 29426
rect 41020 29372 41076 29374
rect 41356 29484 41412 29540
rect 41020 27858 41076 27860
rect 41020 27806 41022 27858
rect 41022 27806 41074 27858
rect 41074 27806 41076 27858
rect 41020 27804 41076 27806
rect 41244 27132 41300 27188
rect 41468 28812 41524 28868
rect 41356 27074 41412 27076
rect 41356 27022 41358 27074
rect 41358 27022 41410 27074
rect 41410 27022 41412 27074
rect 41356 27020 41412 27022
rect 40908 25564 40964 25620
rect 40908 25340 40964 25396
rect 42700 34412 42756 34468
rect 43036 36540 43092 36596
rect 43036 35922 43092 35924
rect 43036 35870 43038 35922
rect 43038 35870 43090 35922
rect 43090 35870 43092 35922
rect 43036 35868 43092 35870
rect 42700 33346 42756 33348
rect 42700 33294 42702 33346
rect 42702 33294 42754 33346
rect 42754 33294 42756 33346
rect 42700 33292 42756 33294
rect 42028 30940 42084 30996
rect 41692 30828 41748 30884
rect 44156 37266 44212 37268
rect 44156 37214 44158 37266
rect 44158 37214 44210 37266
rect 44210 37214 44212 37266
rect 44156 37212 44212 37214
rect 43820 37100 43876 37156
rect 43372 36988 43428 37044
rect 43484 36482 43540 36484
rect 43484 36430 43486 36482
rect 43486 36430 43538 36482
rect 43538 36430 43540 36482
rect 43484 36428 43540 36430
rect 43260 35420 43316 35476
rect 43260 32284 43316 32340
rect 42700 31724 42756 31780
rect 42140 30156 42196 30212
rect 41804 29484 41860 29540
rect 41692 28924 41748 28980
rect 43260 30268 43316 30324
rect 42812 29596 42868 29652
rect 42812 29036 42868 29092
rect 41692 27132 41748 27188
rect 42924 28588 42980 28644
rect 43036 29372 43092 29428
rect 42588 27020 42644 27076
rect 41580 26460 41636 26516
rect 40908 24108 40964 24164
rect 41132 23938 41188 23940
rect 41132 23886 41134 23938
rect 41134 23886 41186 23938
rect 41186 23886 41188 23938
rect 41132 23884 41188 23886
rect 40796 23826 40852 23828
rect 40796 23774 40798 23826
rect 40798 23774 40850 23826
rect 40850 23774 40852 23826
rect 40796 23772 40852 23774
rect 41692 25340 41748 25396
rect 41468 25282 41524 25284
rect 41468 25230 41470 25282
rect 41470 25230 41522 25282
rect 41522 25230 41524 25282
rect 41468 25228 41524 25230
rect 40236 19964 40292 20020
rect 41132 21698 41188 21700
rect 41132 21646 41134 21698
rect 41134 21646 41186 21698
rect 41186 21646 41188 21698
rect 41132 21644 41188 21646
rect 41468 21698 41524 21700
rect 41468 21646 41470 21698
rect 41470 21646 41522 21698
rect 41522 21646 41524 21698
rect 41468 21644 41524 21646
rect 41916 25228 41972 25284
rect 41916 24220 41972 24276
rect 42140 25228 42196 25284
rect 43484 30380 43540 30436
rect 43372 29596 43428 29652
rect 43596 30156 43652 30212
rect 43596 29484 43652 29540
rect 43708 28700 43764 28756
rect 44828 36316 44884 36372
rect 44940 35868 44996 35924
rect 44044 34748 44100 34804
rect 44044 33964 44100 34020
rect 45164 34802 45220 34804
rect 45164 34750 45166 34802
rect 45166 34750 45218 34802
rect 45218 34750 45220 34802
rect 45164 34748 45220 34750
rect 45388 34130 45444 34132
rect 45388 34078 45390 34130
rect 45390 34078 45442 34130
rect 45442 34078 45444 34130
rect 45388 34076 45444 34078
rect 44828 33964 44884 34020
rect 44156 33852 44212 33908
rect 45948 33906 46004 33908
rect 45948 33854 45950 33906
rect 45950 33854 46002 33906
rect 46002 33854 46004 33906
rect 45948 33852 46004 33854
rect 45836 33068 45892 33124
rect 43932 32284 43988 32340
rect 45164 32338 45220 32340
rect 45164 32286 45166 32338
rect 45166 32286 45218 32338
rect 45218 32286 45220 32338
rect 45164 32284 45220 32286
rect 45612 31836 45668 31892
rect 44940 31388 44996 31444
rect 44828 30716 44884 30772
rect 44940 30828 44996 30884
rect 44828 30268 44884 30324
rect 44268 30210 44324 30212
rect 44268 30158 44270 30210
rect 44270 30158 44322 30210
rect 44322 30158 44324 30210
rect 44268 30156 44324 30158
rect 45164 30716 45220 30772
rect 45500 30380 45556 30436
rect 45388 30044 45444 30100
rect 44492 29260 44548 29316
rect 43932 28476 43988 28532
rect 45724 30882 45780 30884
rect 45724 30830 45726 30882
rect 45726 30830 45778 30882
rect 45778 30830 45780 30882
rect 45724 30828 45780 30830
rect 45948 29314 46004 29316
rect 45948 29262 45950 29314
rect 45950 29262 46002 29314
rect 46002 29262 46004 29314
rect 45948 29260 46004 29262
rect 45612 28924 45668 28980
rect 43708 27356 43764 27412
rect 43820 28252 43876 28308
rect 40572 19852 40628 19908
rect 40348 19628 40404 19684
rect 41356 19964 41412 20020
rect 42140 20690 42196 20692
rect 42140 20638 42142 20690
rect 42142 20638 42194 20690
rect 42194 20638 42196 20690
rect 42140 20636 42196 20638
rect 42028 20188 42084 20244
rect 40908 19628 40964 19684
rect 40236 19180 40292 19236
rect 40460 19404 40516 19460
rect 39900 16940 39956 16996
rect 39340 15372 39396 15428
rect 40124 15932 40180 15988
rect 39340 14530 39396 14532
rect 39340 14478 39342 14530
rect 39342 14478 39394 14530
rect 39394 14478 39396 14530
rect 39340 14476 39396 14478
rect 39228 13804 39284 13860
rect 38780 12908 38836 12964
rect 38556 12796 38612 12852
rect 38108 12124 38164 12180
rect 38668 12236 38724 12292
rect 38444 12124 38500 12180
rect 38556 12012 38612 12068
rect 37548 9154 37604 9156
rect 37548 9102 37550 9154
rect 37550 9102 37602 9154
rect 37602 9102 37604 9154
rect 37548 9100 37604 9102
rect 37884 9100 37940 9156
rect 38556 9436 38612 9492
rect 38556 8876 38612 8932
rect 34860 7308 34916 7364
rect 36204 7474 36260 7476
rect 36204 7422 36206 7474
rect 36206 7422 36258 7474
rect 36258 7422 36260 7474
rect 36204 7420 36260 7422
rect 35644 7308 35700 7364
rect 39900 13244 39956 13300
rect 42140 19292 42196 19348
rect 41356 18562 41412 18564
rect 41356 18510 41358 18562
rect 41358 18510 41410 18562
rect 41410 18510 41412 18562
rect 41356 18508 41412 18510
rect 42028 17164 42084 17220
rect 42476 23884 42532 23940
rect 43036 23938 43092 23940
rect 43036 23886 43038 23938
rect 43038 23886 43090 23938
rect 43090 23886 43092 23938
rect 43036 23884 43092 23886
rect 43036 23100 43092 23156
rect 42588 22316 42644 22372
rect 42700 21644 42756 21700
rect 42476 20636 42532 20692
rect 42812 20130 42868 20132
rect 42812 20078 42814 20130
rect 42814 20078 42866 20130
rect 42866 20078 42868 20130
rect 42812 20076 42868 20078
rect 42588 19122 42644 19124
rect 42588 19070 42590 19122
rect 42590 19070 42642 19122
rect 42642 19070 42644 19122
rect 42588 19068 42644 19070
rect 42252 17724 42308 17780
rect 41244 16828 41300 16884
rect 40796 15874 40852 15876
rect 40796 15822 40798 15874
rect 40798 15822 40850 15874
rect 40850 15822 40852 15874
rect 40796 15820 40852 15822
rect 40348 13916 40404 13972
rect 41132 14476 41188 14532
rect 40908 13244 40964 13300
rect 40124 12908 40180 12964
rect 41916 16098 41972 16100
rect 41916 16046 41918 16098
rect 41918 16046 41970 16098
rect 41970 16046 41972 16098
rect 41916 16044 41972 16046
rect 42364 16828 42420 16884
rect 41356 15036 41412 15092
rect 44044 28252 44100 28308
rect 44604 28700 44660 28756
rect 44940 28530 44996 28532
rect 44940 28478 44942 28530
rect 44942 28478 44994 28530
rect 44994 28478 44996 28530
rect 44940 28476 44996 28478
rect 44828 28252 44884 28308
rect 44156 26908 44212 26964
rect 44716 26908 44772 26964
rect 44492 24834 44548 24836
rect 44492 24782 44494 24834
rect 44494 24782 44546 24834
rect 44546 24782 44548 24834
rect 44492 24780 44548 24782
rect 45052 26908 45108 26964
rect 45052 24780 45108 24836
rect 44044 24556 44100 24612
rect 44940 24668 44996 24724
rect 44828 24556 44884 24612
rect 44940 23884 44996 23940
rect 44492 23772 44548 23828
rect 44716 23548 44772 23604
rect 43484 22370 43540 22372
rect 43484 22318 43486 22370
rect 43486 22318 43538 22370
rect 43538 22318 43540 22370
rect 43484 22316 43540 22318
rect 43596 21644 43652 21700
rect 45948 24444 46004 24500
rect 45500 23154 45556 23156
rect 45500 23102 45502 23154
rect 45502 23102 45554 23154
rect 45554 23102 45556 23154
rect 45500 23100 45556 23102
rect 43260 20130 43316 20132
rect 43260 20078 43262 20130
rect 43262 20078 43314 20130
rect 43314 20078 43316 20130
rect 43260 20076 43316 20078
rect 43596 18396 43652 18452
rect 43484 16940 43540 16996
rect 43372 16828 43428 16884
rect 44940 18396 44996 18452
rect 44380 17164 44436 17220
rect 45948 18450 46004 18452
rect 45948 18398 45950 18450
rect 45950 18398 46002 18450
rect 46002 18398 46004 18450
rect 45948 18396 46004 18398
rect 45052 16828 45108 16884
rect 45276 16044 45332 16100
rect 43148 14252 43204 14308
rect 43708 13746 43764 13748
rect 43708 13694 43710 13746
rect 43710 13694 43762 13746
rect 43762 13694 43764 13746
rect 43708 13692 43764 13694
rect 41804 12402 41860 12404
rect 41804 12350 41806 12402
rect 41806 12350 41858 12402
rect 41858 12350 41860 12402
rect 41804 12348 41860 12350
rect 41804 12124 41860 12180
rect 41580 11116 41636 11172
rect 39900 9826 39956 9828
rect 39900 9774 39902 9826
rect 39902 9774 39954 9826
rect 39954 9774 39956 9826
rect 39900 9772 39956 9774
rect 41580 9212 41636 9268
rect 41244 9154 41300 9156
rect 41244 9102 41246 9154
rect 41246 9102 41298 9154
rect 41298 9102 41300 9154
rect 41244 9100 41300 9102
rect 43036 12962 43092 12964
rect 43036 12910 43038 12962
rect 43038 12910 43090 12962
rect 43090 12910 43092 12962
rect 43036 12908 43092 12910
rect 45836 12908 45892 12964
rect 42364 12178 42420 12180
rect 42364 12126 42366 12178
rect 42366 12126 42418 12178
rect 42418 12126 42420 12178
rect 42364 12124 42420 12126
rect 42700 12012 42756 12068
rect 42028 11116 42084 11172
rect 43372 9266 43428 9268
rect 43372 9214 43374 9266
rect 43374 9214 43426 9266
rect 43426 9214 43428 9266
rect 43372 9212 43428 9214
rect 41580 8930 41636 8932
rect 41580 8878 41582 8930
rect 41582 8878 41634 8930
rect 41634 8878 41636 8930
rect 41580 8876 41636 8878
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 21196 4114 21252 4116
rect 21196 4062 21198 4114
rect 21198 4062 21250 4114
rect 21250 4062 21252 4114
rect 21196 4060 21252 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
<< metal3 >>
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 1698 43708 1708 43764
rect 1764 43708 1774 43764
rect 1708 43652 1764 43708
rect 700 43596 1764 43652
rect 700 43316 756 43596
rect 22866 43484 22876 43540
rect 22932 43484 25340 43540
rect 25396 43484 25406 43540
rect 29474 43484 29484 43540
rect 29540 43484 30492 43540
rect 30548 43484 30558 43540
rect 700 43260 980 43316
rect 0 43092 800 43120
rect 924 43092 980 43260
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 0 43036 980 43092
rect 0 43008 800 43036
rect 21970 42700 21980 42756
rect 22036 42700 26124 42756
rect 26180 42700 26190 42756
rect 28354 42700 28364 42756
rect 28420 42700 30492 42756
rect 30548 42700 30558 42756
rect 19842 42588 19852 42644
rect 19908 42588 23324 42644
rect 23380 42588 23390 42644
rect 1698 42476 1708 42532
rect 1764 42476 1774 42532
rect 20132 42476 20188 42588
rect 20244 42476 20254 42532
rect 20402 42476 20412 42532
rect 20468 42476 25676 42532
rect 25732 42476 25742 42532
rect 28018 42476 28028 42532
rect 28084 42476 28364 42532
rect 28420 42476 28430 42532
rect 0 42420 800 42448
rect 1708 42420 1764 42476
rect 0 42364 1764 42420
rect 0 42336 800 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 20412 42196 20468 42476
rect 47200 42420 48000 42448
rect 46162 42364 46172 42420
rect 46228 42364 48000 42420
rect 47200 42336 48000 42364
rect 19506 42140 19516 42196
rect 19572 42140 20468 42196
rect 13570 42028 13580 42084
rect 13636 42028 17388 42084
rect 17444 42028 17454 42084
rect 22082 42028 22092 42084
rect 22148 42028 22428 42084
rect 22484 42028 23436 42084
rect 23492 42028 25564 42084
rect 25620 42028 26908 42084
rect 26964 42028 26974 42084
rect 31714 42028 31724 42084
rect 31780 42028 33516 42084
rect 33572 42028 33582 42084
rect 24098 41916 24108 41972
rect 24164 41916 25788 41972
rect 25844 41916 26460 41972
rect 26516 41916 26526 41972
rect 28690 41916 28700 41972
rect 28756 41916 30044 41972
rect 30100 41916 32508 41972
rect 32564 41916 33628 41972
rect 33684 41916 33694 41972
rect 16034 41804 16044 41860
rect 16100 41804 17948 41860
rect 18004 41804 18014 41860
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 25554 41356 25564 41412
rect 25620 41356 27244 41412
rect 27300 41356 27310 41412
rect 13682 41132 13692 41188
rect 13748 41132 18508 41188
rect 18564 41132 19404 41188
rect 19460 41132 19628 41188
rect 19684 41132 19694 41188
rect 27122 41132 27132 41188
rect 27188 41132 29484 41188
rect 29540 41132 29550 41188
rect 29922 41132 29932 41188
rect 29988 41132 31724 41188
rect 31780 41132 31790 41188
rect 20738 41020 20748 41076
rect 20804 41020 22876 41076
rect 22932 41020 22942 41076
rect 28466 41020 28476 41076
rect 28532 41020 30604 41076
rect 30660 41020 30670 41076
rect 23986 40908 23996 40964
rect 24052 40908 30156 40964
rect 30212 40908 30222 40964
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 17938 40684 17948 40740
rect 18004 40684 19628 40740
rect 19684 40684 19694 40740
rect 11890 40572 11900 40628
rect 11956 40572 16044 40628
rect 16100 40572 21308 40628
rect 21364 40572 21374 40628
rect 28242 40572 28252 40628
rect 28308 40572 31724 40628
rect 31780 40572 35084 40628
rect 35140 40572 35150 40628
rect 15138 40460 15148 40516
rect 15204 40460 16492 40516
rect 16548 40460 16558 40516
rect 22754 40460 22764 40516
rect 22820 40460 27132 40516
rect 27188 40460 27198 40516
rect 30482 40460 30492 40516
rect 30548 40460 31948 40516
rect 31892 40404 31948 40460
rect 12898 40348 12908 40404
rect 12964 40348 13692 40404
rect 13748 40348 14588 40404
rect 14644 40348 17388 40404
rect 17444 40348 17454 40404
rect 20626 40348 20636 40404
rect 20692 40348 21644 40404
rect 21700 40348 23884 40404
rect 23940 40348 23950 40404
rect 25442 40348 25452 40404
rect 25508 40348 28476 40404
rect 28532 40348 28542 40404
rect 29698 40348 29708 40404
rect 29764 40348 31276 40404
rect 31332 40348 31342 40404
rect 31892 40348 35532 40404
rect 35588 40348 35598 40404
rect 16156 40292 16212 40348
rect 11442 40236 11452 40292
rect 11508 40236 12796 40292
rect 12852 40236 12862 40292
rect 13458 40236 13468 40292
rect 13524 40236 15036 40292
rect 15092 40236 15932 40292
rect 15988 40236 15998 40292
rect 16146 40236 16156 40292
rect 16212 40236 16222 40292
rect 12114 40124 12124 40180
rect 12180 40124 14364 40180
rect 14420 40124 14430 40180
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 32274 39788 32284 39844
rect 32340 39788 34188 39844
rect 34244 39788 34254 39844
rect 19170 39676 19180 39732
rect 19236 39676 22092 39732
rect 22148 39676 27356 39732
rect 27412 39676 27422 39732
rect 14354 39564 14364 39620
rect 14420 39564 15596 39620
rect 15652 39564 15662 39620
rect 17490 39564 17500 39620
rect 17556 39564 19404 39620
rect 19460 39564 19470 39620
rect 27570 39564 27580 39620
rect 27636 39564 29708 39620
rect 29764 39564 30044 39620
rect 30100 39564 30110 39620
rect 15362 39452 15372 39508
rect 15428 39452 27692 39508
rect 27748 39452 29372 39508
rect 29428 39452 29438 39508
rect 7634 39340 7644 39396
rect 7700 39340 15260 39396
rect 15316 39340 21756 39396
rect 21812 39340 21822 39396
rect 22194 39340 22204 39396
rect 22260 39340 29148 39396
rect 29204 39340 29214 39396
rect 33170 39340 33180 39396
rect 33236 39340 34748 39396
rect 34804 39340 34814 39396
rect 12898 39228 12908 39284
rect 12964 39228 13692 39284
rect 13748 39228 13758 39284
rect 28018 39228 28028 39284
rect 28084 39228 33068 39284
rect 33124 39228 33134 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 11218 39004 11228 39060
rect 11284 39004 20188 39060
rect 37762 39004 37772 39060
rect 37828 39004 39452 39060
rect 39508 39004 39518 39060
rect 20132 38948 20188 39004
rect 9202 38892 9212 38948
rect 9268 38892 11676 38948
rect 11732 38892 12572 38948
rect 12628 38892 13468 38948
rect 13524 38892 13534 38948
rect 14354 38892 14364 38948
rect 14420 38892 15372 38948
rect 15428 38892 16716 38948
rect 16772 38892 16782 38948
rect 20132 38892 20972 38948
rect 21028 38892 21038 38948
rect 30706 38892 30716 38948
rect 30772 38892 36316 38948
rect 36372 38892 36382 38948
rect 15026 38780 15036 38836
rect 15092 38780 15484 38836
rect 15540 38780 16268 38836
rect 16324 38780 16828 38836
rect 16884 38780 16894 38836
rect 17826 38780 17836 38836
rect 17892 38780 22204 38836
rect 22260 38780 22270 38836
rect 32498 38780 32508 38836
rect 32564 38780 33516 38836
rect 33572 38780 33582 38836
rect 37650 38780 37660 38836
rect 37716 38780 38556 38836
rect 38612 38780 38892 38836
rect 38948 38780 38958 38836
rect 39666 38780 39676 38836
rect 39732 38780 39742 38836
rect 39676 38724 39732 38780
rect 13794 38668 13804 38724
rect 13860 38668 17388 38724
rect 17444 38668 17454 38724
rect 24098 38668 24108 38724
rect 24164 38668 25452 38724
rect 25508 38668 25518 38724
rect 30034 38668 30044 38724
rect 30100 38668 39732 38724
rect 29250 38556 29260 38612
rect 29316 38556 30828 38612
rect 30884 38556 32284 38612
rect 32340 38556 32350 38612
rect 38546 38556 38556 38612
rect 38612 38556 39228 38612
rect 39284 38556 40908 38612
rect 40964 38556 40974 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 16482 38220 16492 38276
rect 16548 38220 19068 38276
rect 19124 38220 22428 38276
rect 22484 38220 22494 38276
rect 23762 38220 23772 38276
rect 23828 38220 24556 38276
rect 24612 38220 26236 38276
rect 26292 38220 26302 38276
rect 19170 38108 19180 38164
rect 19236 38108 20188 38164
rect 20244 38108 24052 38164
rect 12786 37996 12796 38052
rect 12852 37996 15596 38052
rect 15652 37996 15662 38052
rect 18834 37996 18844 38052
rect 18900 37996 22988 38052
rect 23044 37996 23054 38052
rect 23996 37940 24052 38108
rect 39442 37996 39452 38052
rect 39508 37996 40908 38052
rect 40964 37996 40974 38052
rect 15092 37884 21308 37940
rect 21364 37884 21374 37940
rect 23986 37884 23996 37940
rect 24052 37884 24062 37940
rect 25890 37884 25900 37940
rect 25956 37884 27804 37940
rect 27860 37884 27870 37940
rect 36082 37884 36092 37940
rect 36148 37884 36988 37940
rect 37044 37884 37054 37940
rect 15092 37828 15148 37884
rect 14700 37772 15148 37828
rect 19842 37772 19852 37828
rect 19908 37772 21644 37828
rect 21700 37772 21710 37828
rect 23426 37772 23436 37828
rect 23492 37772 24220 37828
rect 24276 37772 24286 37828
rect 24546 37772 24556 37828
rect 24612 37772 25228 37828
rect 25284 37772 26572 37828
rect 26628 37772 26638 37828
rect 14700 37492 14756 37772
rect 24220 37716 24276 37772
rect 24220 37660 26124 37716
rect 26180 37660 26190 37716
rect 37426 37660 37436 37716
rect 37492 37660 38444 37716
rect 38500 37660 38510 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 13010 37436 13020 37492
rect 13076 37436 14252 37492
rect 14308 37436 14700 37492
rect 14756 37436 14766 37492
rect 21634 37436 21644 37492
rect 21700 37436 25788 37492
rect 25844 37436 25854 37492
rect 15138 37324 15148 37380
rect 15204 37324 17724 37380
rect 17780 37324 20412 37380
rect 20468 37324 20478 37380
rect 31266 37324 31276 37380
rect 31332 37324 32396 37380
rect 32452 37324 33516 37380
rect 33572 37324 33582 37380
rect 36082 37324 36092 37380
rect 36148 37324 37548 37380
rect 37604 37324 41244 37380
rect 41300 37324 41310 37380
rect 14578 37212 14588 37268
rect 14644 37212 15708 37268
rect 15764 37212 15774 37268
rect 16370 37212 16380 37268
rect 16436 37212 17836 37268
rect 17892 37212 17902 37268
rect 23986 37212 23996 37268
rect 24052 37212 25452 37268
rect 25508 37212 26460 37268
rect 26516 37212 26526 37268
rect 37090 37212 37100 37268
rect 37156 37212 39844 37268
rect 40002 37212 40012 37268
rect 40068 37212 41356 37268
rect 41412 37212 41422 37268
rect 44146 37212 44156 37268
rect 44212 37212 44222 37268
rect 39788 37156 39844 37212
rect 40684 37156 40740 37212
rect 16594 37100 16604 37156
rect 16660 37100 17388 37156
rect 17444 37100 17454 37156
rect 20066 37100 20076 37156
rect 20132 37100 21084 37156
rect 21140 37100 21150 37156
rect 24434 37100 24444 37156
rect 24500 37100 25340 37156
rect 25396 37100 27132 37156
rect 27188 37100 27198 37156
rect 30930 37100 30940 37156
rect 30996 37100 31612 37156
rect 31668 37100 35420 37156
rect 35476 37100 35980 37156
rect 36036 37100 36046 37156
rect 37426 37100 37436 37156
rect 37492 37100 38108 37156
rect 38164 37100 38892 37156
rect 38948 37100 39228 37156
rect 39284 37100 39294 37156
rect 39788 37100 40348 37156
rect 40404 37100 40414 37156
rect 40674 37100 40684 37156
rect 40740 37100 40750 37156
rect 42018 37100 42028 37156
rect 42084 37100 43820 37156
rect 43876 37100 43886 37156
rect 44156 37044 44212 37212
rect 15026 36988 15036 37044
rect 15092 36876 15148 37044
rect 15250 36988 15260 37044
rect 15316 36988 16268 37044
rect 16324 36988 16492 37044
rect 16548 36988 16558 37044
rect 19618 36988 19628 37044
rect 19684 36988 21308 37044
rect 21364 36988 21476 37044
rect 22306 36988 22316 37044
rect 22372 36988 23548 37044
rect 23604 36988 24556 37044
rect 24612 36988 24622 37044
rect 33954 36988 33964 37044
rect 34020 36988 34860 37044
rect 34916 36988 35868 37044
rect 35924 36988 36484 37044
rect 36642 36988 36652 37044
rect 36708 36988 37100 37044
rect 37156 36988 37996 37044
rect 38052 36988 38556 37044
rect 38612 36988 39564 37044
rect 39620 36988 39630 37044
rect 40450 36988 40460 37044
rect 40516 36988 41356 37044
rect 41412 36988 41422 37044
rect 43362 36988 43372 37044
rect 43428 36988 44212 37044
rect 21420 36932 21476 36988
rect 36428 36932 36484 36988
rect 15204 36876 15214 36932
rect 21420 36876 22092 36932
rect 22148 36876 22158 36932
rect 22754 36876 22764 36932
rect 22820 36876 26348 36932
rect 26404 36876 29372 36932
rect 29428 36876 29438 36932
rect 36428 36876 42364 36932
rect 42420 36876 42430 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 15810 36764 15820 36820
rect 15876 36764 17612 36820
rect 17668 36764 17678 36820
rect 24098 36652 24108 36708
rect 24164 36652 27692 36708
rect 27748 36652 27758 36708
rect 13682 36540 13692 36596
rect 13748 36540 15484 36596
rect 15540 36540 15550 36596
rect 25666 36540 25676 36596
rect 25732 36540 26908 36596
rect 39330 36540 39340 36596
rect 39396 36540 42476 36596
rect 42532 36540 43036 36596
rect 43092 36540 43102 36596
rect 26852 36484 26908 36540
rect 9426 36428 9436 36484
rect 9492 36428 11116 36484
rect 11172 36428 11182 36484
rect 19730 36428 19740 36484
rect 19796 36428 21644 36484
rect 21700 36428 24892 36484
rect 24948 36428 24958 36484
rect 26852 36428 30604 36484
rect 30660 36428 30670 36484
rect 34178 36428 34188 36484
rect 34244 36428 36204 36484
rect 36260 36428 36270 36484
rect 38210 36428 38220 36484
rect 38276 36428 39788 36484
rect 39844 36428 42700 36484
rect 42756 36428 43484 36484
rect 43540 36428 43708 36484
rect 43652 36372 43708 36428
rect 2034 36316 2044 36372
rect 2100 36316 6300 36372
rect 6356 36316 6366 36372
rect 9650 36316 9660 36372
rect 9716 36316 10108 36372
rect 10164 36316 10892 36372
rect 10948 36316 15260 36372
rect 15316 36316 15326 36372
rect 19506 36316 19516 36372
rect 19572 36316 21868 36372
rect 21924 36316 21934 36372
rect 22082 36316 22092 36372
rect 22148 36316 22428 36372
rect 22484 36316 22494 36372
rect 28466 36316 28476 36372
rect 28532 36316 29148 36372
rect 29204 36316 29214 36372
rect 37650 36316 37660 36372
rect 37716 36316 38108 36372
rect 38164 36316 38174 36372
rect 43652 36316 44828 36372
rect 44884 36316 44894 36372
rect 5506 36204 5516 36260
rect 5572 36204 6972 36260
rect 7028 36204 7038 36260
rect 10770 36204 10780 36260
rect 10836 36204 11228 36260
rect 11284 36204 15372 36260
rect 15428 36204 15438 36260
rect 22530 36204 22540 36260
rect 22596 36204 22876 36260
rect 22932 36204 22942 36260
rect 26674 36204 26684 36260
rect 26740 36204 30156 36260
rect 30212 36204 30222 36260
rect 37538 36204 37548 36260
rect 37604 36204 40124 36260
rect 40180 36204 41356 36260
rect 41412 36204 41422 36260
rect 5170 36092 5180 36148
rect 5236 36092 5964 36148
rect 6020 36092 6748 36148
rect 6804 36092 7980 36148
rect 8036 36092 8046 36148
rect 12898 36092 12908 36148
rect 12964 36092 16492 36148
rect 16548 36092 16558 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 14354 35980 14364 36036
rect 14420 35980 16604 36036
rect 16660 35980 16670 36036
rect 27794 35980 27804 36036
rect 27860 35980 28588 36036
rect 28644 35980 39900 36036
rect 39956 35980 39966 36036
rect 4834 35868 4844 35924
rect 4900 35868 6748 35924
rect 6804 35868 6814 35924
rect 41906 35868 41916 35924
rect 41972 35868 43036 35924
rect 43092 35868 44940 35924
rect 44996 35868 45006 35924
rect 22194 35756 22204 35812
rect 22260 35756 23548 35812
rect 23604 35756 23614 35812
rect 3154 35644 3164 35700
rect 3220 35644 3836 35700
rect 3892 35644 3902 35700
rect 4498 35644 4508 35700
rect 4564 35644 5516 35700
rect 5572 35644 5582 35700
rect 20402 35644 20412 35700
rect 20468 35644 21532 35700
rect 21588 35644 21598 35700
rect 5618 35532 5628 35588
rect 5684 35532 8540 35588
rect 8596 35532 8606 35588
rect 3490 35420 3500 35476
rect 3556 35420 4900 35476
rect 6178 35420 6188 35476
rect 6244 35420 7756 35476
rect 7812 35420 7822 35476
rect 15586 35420 15596 35476
rect 15652 35420 18284 35476
rect 18340 35420 18350 35476
rect 22866 35420 22876 35476
rect 22932 35420 24332 35476
rect 24388 35420 24398 35476
rect 25554 35420 25564 35476
rect 25620 35420 27020 35476
rect 27076 35420 27086 35476
rect 41458 35420 41468 35476
rect 41524 35420 43260 35476
rect 43316 35420 43326 35476
rect 4844 35364 4900 35420
rect 4844 35308 8204 35364
rect 8260 35308 8270 35364
rect 27570 35308 27580 35364
rect 27636 35308 28252 35364
rect 28308 35308 34300 35364
rect 34356 35308 34366 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 30156 35252 30212 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 22194 35196 22204 35252
rect 22260 35196 22876 35252
rect 22932 35196 22942 35252
rect 27122 35196 27132 35252
rect 27188 35196 29148 35252
rect 29204 35196 29214 35252
rect 30146 35196 30156 35252
rect 30212 35196 30222 35252
rect 38658 35196 38668 35252
rect 38724 35196 39788 35252
rect 39844 35196 39854 35252
rect 4946 35084 4956 35140
rect 5012 35084 6076 35140
rect 6132 35084 6142 35140
rect 7858 35084 7868 35140
rect 7924 35084 9212 35140
rect 9268 35084 9278 35140
rect 14578 35084 14588 35140
rect 14644 35084 15148 35140
rect 33618 35084 33628 35140
rect 33684 35084 39452 35140
rect 39508 35084 39518 35140
rect 3042 34972 3052 35028
rect 3108 34972 5404 35028
rect 5460 34972 5470 35028
rect 13010 34972 13020 35028
rect 13076 34972 14476 35028
rect 14532 34972 14542 35028
rect 15092 34916 15148 35084
rect 22614 34972 22652 35028
rect 22708 34972 22718 35028
rect 26338 34972 26348 35028
rect 26404 34972 26572 35028
rect 26628 34972 26638 35028
rect 15092 34860 15372 34916
rect 15428 34860 15438 34916
rect 34738 34860 34748 34916
rect 34804 34860 38668 34916
rect 38724 34860 38734 34916
rect 8194 34748 8204 34804
rect 8260 34748 8540 34804
rect 8596 34748 9884 34804
rect 9940 34748 9950 34804
rect 37650 34748 37660 34804
rect 37716 34748 39676 34804
rect 39732 34748 39742 34804
rect 40002 34748 40012 34804
rect 40068 34748 41412 34804
rect 41570 34748 41580 34804
rect 41636 34748 44044 34804
rect 44100 34748 44110 34804
rect 45154 34748 45164 34804
rect 45220 34748 45230 34804
rect 41356 34692 41412 34748
rect 45164 34692 45220 34748
rect 4386 34636 4396 34692
rect 4452 34636 5068 34692
rect 5124 34636 5964 34692
rect 6020 34636 8316 34692
rect 8372 34636 8382 34692
rect 20850 34636 20860 34692
rect 20916 34636 21756 34692
rect 21812 34636 21980 34692
rect 22036 34636 23772 34692
rect 23828 34636 23838 34692
rect 37090 34636 37100 34692
rect 37156 34636 39340 34692
rect 39396 34636 41132 34692
rect 41188 34636 41198 34692
rect 41356 34636 45220 34692
rect 22082 34524 22092 34580
rect 22148 34524 23212 34580
rect 23268 34524 23278 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 35746 34412 35756 34468
rect 35812 34412 37212 34468
rect 37268 34412 42700 34468
rect 42756 34412 42766 34468
rect 0 34356 800 34384
rect 0 34300 1708 34356
rect 1764 34300 2492 34356
rect 2548 34300 2558 34356
rect 39442 34300 39452 34356
rect 39508 34300 40460 34356
rect 40516 34300 40526 34356
rect 0 34272 800 34300
rect 15586 34188 15596 34244
rect 15652 34188 16156 34244
rect 16212 34188 16828 34244
rect 16884 34188 16894 34244
rect 22418 34188 22428 34244
rect 22484 34188 22652 34244
rect 22708 34188 23660 34244
rect 23716 34188 25228 34244
rect 25284 34188 25294 34244
rect 39106 34188 39116 34244
rect 39172 34188 43708 34244
rect 43652 34132 43708 34188
rect 17490 34076 17500 34132
rect 17556 34076 18172 34132
rect 18228 34076 19292 34132
rect 19348 34076 19358 34132
rect 37426 34076 37436 34132
rect 37492 34076 39004 34132
rect 39060 34076 39070 34132
rect 39778 34076 39788 34132
rect 39844 34076 40908 34132
rect 40964 34076 40974 34132
rect 43652 34076 45388 34132
rect 45444 34076 45454 34132
rect 36978 33964 36988 34020
rect 37044 33964 37996 34020
rect 38052 33964 38062 34020
rect 38612 33964 38892 34020
rect 38948 33964 38958 34020
rect 44034 33964 44044 34020
rect 44100 33964 44828 34020
rect 44884 33964 44894 34020
rect 38612 33908 38668 33964
rect 4274 33852 4284 33908
rect 4340 33852 5292 33908
rect 5348 33852 5358 33908
rect 6066 33852 6076 33908
rect 6132 33852 6636 33908
rect 6692 33852 9548 33908
rect 9604 33852 9614 33908
rect 19282 33852 19292 33908
rect 19348 33852 23212 33908
rect 23268 33852 26348 33908
rect 26404 33852 26414 33908
rect 38098 33852 38108 33908
rect 38164 33852 38332 33908
rect 38388 33852 38668 33908
rect 44146 33852 44156 33908
rect 44212 33852 45948 33908
rect 46004 33852 46014 33908
rect 28018 33740 28028 33796
rect 28084 33740 29484 33796
rect 29540 33740 29550 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 16034 33628 16044 33684
rect 16100 33628 17612 33684
rect 17668 33628 21868 33684
rect 21924 33628 22652 33684
rect 22708 33628 22718 33684
rect 24434 33628 24444 33684
rect 24500 33628 25508 33684
rect 37202 33628 37212 33684
rect 37268 33628 38108 33684
rect 38164 33628 38174 33684
rect 25452 33572 25508 33628
rect 2146 33516 2156 33572
rect 2212 33516 4172 33572
rect 4228 33516 4238 33572
rect 12786 33516 12796 33572
rect 12852 33516 15820 33572
rect 15876 33516 16940 33572
rect 16996 33516 17006 33572
rect 25452 33516 25564 33572
rect 25620 33516 25630 33572
rect 4050 33404 4060 33460
rect 4116 33404 6188 33460
rect 6244 33404 10556 33460
rect 10612 33404 10622 33460
rect 11330 33404 11340 33460
rect 11396 33404 13356 33460
rect 13412 33404 13916 33460
rect 13972 33404 14924 33460
rect 14980 33404 14990 33460
rect 23986 33404 23996 33460
rect 24052 33404 25676 33460
rect 25732 33404 25742 33460
rect 28578 33404 28588 33460
rect 28644 33404 29260 33460
rect 29316 33404 29326 33460
rect 4834 33292 4844 33348
rect 4900 33292 5628 33348
rect 5684 33292 5694 33348
rect 15026 33292 15036 33348
rect 15092 33292 17276 33348
rect 17332 33292 17342 33348
rect 21634 33292 21644 33348
rect 21700 33292 22428 33348
rect 22484 33292 25228 33348
rect 25284 33292 25294 33348
rect 29698 33292 29708 33348
rect 29764 33292 32060 33348
rect 32116 33292 32956 33348
rect 33012 33292 33022 33348
rect 38658 33292 38668 33348
rect 38724 33292 39116 33348
rect 39172 33292 42700 33348
rect 42756 33292 42766 33348
rect 2034 33180 2044 33236
rect 2100 33180 3724 33236
rect 3780 33180 3790 33236
rect 9538 33180 9548 33236
rect 9604 33180 10332 33236
rect 10388 33180 10398 33236
rect 21410 33180 21420 33236
rect 21476 33180 22204 33236
rect 22260 33180 22270 33236
rect 26562 33180 26572 33236
rect 26628 33180 28252 33236
rect 28308 33180 29036 33236
rect 29092 33180 29102 33236
rect 8642 33068 8652 33124
rect 8708 33068 10108 33124
rect 10164 33068 10174 33124
rect 22754 33068 22764 33124
rect 22820 33068 23324 33124
rect 23380 33068 23390 33124
rect 24546 33068 24556 33124
rect 24612 33068 25452 33124
rect 25508 33068 26348 33124
rect 26404 33068 26414 33124
rect 28690 33068 28700 33124
rect 28756 33068 29372 33124
rect 29428 33068 29438 33124
rect 37650 33068 37660 33124
rect 37716 33068 38220 33124
rect 38276 33068 45836 33124
rect 45892 33068 45902 33124
rect 3714 32956 3724 33012
rect 3780 32956 4844 33012
rect 4900 32956 4910 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 14466 32844 14476 32900
rect 14532 32844 16156 32900
rect 16212 32844 16222 32900
rect 3826 32732 3836 32788
rect 3892 32732 5404 32788
rect 5460 32732 5470 32788
rect 6962 32732 6972 32788
rect 7028 32732 8540 32788
rect 8596 32732 8606 32788
rect 11666 32620 11676 32676
rect 11732 32620 22204 32676
rect 22260 32620 22270 32676
rect 12562 32508 12572 32564
rect 12628 32508 13692 32564
rect 13748 32508 14700 32564
rect 14756 32508 14766 32564
rect 20290 32508 20300 32564
rect 20356 32508 21420 32564
rect 21476 32508 21486 32564
rect 24434 32508 24444 32564
rect 24500 32508 25900 32564
rect 25956 32508 25966 32564
rect 26852 32508 28028 32564
rect 28084 32508 28094 32564
rect 32386 32508 32396 32564
rect 32452 32508 33516 32564
rect 33572 32508 33582 32564
rect 36754 32508 36764 32564
rect 36820 32508 38332 32564
rect 38388 32508 39564 32564
rect 39620 32508 39630 32564
rect 26852 32452 26908 32508
rect 10546 32396 10556 32452
rect 10612 32396 11564 32452
rect 11620 32396 12012 32452
rect 12068 32396 12078 32452
rect 19282 32396 19292 32452
rect 19348 32396 20412 32452
rect 20468 32396 20478 32452
rect 25554 32396 25564 32452
rect 25620 32396 26908 32452
rect 27010 32396 27020 32452
rect 27076 32396 27086 32452
rect 32610 32396 32620 32452
rect 32676 32396 36428 32452
rect 36484 32396 36494 32452
rect 36978 32396 36988 32452
rect 37044 32396 38892 32452
rect 38948 32396 38958 32452
rect 16930 32284 16940 32340
rect 16996 32284 22204 32340
rect 22260 32284 22270 32340
rect 12898 32172 12908 32228
rect 12964 32172 13580 32228
rect 13636 32172 17276 32228
rect 17332 32172 17342 32228
rect 20402 32172 20412 32228
rect 20468 32172 21644 32228
rect 21700 32172 21710 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 21186 32060 21196 32116
rect 21252 32060 25340 32116
rect 25396 32060 25406 32116
rect 13682 31948 13692 32004
rect 13748 31948 15036 32004
rect 15092 31948 15102 32004
rect 18722 31948 18732 32004
rect 18788 31948 20972 32004
rect 21028 31948 21038 32004
rect 16594 31836 16604 31892
rect 16660 31836 19404 31892
rect 19460 31836 19908 31892
rect 19852 31780 19908 31836
rect 21756 31780 21812 32060
rect 27020 32004 27076 32396
rect 34290 32284 34300 32340
rect 34356 32284 38780 32340
rect 38836 32284 38846 32340
rect 43250 32284 43260 32340
rect 43316 32284 43932 32340
rect 43988 32284 45164 32340
rect 45220 32284 45230 32340
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 36418 32060 36428 32116
rect 36484 32060 36932 32116
rect 36876 32004 36932 32060
rect 27010 31948 27020 32004
rect 27076 31948 27086 32004
rect 27234 31948 27244 32004
rect 27300 31948 28700 32004
rect 28756 31948 28766 32004
rect 36876 31948 38668 32004
rect 38612 31892 38668 31948
rect 22082 31836 22092 31892
rect 22148 31836 22158 31892
rect 27794 31836 27804 31892
rect 27860 31836 29260 31892
rect 29316 31836 29326 31892
rect 35746 31836 35756 31892
rect 35812 31836 36540 31892
rect 36596 31836 36606 31892
rect 37538 31836 37548 31892
rect 37604 31836 37614 31892
rect 38612 31836 41580 31892
rect 41636 31836 41646 31892
rect 43652 31836 45612 31892
rect 45668 31836 45678 31892
rect 11554 31724 11564 31780
rect 11620 31724 12236 31780
rect 12292 31724 12302 31780
rect 17602 31724 17612 31780
rect 17668 31724 18956 31780
rect 19012 31724 19022 31780
rect 19842 31724 19852 31780
rect 19908 31724 21756 31780
rect 21812 31724 21822 31780
rect 22092 31668 22148 31836
rect 23426 31724 23436 31780
rect 23492 31724 25228 31780
rect 25284 31724 25294 31780
rect 28354 31724 28364 31780
rect 28420 31724 29596 31780
rect 29652 31724 30268 31780
rect 30324 31724 30334 31780
rect 3938 31612 3948 31668
rect 4004 31612 5516 31668
rect 5572 31612 5582 31668
rect 11218 31612 11228 31668
rect 11284 31612 11900 31668
rect 11956 31612 13580 31668
rect 13636 31612 13646 31668
rect 15362 31612 15372 31668
rect 15428 31612 17948 31668
rect 18004 31612 18014 31668
rect 21634 31612 21644 31668
rect 21700 31612 22148 31668
rect 37548 31668 37604 31836
rect 43652 31780 43708 31836
rect 37874 31724 37884 31780
rect 37940 31724 39452 31780
rect 39508 31724 42700 31780
rect 42756 31724 43708 31780
rect 37548 31612 39004 31668
rect 39060 31612 39070 31668
rect 2482 31500 2492 31556
rect 2548 31500 3836 31556
rect 3892 31500 3902 31556
rect 8306 31500 8316 31556
rect 8372 31500 9212 31556
rect 9268 31500 10444 31556
rect 10500 31500 10510 31556
rect 14466 31500 14476 31556
rect 14532 31500 15148 31556
rect 25554 31500 25564 31556
rect 25620 31500 26124 31556
rect 26180 31500 26190 31556
rect 27570 31500 27580 31556
rect 27636 31500 29484 31556
rect 29540 31500 39564 31556
rect 39620 31500 40236 31556
rect 40292 31500 43708 31556
rect 15092 31332 15148 31500
rect 43652 31444 43708 31500
rect 26786 31388 26796 31444
rect 26852 31388 29372 31444
rect 29428 31388 30828 31444
rect 30884 31388 30894 31444
rect 43652 31388 44940 31444
rect 44996 31388 45006 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 15092 31276 15372 31332
rect 15428 31276 15438 31332
rect 36530 31276 36540 31332
rect 36596 31276 37324 31332
rect 37380 31276 37390 31332
rect 7410 31164 7420 31220
rect 7476 31164 8204 31220
rect 8260 31164 8270 31220
rect 20738 31164 20748 31220
rect 20804 31164 22540 31220
rect 22596 31164 24108 31220
rect 24164 31164 24174 31220
rect 25554 31164 25564 31220
rect 25620 31164 26684 31220
rect 26740 31164 26750 31220
rect 15026 31052 15036 31108
rect 15092 31052 15708 31108
rect 15764 31052 16828 31108
rect 16884 31052 16894 31108
rect 28018 31052 28028 31108
rect 28084 31052 28812 31108
rect 28868 31052 28878 31108
rect 34626 31052 34636 31108
rect 34692 31052 37548 31108
rect 37604 31052 37614 31108
rect 12226 30940 12236 30996
rect 12292 30940 16044 30996
rect 16100 30940 16110 30996
rect 37548 30884 37604 31052
rect 38210 30940 38220 30996
rect 38276 30940 42028 30996
rect 42084 30940 42094 30996
rect 16370 30828 16380 30884
rect 16436 30828 17612 30884
rect 17668 30828 17678 30884
rect 24322 30828 24332 30884
rect 24388 30828 25228 30884
rect 25284 30828 25294 30884
rect 35522 30828 35532 30884
rect 35588 30828 36092 30884
rect 36148 30828 36158 30884
rect 36866 30828 36876 30884
rect 36932 30828 37324 30884
rect 37380 30828 37390 30884
rect 37548 30828 41692 30884
rect 41748 30828 41758 30884
rect 44930 30828 44940 30884
rect 44996 30828 45724 30884
rect 45780 30828 45790 30884
rect 44818 30716 44828 30772
rect 44884 30716 45164 30772
rect 45220 30716 45230 30772
rect 21970 30604 21980 30660
rect 22036 30604 22428 30660
rect 22484 30604 26572 30660
rect 26628 30604 26638 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 36754 30380 36764 30436
rect 36820 30380 38108 30436
rect 38164 30380 38174 30436
rect 43474 30380 43484 30436
rect 43540 30380 45500 30436
rect 45556 30380 45566 30436
rect 25330 30268 25340 30324
rect 25396 30268 26348 30324
rect 26404 30268 26796 30324
rect 26852 30268 26862 30324
rect 43250 30268 43260 30324
rect 43316 30268 44828 30324
rect 44884 30268 44894 30324
rect 2258 30156 2268 30212
rect 2324 30156 3724 30212
rect 3780 30156 3790 30212
rect 10770 30156 10780 30212
rect 10836 30156 12124 30212
rect 12180 30156 13356 30212
rect 13412 30156 13422 30212
rect 15474 30156 15484 30212
rect 15540 30156 17388 30212
rect 17444 30156 17454 30212
rect 19506 30156 19516 30212
rect 19572 30156 20188 30212
rect 20244 30156 20254 30212
rect 22082 30156 22092 30212
rect 22148 30156 22158 30212
rect 24546 30156 24556 30212
rect 24612 30156 25788 30212
rect 25844 30156 25854 30212
rect 27122 30156 27132 30212
rect 27188 30156 27692 30212
rect 27748 30156 27758 30212
rect 28354 30156 28364 30212
rect 28420 30156 29148 30212
rect 29204 30156 29214 30212
rect 37314 30156 37324 30212
rect 37380 30156 37884 30212
rect 37940 30156 37950 30212
rect 41458 30156 41468 30212
rect 41524 30156 42140 30212
rect 42196 30156 42206 30212
rect 43586 30156 43596 30212
rect 43652 30156 44268 30212
rect 44324 30156 44334 30212
rect 22092 30100 22148 30156
rect 3826 30044 3836 30100
rect 3892 30044 5404 30100
rect 5460 30044 5470 30100
rect 12786 30044 12796 30100
rect 12852 30044 13468 30100
rect 13524 30044 15820 30100
rect 15876 30044 15886 30100
rect 22092 30044 26908 30100
rect 34738 30044 34748 30100
rect 34804 30044 35756 30100
rect 35812 30044 35822 30100
rect 38882 30044 38892 30100
rect 38948 30044 41020 30100
rect 41076 30044 45388 30100
rect 45444 30044 45454 30100
rect 17826 29932 17836 29988
rect 17892 29932 19628 29988
rect 19684 29932 19694 29988
rect 21746 29932 21756 29988
rect 21812 29932 22540 29988
rect 22596 29932 22606 29988
rect 23090 29820 23100 29876
rect 23156 29820 24332 29876
rect 24388 29820 25788 29876
rect 25844 29820 25854 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 26852 29764 26908 30044
rect 28242 29932 28252 29988
rect 28308 29932 30604 29988
rect 30660 29932 33180 29988
rect 33236 29932 33246 29988
rect 20290 29708 20300 29764
rect 20356 29708 21196 29764
rect 21252 29708 23884 29764
rect 23940 29708 23950 29764
rect 26852 29708 28588 29764
rect 28644 29708 28654 29764
rect 5058 29596 5068 29652
rect 5124 29596 5628 29652
rect 5684 29596 5694 29652
rect 14914 29596 14924 29652
rect 14980 29596 16492 29652
rect 16548 29596 16558 29652
rect 17714 29596 17724 29652
rect 17780 29596 33068 29652
rect 33124 29596 33134 29652
rect 34738 29596 34748 29652
rect 34804 29596 35532 29652
rect 35588 29596 35598 29652
rect 38882 29596 38892 29652
rect 38948 29596 39900 29652
rect 39956 29596 42812 29652
rect 42868 29596 43372 29652
rect 43428 29596 43438 29652
rect 13906 29484 13916 29540
rect 13972 29484 15932 29540
rect 15988 29484 16716 29540
rect 16772 29484 16782 29540
rect 18498 29484 18508 29540
rect 18564 29484 22708 29540
rect 23650 29484 23660 29540
rect 23716 29484 24892 29540
rect 24948 29484 24958 29540
rect 25778 29484 25788 29540
rect 25844 29484 27804 29540
rect 27860 29484 27870 29540
rect 28466 29484 28476 29540
rect 28532 29484 30380 29540
rect 30436 29484 30446 29540
rect 32050 29484 32060 29540
rect 32116 29484 33516 29540
rect 33572 29484 33582 29540
rect 36306 29484 36316 29540
rect 36372 29484 38220 29540
rect 38276 29484 38286 29540
rect 41346 29484 41356 29540
rect 41412 29484 41804 29540
rect 41860 29484 43596 29540
rect 43652 29484 43662 29540
rect 22652 29428 22708 29484
rect 15092 29372 20860 29428
rect 20916 29372 20926 29428
rect 22642 29372 22652 29428
rect 22708 29372 22718 29428
rect 23426 29372 23436 29428
rect 23492 29372 24556 29428
rect 24612 29372 24622 29428
rect 29250 29372 29260 29428
rect 29316 29372 29932 29428
rect 29988 29372 34748 29428
rect 34804 29372 34814 29428
rect 37202 29372 37212 29428
rect 37268 29372 39340 29428
rect 39396 29372 39406 29428
rect 41010 29372 41020 29428
rect 41076 29372 43036 29428
rect 43092 29372 43102 29428
rect 15092 29316 15148 29372
rect 24556 29316 24612 29372
rect 14130 29260 14140 29316
rect 14196 29260 15148 29316
rect 19394 29260 19404 29316
rect 19460 29260 20188 29316
rect 20244 29260 20254 29316
rect 22306 29260 22316 29316
rect 22372 29260 23100 29316
rect 23156 29260 23166 29316
rect 24556 29260 25564 29316
rect 25620 29260 25630 29316
rect 44482 29260 44492 29316
rect 44548 29260 45948 29316
rect 46004 29260 46014 29316
rect 22978 29148 22988 29204
rect 23044 29148 23436 29204
rect 23492 29148 33404 29204
rect 33460 29148 33470 29204
rect 11666 29036 11676 29092
rect 11732 29036 14140 29092
rect 14196 29036 14206 29092
rect 14914 29036 14924 29092
rect 14980 29036 21980 29092
rect 22036 29036 22046 29092
rect 28578 29036 28588 29092
rect 28644 29036 33964 29092
rect 34020 29036 34860 29092
rect 34916 29036 34926 29092
rect 36418 29036 36428 29092
rect 36484 29036 37772 29092
rect 37828 29036 40796 29092
rect 40852 29036 42812 29092
rect 42868 29036 42878 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 28130 28924 28140 28980
rect 28196 28924 28924 28980
rect 28980 28924 31164 28980
rect 31220 28924 33628 28980
rect 33684 28924 33694 28980
rect 35532 28924 37100 28980
rect 37156 28924 37166 28980
rect 38994 28924 39004 28980
rect 39060 28924 41692 28980
rect 41748 28924 45612 28980
rect 45668 28924 45678 28980
rect 35532 28868 35588 28924
rect 26852 28812 35588 28868
rect 35858 28812 35868 28868
rect 35924 28812 36540 28868
rect 36596 28812 41468 28868
rect 41524 28812 41534 28868
rect 1810 28588 1820 28644
rect 1876 28588 2268 28644
rect 2324 28588 5628 28644
rect 5684 28588 5694 28644
rect 22306 28588 22316 28644
rect 22372 28588 23324 28644
rect 23380 28588 23884 28644
rect 23940 28588 23950 28644
rect 26852 28532 26908 28812
rect 28354 28700 28364 28756
rect 28420 28700 30548 28756
rect 32274 28700 32284 28756
rect 32340 28700 32956 28756
rect 33012 28700 33022 28756
rect 43698 28700 43708 28756
rect 43764 28700 44604 28756
rect 44660 28700 44670 28756
rect 30492 28644 30548 28700
rect 27682 28588 27692 28644
rect 27748 28588 29260 28644
rect 29316 28588 29326 28644
rect 30482 28588 30492 28644
rect 30548 28588 31836 28644
rect 31892 28588 32844 28644
rect 32900 28588 32910 28644
rect 33506 28588 33516 28644
rect 33572 28588 34524 28644
rect 34580 28588 34590 28644
rect 34748 28588 42924 28644
rect 42980 28588 42990 28644
rect 34748 28532 34804 28588
rect 10098 28476 10108 28532
rect 10164 28476 11452 28532
rect 11508 28476 11518 28532
rect 15810 28476 15820 28532
rect 15876 28476 16828 28532
rect 16884 28476 17388 28532
rect 17444 28476 17454 28532
rect 21298 28476 21308 28532
rect 21364 28476 24220 28532
rect 24276 28476 24286 28532
rect 25106 28476 25116 28532
rect 25172 28476 26908 28532
rect 32946 28476 32956 28532
rect 33012 28476 34804 28532
rect 34962 28476 34972 28532
rect 35028 28476 36316 28532
rect 36372 28476 36382 28532
rect 43922 28476 43932 28532
rect 43988 28476 44940 28532
rect 44996 28476 45006 28532
rect 9538 28364 9548 28420
rect 9604 28364 10444 28420
rect 10500 28364 10510 28420
rect 19954 28364 19964 28420
rect 20020 28364 20860 28420
rect 20916 28364 20926 28420
rect 21410 28364 21420 28420
rect 21476 28364 22092 28420
rect 22148 28364 22158 28420
rect 23426 28364 23436 28420
rect 23492 28364 24892 28420
rect 24948 28364 24958 28420
rect 43652 28252 43820 28308
rect 43876 28252 43886 28308
rect 44034 28252 44044 28308
rect 44100 28252 44828 28308
rect 44884 28252 44894 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 43652 28084 43708 28252
rect 4274 28028 4284 28084
rect 4340 28028 10220 28084
rect 10276 28028 10286 28084
rect 18274 28028 18284 28084
rect 18340 28028 20748 28084
rect 20804 28028 20814 28084
rect 23202 28028 23212 28084
rect 23268 28028 23996 28084
rect 24052 28028 24556 28084
rect 24612 28028 25340 28084
rect 25396 28028 25406 28084
rect 33394 28028 33404 28084
rect 33460 28028 33964 28084
rect 34020 28028 34300 28084
rect 34356 28028 34366 28084
rect 34738 28028 34748 28084
rect 34804 28028 38780 28084
rect 38836 28028 43708 28084
rect 4722 27916 4732 27972
rect 4788 27916 6636 27972
rect 6692 27916 6702 27972
rect 26114 27916 26124 27972
rect 26180 27916 27132 27972
rect 27188 27916 27198 27972
rect 28578 27916 28588 27972
rect 28644 27916 29820 27972
rect 29876 27916 34188 27972
rect 34244 27916 34254 27972
rect 16482 27804 16492 27860
rect 16548 27804 17500 27860
rect 17556 27804 19180 27860
rect 19236 27804 19246 27860
rect 21298 27804 21308 27860
rect 21364 27804 21644 27860
rect 21700 27804 21710 27860
rect 21970 27804 21980 27860
rect 22036 27804 23660 27860
rect 23716 27804 23726 27860
rect 29362 27804 29372 27860
rect 29428 27804 32172 27860
rect 32228 27804 32238 27860
rect 33058 27804 33068 27860
rect 33124 27804 34300 27860
rect 34356 27804 34366 27860
rect 37874 27804 37884 27860
rect 37940 27804 40012 27860
rect 40068 27804 41020 27860
rect 41076 27804 41086 27860
rect 17042 27692 17052 27748
rect 17108 27692 28700 27748
rect 28756 27692 28766 27748
rect 30034 27692 30044 27748
rect 30100 27692 31500 27748
rect 31556 27692 31566 27748
rect 39554 27692 39564 27748
rect 39620 27692 40684 27748
rect 40740 27692 40750 27748
rect 0 27636 800 27664
rect 0 27580 1932 27636
rect 1988 27580 1998 27636
rect 16594 27580 16604 27636
rect 16660 27580 18284 27636
rect 18340 27580 18350 27636
rect 18610 27580 18620 27636
rect 18676 27580 22204 27636
rect 22260 27580 22270 27636
rect 24210 27580 24220 27636
rect 24276 27580 24668 27636
rect 24724 27580 25004 27636
rect 25060 27580 25070 27636
rect 29138 27580 29148 27636
rect 29204 27580 38668 27636
rect 38724 27580 38734 27636
rect 0 27552 800 27580
rect 12338 27468 12348 27524
rect 12404 27468 32396 27524
rect 32452 27468 33852 27524
rect 33908 27468 33918 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 9874 27356 9884 27412
rect 9940 27356 13692 27412
rect 13748 27356 13758 27412
rect 19506 27356 19516 27412
rect 19572 27356 21532 27412
rect 21588 27356 24332 27412
rect 24388 27356 32172 27412
rect 32228 27356 32238 27412
rect 39330 27356 39340 27412
rect 39396 27356 43708 27412
rect 43764 27356 43774 27412
rect 13234 27244 13244 27300
rect 13300 27244 13804 27300
rect 13860 27244 14812 27300
rect 14868 27244 14878 27300
rect 18722 27244 18732 27300
rect 18788 27244 21756 27300
rect 21812 27244 21822 27300
rect 37426 27244 37436 27300
rect 37492 27244 37772 27300
rect 37828 27244 37838 27300
rect 1922 27132 1932 27188
rect 1988 27132 1998 27188
rect 12674 27132 12684 27188
rect 12740 27132 16492 27188
rect 16548 27132 16558 27188
rect 17490 27132 17500 27188
rect 17556 27132 22092 27188
rect 22148 27132 22158 27188
rect 25106 27132 25116 27188
rect 25172 27132 25182 27188
rect 30258 27132 30268 27188
rect 30324 27132 30716 27188
rect 30772 27132 30782 27188
rect 35186 27132 35196 27188
rect 35252 27132 40012 27188
rect 40068 27132 41244 27188
rect 41300 27132 41692 27188
rect 41748 27132 41758 27188
rect 0 26964 800 26992
rect 1932 26964 1988 27132
rect 25116 27076 25172 27132
rect 4274 27020 4284 27076
rect 4340 27020 9548 27076
rect 9604 27020 9614 27076
rect 11778 27020 11788 27076
rect 11844 27020 19404 27076
rect 19460 27020 19470 27076
rect 20514 27020 20524 27076
rect 20580 27020 22428 27076
rect 22484 27020 23100 27076
rect 23156 27020 23166 27076
rect 23986 27020 23996 27076
rect 24052 27020 25172 27076
rect 25330 27020 25340 27076
rect 25396 27020 26908 27076
rect 26964 27020 26974 27076
rect 28578 27020 28588 27076
rect 28644 27020 29148 27076
rect 29204 27020 29214 27076
rect 29810 27020 29820 27076
rect 29876 27020 30380 27076
rect 30436 27020 30446 27076
rect 31154 27020 31164 27076
rect 31220 27020 31836 27076
rect 31892 27020 31902 27076
rect 34066 27020 34076 27076
rect 34132 27020 34524 27076
rect 34580 27020 34590 27076
rect 36082 27020 36092 27076
rect 36148 27020 37324 27076
rect 37380 27020 37390 27076
rect 38210 27020 38220 27076
rect 38276 27020 39228 27076
rect 39284 27020 39676 27076
rect 39732 27020 39742 27076
rect 41346 27020 41356 27076
rect 41412 27020 42588 27076
rect 42644 27020 42654 27076
rect 0 26908 1988 26964
rect 2370 26908 2380 26964
rect 2436 26908 3164 26964
rect 3220 26908 4620 26964
rect 4676 26908 4686 26964
rect 9986 26908 9996 26964
rect 10052 26908 11116 26964
rect 11172 26908 11182 26964
rect 16258 26908 16268 26964
rect 16324 26908 17052 26964
rect 17108 26908 18620 26964
rect 18676 26908 18686 26964
rect 23538 26908 23548 26964
rect 23604 26908 24276 26964
rect 24770 26908 24780 26964
rect 24836 26908 25452 26964
rect 25508 26908 26348 26964
rect 26404 26908 26414 26964
rect 26562 26908 26572 26964
rect 26628 26908 31724 26964
rect 31780 26908 31790 26964
rect 38098 26908 38108 26964
rect 38164 26908 39004 26964
rect 39060 26908 39070 26964
rect 40114 26908 40124 26964
rect 40180 26908 44156 26964
rect 44212 26908 44716 26964
rect 44772 26908 45052 26964
rect 45108 26908 45118 26964
rect 0 26880 800 26908
rect 24210 26852 24220 26908
rect 24276 26852 24286 26908
rect 16930 26796 16940 26852
rect 16996 26796 21980 26852
rect 22036 26796 22046 26852
rect 26786 26796 26796 26852
rect 26852 26796 35084 26852
rect 35140 26796 35150 26852
rect 19282 26684 19292 26740
rect 19348 26684 19358 26740
rect 28354 26684 28364 26740
rect 28420 26684 33068 26740
rect 33124 26684 33134 26740
rect 19292 26516 19348 26684
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 24434 26572 24444 26628
rect 24500 26572 25116 26628
rect 25172 26572 25182 26628
rect 29922 26572 29932 26628
rect 29988 26572 31724 26628
rect 31780 26572 31790 26628
rect 35746 26572 35756 26628
rect 35812 26572 40124 26628
rect 40180 26572 40190 26628
rect 17938 26460 17948 26516
rect 18004 26460 20972 26516
rect 21028 26460 21038 26516
rect 24770 26460 24780 26516
rect 24836 26460 25788 26516
rect 25844 26460 25854 26516
rect 28018 26460 28028 26516
rect 28084 26460 28476 26516
rect 28532 26460 28542 26516
rect 34514 26460 34524 26516
rect 34580 26460 37100 26516
rect 37156 26460 37166 26516
rect 38770 26460 38780 26516
rect 38836 26460 39676 26516
rect 39732 26460 41580 26516
rect 41636 26460 41646 26516
rect 10210 26348 10220 26404
rect 10276 26348 11004 26404
rect 11060 26348 11676 26404
rect 11732 26348 11742 26404
rect 21970 26348 21980 26404
rect 22036 26348 23996 26404
rect 24052 26348 24062 26404
rect 28690 26348 28700 26404
rect 28756 26348 33292 26404
rect 33348 26348 33358 26404
rect 0 26292 800 26320
rect 0 26236 1932 26292
rect 1988 26236 1998 26292
rect 7746 26236 7756 26292
rect 7812 26236 8204 26292
rect 8260 26236 8270 26292
rect 8642 26236 8652 26292
rect 8708 26236 9996 26292
rect 10052 26236 10062 26292
rect 21746 26236 21756 26292
rect 21812 26236 23100 26292
rect 23156 26236 23548 26292
rect 23604 26236 23614 26292
rect 27458 26236 27468 26292
rect 27524 26236 28252 26292
rect 28308 26236 28318 26292
rect 30930 26236 30940 26292
rect 30996 26236 34300 26292
rect 34356 26236 34366 26292
rect 0 26208 800 26236
rect 8530 26124 8540 26180
rect 8596 26124 10052 26180
rect 18610 26124 18620 26180
rect 18676 26124 26124 26180
rect 26180 26124 26190 26180
rect 28354 26124 28364 26180
rect 28420 26124 34412 26180
rect 34468 26124 34478 26180
rect 9996 26068 10052 26124
rect 5058 26012 5068 26068
rect 5124 26012 6972 26068
rect 7028 26012 9212 26068
rect 9268 26012 9278 26068
rect 9986 26012 9996 26068
rect 10052 26012 18508 26068
rect 18564 26012 18574 26068
rect 20962 26012 20972 26068
rect 21028 26012 21308 26068
rect 21364 26012 22428 26068
rect 22484 26012 22494 26068
rect 24098 26012 24108 26068
rect 24164 26012 26236 26068
rect 26292 26012 26302 26068
rect 32386 26012 32396 26068
rect 32452 26012 32844 26068
rect 32900 26012 32910 26068
rect 17602 25900 17612 25956
rect 17668 25900 21644 25956
rect 21700 25900 22540 25956
rect 22596 25900 22606 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 4834 25788 4844 25844
rect 4900 25788 6188 25844
rect 6244 25788 8092 25844
rect 8148 25788 8158 25844
rect 2706 25676 2716 25732
rect 2772 25676 4620 25732
rect 4676 25676 4686 25732
rect 33842 25676 33852 25732
rect 33908 25676 35196 25732
rect 35252 25676 35262 25732
rect 0 25620 800 25648
rect 0 25564 2828 25620
rect 2884 25564 2894 25620
rect 4274 25564 4284 25620
rect 4340 25564 12460 25620
rect 12516 25564 12526 25620
rect 24994 25564 25004 25620
rect 25060 25564 26348 25620
rect 26404 25564 26414 25620
rect 27906 25564 27916 25620
rect 27972 25564 28364 25620
rect 28420 25564 28430 25620
rect 36428 25564 37772 25620
rect 37828 25564 37838 25620
rect 40114 25564 40124 25620
rect 40180 25564 40908 25620
rect 40964 25564 40974 25620
rect 0 25536 800 25564
rect 36428 25508 36484 25564
rect 6626 25452 6636 25508
rect 6692 25452 7756 25508
rect 7812 25452 7822 25508
rect 13468 25452 19852 25508
rect 19908 25452 19918 25508
rect 21634 25452 21644 25508
rect 21700 25452 22316 25508
rect 22372 25452 22382 25508
rect 23762 25452 23772 25508
rect 23828 25452 25564 25508
rect 25620 25452 25630 25508
rect 33740 25452 36428 25508
rect 36484 25452 36494 25508
rect 36754 25452 36764 25508
rect 36820 25452 41972 25508
rect 4722 25340 4732 25396
rect 4788 25340 10892 25396
rect 10948 25340 10958 25396
rect 3612 25228 5852 25284
rect 5908 25228 5918 25284
rect 10770 25228 10780 25284
rect 10836 25228 12796 25284
rect 12852 25228 12862 25284
rect 0 24948 800 24976
rect 3612 24948 3668 25228
rect 13468 25172 13524 25452
rect 33740 25396 33796 25452
rect 17714 25340 17724 25396
rect 17780 25340 21308 25396
rect 21364 25340 22652 25396
rect 22708 25340 22718 25396
rect 23426 25340 23436 25396
rect 23492 25340 27020 25396
rect 27076 25340 27086 25396
rect 28364 25340 33740 25396
rect 33796 25340 33806 25396
rect 34290 25340 34300 25396
rect 34356 25340 35644 25396
rect 35700 25340 35710 25396
rect 38612 25340 40684 25396
rect 40740 25340 40750 25396
rect 40898 25340 40908 25396
rect 40964 25340 41692 25396
rect 41748 25340 41758 25396
rect 28364 25284 28420 25340
rect 38612 25284 38668 25340
rect 41916 25284 41972 25452
rect 19628 25228 20244 25284
rect 25666 25228 25676 25284
rect 25732 25228 26236 25284
rect 26292 25228 26908 25284
rect 26964 25228 26974 25284
rect 27570 25228 27580 25284
rect 27636 25228 28364 25284
rect 28420 25228 28430 25284
rect 28578 25228 28588 25284
rect 28644 25228 32284 25284
rect 32340 25228 32350 25284
rect 33628 25228 38668 25284
rect 40226 25228 40236 25284
rect 40292 25228 41468 25284
rect 41524 25228 41534 25284
rect 41906 25228 41916 25284
rect 41972 25228 42140 25284
rect 42196 25228 42206 25284
rect 10546 25116 10556 25172
rect 10612 25116 13524 25172
rect 14018 25116 14028 25172
rect 14084 25116 15372 25172
rect 15428 25116 15438 25172
rect 18834 25116 18844 25172
rect 18900 25116 19404 25172
rect 19460 25116 19470 25172
rect 19628 25060 19684 25228
rect 20188 25172 20244 25228
rect 33628 25172 33684 25228
rect 20188 25116 23660 25172
rect 23716 25116 23996 25172
rect 24052 25116 27132 25172
rect 27188 25116 27198 25172
rect 27458 25116 27468 25172
rect 27524 25116 33684 25172
rect 37426 25116 37436 25172
rect 37492 25116 37660 25172
rect 37716 25116 37726 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 15092 25004 19684 25060
rect 20178 25004 20188 25060
rect 20244 25004 22764 25060
rect 22820 25004 22830 25060
rect 15092 24948 15148 25004
rect 0 24892 3668 24948
rect 14466 24892 14476 24948
rect 14532 24892 15148 24948
rect 19730 24892 19740 24948
rect 19796 24892 20412 24948
rect 20468 24892 20478 24948
rect 0 24864 800 24892
rect 4274 24780 4284 24836
rect 4340 24780 6972 24836
rect 7028 24780 7038 24836
rect 8418 24780 8428 24836
rect 8484 24780 11340 24836
rect 11396 24780 12348 24836
rect 12404 24780 12414 24836
rect 13468 24780 20188 24836
rect 20244 24780 20254 24836
rect 44482 24780 44492 24836
rect 44548 24780 45052 24836
rect 45108 24780 45118 24836
rect 9986 24668 9996 24724
rect 10052 24668 13244 24724
rect 13300 24668 13310 24724
rect 13468 24612 13524 24780
rect 15138 24668 15148 24724
rect 15204 24668 18620 24724
rect 18676 24668 23324 24724
rect 23380 24668 23390 24724
rect 24210 24668 24220 24724
rect 24276 24668 26124 24724
rect 26180 24668 26190 24724
rect 29586 24668 29596 24724
rect 29652 24668 30044 24724
rect 30100 24668 30110 24724
rect 38322 24668 38332 24724
rect 38388 24668 40012 24724
rect 40068 24668 44940 24724
rect 44996 24668 45006 24724
rect 1810 24556 1820 24612
rect 1876 24556 5852 24612
rect 5908 24556 7980 24612
rect 8036 24556 8046 24612
rect 8866 24556 8876 24612
rect 8932 24556 11900 24612
rect 11956 24556 13524 24612
rect 15092 24556 22316 24612
rect 22372 24556 22382 24612
rect 26786 24556 26796 24612
rect 26852 24556 39116 24612
rect 39172 24556 39182 24612
rect 44034 24556 44044 24612
rect 44100 24556 44828 24612
rect 44884 24556 44894 24612
rect 15092 24388 15148 24556
rect 37426 24444 37436 24500
rect 37492 24444 38108 24500
rect 38164 24444 38174 24500
rect 38434 24444 38444 24500
rect 38500 24444 45948 24500
rect 46004 24444 46014 24500
rect 38108 24388 38164 24444
rect 10770 24332 10780 24388
rect 10836 24332 15148 24388
rect 17154 24332 17164 24388
rect 17220 24332 31500 24388
rect 31556 24332 31566 24388
rect 38108 24332 39788 24388
rect 39844 24332 39854 24388
rect 0 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 0 24220 2044 24276
rect 2100 24220 2110 24276
rect 21298 24220 21308 24276
rect 21364 24220 26460 24276
rect 26516 24220 26526 24276
rect 38770 24220 38780 24276
rect 38836 24220 39116 24276
rect 39172 24220 39182 24276
rect 41906 24220 41916 24276
rect 41972 24220 41982 24276
rect 0 24192 800 24220
rect 12002 24108 12012 24164
rect 12068 24108 15148 24164
rect 16706 24108 16716 24164
rect 16772 24108 18620 24164
rect 18676 24108 27356 24164
rect 27412 24108 27422 24164
rect 31826 24108 31836 24164
rect 31892 24108 37660 24164
rect 37716 24108 37726 24164
rect 38434 24108 38444 24164
rect 38500 24108 40908 24164
rect 40964 24108 40974 24164
rect 15092 24052 15148 24108
rect 41916 24052 41972 24220
rect 15092 23996 19292 24052
rect 19348 23996 19358 24052
rect 24434 23996 24444 24052
rect 24500 23996 26684 24052
rect 26740 23996 26750 24052
rect 27794 23996 27804 24052
rect 27860 23996 41972 24052
rect 13010 23884 13020 23940
rect 13076 23884 14252 23940
rect 14308 23884 14700 23940
rect 14756 23884 14766 23940
rect 15362 23884 15372 23940
rect 15428 23884 15708 23940
rect 15764 23884 15774 23940
rect 19394 23884 19404 23940
rect 19460 23884 20188 23940
rect 20244 23884 20254 23940
rect 23314 23884 23324 23940
rect 23380 23884 24220 23940
rect 24276 23884 24286 23940
rect 26450 23884 26460 23940
rect 26516 23884 26908 23940
rect 29026 23884 29036 23940
rect 29092 23884 29932 23940
rect 29988 23884 29998 23940
rect 30370 23884 30380 23940
rect 30436 23884 31052 23940
rect 31108 23884 32620 23940
rect 32676 23884 32686 23940
rect 37762 23884 37772 23940
rect 37828 23884 39116 23940
rect 39172 23884 39620 23940
rect 40226 23884 40236 23940
rect 40292 23884 41132 23940
rect 41188 23884 41198 23940
rect 42466 23884 42476 23940
rect 42532 23884 43036 23940
rect 43092 23884 44940 23940
rect 44996 23884 45006 23940
rect 26852 23828 26908 23884
rect 6178 23772 6188 23828
rect 6244 23772 8652 23828
rect 8708 23772 8718 23828
rect 8978 23772 8988 23828
rect 9044 23772 9660 23828
rect 9716 23772 23548 23828
rect 23604 23772 23614 23828
rect 25218 23772 25228 23828
rect 25284 23772 26348 23828
rect 26404 23772 26414 23828
rect 26852 23772 32732 23828
rect 32788 23772 32798 23828
rect 35410 23772 35420 23828
rect 35476 23772 36988 23828
rect 37044 23772 37884 23828
rect 37940 23772 39004 23828
rect 39060 23772 39070 23828
rect 39564 23716 39620 23884
rect 39778 23772 39788 23828
rect 39844 23772 40796 23828
rect 40852 23772 44492 23828
rect 44548 23772 44558 23828
rect 6626 23660 6636 23716
rect 6692 23660 6702 23716
rect 15698 23660 15708 23716
rect 15764 23660 18172 23716
rect 18228 23660 19292 23716
rect 19348 23660 19740 23716
rect 19796 23660 19806 23716
rect 22754 23660 22764 23716
rect 22820 23660 23436 23716
rect 23492 23660 23502 23716
rect 25666 23660 25676 23716
rect 25732 23660 27692 23716
rect 27748 23660 27758 23716
rect 29362 23660 29372 23716
rect 29428 23660 31388 23716
rect 31444 23660 31454 23716
rect 36194 23660 36204 23716
rect 36260 23660 37212 23716
rect 37268 23660 38556 23716
rect 38612 23660 38622 23716
rect 39564 23660 44772 23716
rect 0 23604 800 23632
rect 6636 23604 6692 23660
rect 44716 23604 44772 23660
rect 0 23548 6692 23604
rect 8372 23548 8820 23604
rect 11890 23548 11900 23604
rect 11956 23548 12796 23604
rect 12852 23548 14644 23604
rect 44706 23548 44716 23604
rect 44772 23548 44782 23604
rect 0 23520 800 23548
rect 8372 23492 8428 23548
rect 6962 23436 6972 23492
rect 7028 23436 8428 23492
rect 8764 23492 8820 23548
rect 8764 23436 10444 23492
rect 10500 23436 10510 23492
rect 12562 23436 12572 23492
rect 12628 23436 12908 23492
rect 12964 23436 14364 23492
rect 14420 23436 14430 23492
rect 14588 23380 14644 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 14914 23436 14924 23492
rect 14980 23436 15372 23492
rect 15428 23436 15438 23492
rect 15670 23436 15708 23492
rect 15764 23436 15774 23492
rect 20514 23436 20524 23492
rect 20580 23436 22988 23492
rect 23044 23436 23054 23492
rect 30594 23436 30604 23492
rect 30660 23436 33180 23492
rect 33236 23436 33246 23492
rect 4946 23324 4956 23380
rect 5012 23324 5852 23380
rect 5908 23324 5918 23380
rect 6402 23324 6412 23380
rect 6468 23324 7644 23380
rect 7700 23324 7710 23380
rect 14588 23324 20748 23380
rect 20804 23324 20814 23380
rect 24546 23324 24556 23380
rect 24612 23324 26908 23380
rect 27234 23324 27244 23380
rect 27300 23324 27916 23380
rect 27972 23324 29372 23380
rect 29428 23324 29438 23380
rect 31490 23324 31500 23380
rect 31556 23324 32284 23380
rect 32340 23324 32350 23380
rect 26852 23268 26908 23324
rect 6850 23212 6860 23268
rect 6916 23212 9436 23268
rect 9492 23212 9502 23268
rect 9874 23212 9884 23268
rect 9940 23212 10668 23268
rect 10724 23212 10734 23268
rect 14466 23212 14476 23268
rect 14532 23212 15036 23268
rect 15092 23212 16660 23268
rect 18498 23212 18508 23268
rect 18564 23212 20300 23268
rect 20356 23212 21756 23268
rect 21812 23212 21822 23268
rect 25750 23212 25788 23268
rect 25844 23212 25854 23268
rect 26852 23212 37100 23268
rect 37156 23212 37166 23268
rect 10434 23100 10444 23156
rect 10500 23100 10780 23156
rect 10836 23100 10846 23156
rect 13906 23100 13916 23156
rect 13972 23100 15596 23156
rect 15652 23100 15662 23156
rect 16604 23044 16660 23212
rect 17938 23100 17948 23156
rect 18004 23100 21420 23156
rect 21476 23100 21486 23156
rect 22166 23100 22204 23156
rect 22260 23100 22270 23156
rect 32610 23100 32620 23156
rect 32676 23100 33180 23156
rect 33236 23100 33852 23156
rect 33908 23100 33918 23156
rect 34066 23100 34076 23156
rect 34132 23100 36204 23156
rect 36260 23100 36270 23156
rect 43026 23100 43036 23156
rect 43092 23100 45500 23156
rect 45556 23100 45566 23156
rect 34076 23044 34132 23100
rect 2370 22988 2380 23044
rect 2436 22988 8540 23044
rect 8596 22988 8606 23044
rect 16594 22988 16604 23044
rect 16660 22988 25452 23044
rect 25508 22988 25518 23044
rect 25788 22988 26124 23044
rect 26180 22988 26684 23044
rect 26740 22988 26750 23044
rect 33618 22988 33628 23044
rect 33684 22988 34132 23044
rect 0 22932 800 22960
rect 25788 22932 25844 22988
rect 0 22876 2716 22932
rect 2772 22876 2782 22932
rect 22866 22876 22876 22932
rect 22932 22876 23436 22932
rect 23492 22876 23502 22932
rect 25330 22876 25340 22932
rect 25396 22876 25844 22932
rect 26002 22876 26012 22932
rect 26068 22876 26796 22932
rect 26852 22876 26862 22932
rect 33506 22876 33516 22932
rect 33572 22876 35868 22932
rect 35924 22876 35934 22932
rect 0 22848 800 22876
rect 15670 22764 15708 22820
rect 15764 22764 15774 22820
rect 23174 22764 23212 22820
rect 23268 22764 23278 22820
rect 24668 22764 27244 22820
rect 27300 22764 27310 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 24668 22708 24724 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 21410 22652 21420 22708
rect 21476 22652 23548 22708
rect 23604 22652 23772 22708
rect 23828 22652 23838 22708
rect 24658 22652 24668 22708
rect 24724 22652 24734 22708
rect 11666 22540 11676 22596
rect 11732 22540 12236 22596
rect 12292 22540 28364 22596
rect 28420 22540 28430 22596
rect 15698 22428 15708 22484
rect 15764 22428 16492 22484
rect 16548 22428 16558 22484
rect 20514 22428 20524 22484
rect 20580 22428 23324 22484
rect 23380 22428 23390 22484
rect 30146 22428 30156 22484
rect 30212 22428 30604 22484
rect 30660 22428 30670 22484
rect 35186 22428 35196 22484
rect 35252 22428 38668 22484
rect 38724 22428 38892 22484
rect 38948 22428 38958 22484
rect 4722 22316 4732 22372
rect 4788 22316 5964 22372
rect 6020 22316 6030 22372
rect 6402 22316 6412 22372
rect 6468 22316 8428 22372
rect 8484 22316 8494 22372
rect 17826 22316 17836 22372
rect 17892 22316 19964 22372
rect 20020 22316 20030 22372
rect 20626 22316 20636 22372
rect 20692 22316 21420 22372
rect 21476 22316 21486 22372
rect 21858 22316 21868 22372
rect 21924 22316 26908 22372
rect 26964 22316 26974 22372
rect 27570 22316 27580 22372
rect 27636 22316 29036 22372
rect 29092 22316 29102 22372
rect 29250 22316 29260 22372
rect 29316 22316 29820 22372
rect 29876 22316 29886 22372
rect 33506 22316 33516 22372
rect 33572 22316 35532 22372
rect 35588 22316 35598 22372
rect 42578 22316 42588 22372
rect 42644 22316 43484 22372
rect 43540 22316 43550 22372
rect 7074 22204 7084 22260
rect 7140 22204 12796 22260
rect 12852 22204 18396 22260
rect 18452 22204 18462 22260
rect 24322 22204 24332 22260
rect 24388 22204 26908 22260
rect 27906 22204 27916 22260
rect 27972 22204 29148 22260
rect 29204 22204 29214 22260
rect 32274 22204 32284 22260
rect 32340 22204 34972 22260
rect 35028 22204 35038 22260
rect 35858 22204 35868 22260
rect 35924 22204 37884 22260
rect 37940 22204 37950 22260
rect 26852 22148 26908 22204
rect 4274 22092 4284 22148
rect 4340 22092 8204 22148
rect 8260 22092 8270 22148
rect 12450 22092 12460 22148
rect 12516 22092 13580 22148
rect 13636 22092 13646 22148
rect 19282 22092 19292 22148
rect 19348 22092 22932 22148
rect 23090 22092 23100 22148
rect 23156 22092 25788 22148
rect 25844 22092 25854 22148
rect 26852 22092 32340 22148
rect 22876 22036 22932 22092
rect 32284 22036 32340 22092
rect 15362 21980 15372 22036
rect 15428 21980 15708 22036
rect 15764 21980 15774 22036
rect 16034 21980 16044 22036
rect 16100 21980 18172 22036
rect 18228 21980 18238 22036
rect 22876 21980 24444 22036
rect 24500 21980 25004 22036
rect 25060 21980 25070 22036
rect 26114 21980 26124 22036
rect 26180 21980 26684 22036
rect 26740 21980 26750 22036
rect 29026 21980 29036 22036
rect 29092 21980 30716 22036
rect 30772 21980 30782 22036
rect 32274 21980 32284 22036
rect 32340 21980 32350 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 13010 21868 13020 21924
rect 13076 21868 13804 21924
rect 13860 21868 14700 21924
rect 14756 21868 14766 21924
rect 15026 21868 15036 21924
rect 15092 21868 17164 21924
rect 17220 21868 17230 21924
rect 28578 21868 28588 21924
rect 28644 21868 29596 21924
rect 29652 21868 31164 21924
rect 31220 21868 33292 21924
rect 33348 21868 33358 21924
rect 8082 21756 8092 21812
rect 8148 21756 10220 21812
rect 10276 21756 10286 21812
rect 10668 21756 11676 21812
rect 11732 21756 11742 21812
rect 14914 21756 14924 21812
rect 14980 21756 17836 21812
rect 17892 21756 17902 21812
rect 19506 21756 19516 21812
rect 19572 21756 20412 21812
rect 20468 21756 20478 21812
rect 20626 21756 20636 21812
rect 20692 21756 21532 21812
rect 21588 21756 22092 21812
rect 22148 21756 22158 21812
rect 22306 21756 22316 21812
rect 22372 21756 27132 21812
rect 27188 21756 27198 21812
rect 37986 21756 37996 21812
rect 38052 21756 38444 21812
rect 38500 21756 40012 21812
rect 40068 21756 40078 21812
rect 10668 21700 10724 21756
rect 7410 21644 7420 21700
rect 7476 21644 10724 21700
rect 10780 21644 13132 21700
rect 13188 21644 14028 21700
rect 14084 21644 14094 21700
rect 16482 21644 16492 21700
rect 16548 21644 16828 21700
rect 16884 21644 16894 21700
rect 20962 21644 20972 21700
rect 21028 21644 25788 21700
rect 25844 21644 25854 21700
rect 28018 21644 28028 21700
rect 28084 21644 30268 21700
rect 30324 21644 30334 21700
rect 30594 21644 30604 21700
rect 30660 21644 31276 21700
rect 31332 21644 33740 21700
rect 33796 21644 33806 21700
rect 34514 21644 34524 21700
rect 34580 21644 35980 21700
rect 36036 21644 36046 21700
rect 38098 21644 38108 21700
rect 38164 21644 41132 21700
rect 41188 21644 41198 21700
rect 41458 21644 41468 21700
rect 41524 21644 42700 21700
rect 42756 21644 43596 21700
rect 43652 21644 43662 21700
rect 0 21588 800 21616
rect 10780 21588 10836 21644
rect 0 21532 1708 21588
rect 1764 21532 1774 21588
rect 7522 21532 7532 21588
rect 7588 21532 10836 21588
rect 10994 21532 11004 21588
rect 11060 21532 11788 21588
rect 11844 21532 11854 21588
rect 16146 21532 16156 21588
rect 16212 21532 17500 21588
rect 17556 21532 17566 21588
rect 18386 21532 18396 21588
rect 18452 21532 22652 21588
rect 22708 21532 22718 21588
rect 27234 21532 27244 21588
rect 27300 21532 27804 21588
rect 27860 21532 27870 21588
rect 28550 21532 28588 21588
rect 28644 21532 28654 21588
rect 31490 21532 31500 21588
rect 31556 21532 32956 21588
rect 33012 21532 33022 21588
rect 33954 21532 33964 21588
rect 34020 21532 35084 21588
rect 35140 21532 35150 21588
rect 0 21504 800 21532
rect 14354 21420 14364 21476
rect 14420 21420 18284 21476
rect 18340 21420 18350 21476
rect 22082 21420 22092 21476
rect 22148 21420 24892 21476
rect 24948 21420 24958 21476
rect 27010 21420 27020 21476
rect 27076 21420 28364 21476
rect 28420 21420 28430 21476
rect 10210 21308 10220 21364
rect 10276 21308 17388 21364
rect 17444 21308 18060 21364
rect 18116 21308 18126 21364
rect 22530 21308 22540 21364
rect 22596 21308 23324 21364
rect 23380 21308 23390 21364
rect 28690 21308 28700 21364
rect 28756 21308 31164 21364
rect 31220 21308 31230 21364
rect 31388 21308 36204 21364
rect 36260 21308 36270 21364
rect 31388 21252 31444 21308
rect 20850 21196 20860 21252
rect 20916 21196 26572 21252
rect 26628 21196 26638 21252
rect 28354 21196 28364 21252
rect 28420 21196 31444 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 20290 21084 20300 21140
rect 20356 21084 27244 21140
rect 27300 21084 27310 21140
rect 13570 20972 13580 21028
rect 13636 20972 14924 21028
rect 14980 20972 14990 21028
rect 32050 20972 32060 21028
rect 32116 20972 33740 21028
rect 33796 20972 33806 21028
rect 0 20916 800 20944
rect 0 20860 1820 20916
rect 1876 20860 1886 20916
rect 10546 20860 10556 20916
rect 10612 20860 11340 20916
rect 11396 20860 11406 20916
rect 13458 20860 13468 20916
rect 13524 20860 16828 20916
rect 16884 20860 16894 20916
rect 19618 20860 19628 20916
rect 19684 20860 20300 20916
rect 20356 20860 20366 20916
rect 22866 20860 22876 20916
rect 22932 20860 28644 20916
rect 29698 20860 29708 20916
rect 29764 20860 30492 20916
rect 30548 20860 30558 20916
rect 0 20832 800 20860
rect 28588 20804 28644 20860
rect 6290 20748 6300 20804
rect 6356 20748 7532 20804
rect 7588 20748 7598 20804
rect 14130 20748 14140 20804
rect 14196 20748 14812 20804
rect 14868 20748 17164 20804
rect 17220 20748 17230 20804
rect 26114 20748 26124 20804
rect 26180 20748 26796 20804
rect 26852 20748 26862 20804
rect 27122 20748 27132 20804
rect 27188 20748 27804 20804
rect 27860 20748 27870 20804
rect 28578 20748 28588 20804
rect 28644 20748 29260 20804
rect 29316 20748 29326 20804
rect 33282 20748 33292 20804
rect 33348 20748 34524 20804
rect 34580 20748 34590 20804
rect 14914 20636 14924 20692
rect 14980 20636 15148 20692
rect 16034 20636 16044 20692
rect 16100 20636 17276 20692
rect 17332 20636 17342 20692
rect 34402 20636 34412 20692
rect 34468 20636 35980 20692
rect 36036 20636 36046 20692
rect 42130 20636 42140 20692
rect 42196 20636 42476 20692
rect 42532 20636 42542 20692
rect 15092 20580 15148 20636
rect 5058 20524 5068 20580
rect 5124 20524 6636 20580
rect 6692 20524 6702 20580
rect 9874 20524 9884 20580
rect 9940 20524 11004 20580
rect 11060 20524 11070 20580
rect 15092 20524 15932 20580
rect 15988 20524 17388 20580
rect 17444 20524 17454 20580
rect 22082 20524 22092 20580
rect 22148 20524 22204 20580
rect 22260 20524 22270 20580
rect 4274 20412 4284 20468
rect 4340 20412 5964 20468
rect 6020 20412 6860 20468
rect 6916 20412 7644 20468
rect 7700 20412 7710 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 28690 20300 28700 20356
rect 28756 20300 29260 20356
rect 29316 20300 30380 20356
rect 30436 20300 30446 20356
rect 35746 20300 35756 20356
rect 35812 20300 37660 20356
rect 37716 20300 37726 20356
rect 0 20244 800 20272
rect 0 20188 1932 20244
rect 1988 20188 1998 20244
rect 3154 20188 3164 20244
rect 3220 20188 16772 20244
rect 27458 20188 27468 20244
rect 27524 20188 30212 20244
rect 33506 20188 33516 20244
rect 33572 20188 34860 20244
rect 34916 20188 34926 20244
rect 36754 20188 36764 20244
rect 36820 20188 42028 20244
rect 42084 20188 43316 20244
rect 0 20160 800 20188
rect 1698 20076 1708 20132
rect 1764 20076 3388 20132
rect 10434 20076 10444 20132
rect 10500 20076 11676 20132
rect 11732 20076 12572 20132
rect 12628 20076 12638 20132
rect 15092 20076 15260 20132
rect 15316 20076 15326 20132
rect 3332 20020 3388 20076
rect 15092 20020 15148 20076
rect 16716 20020 16772 20188
rect 30156 20132 30212 20188
rect 43260 20132 43316 20188
rect 17378 20076 17388 20132
rect 17444 20076 17454 20132
rect 20066 20076 20076 20132
rect 20132 20076 21084 20132
rect 21140 20076 23772 20132
rect 23828 20076 23838 20132
rect 30156 20076 36092 20132
rect 36148 20076 36158 20132
rect 38210 20076 38220 20132
rect 38276 20076 42812 20132
rect 42868 20076 42878 20132
rect 43250 20076 43260 20132
rect 43316 20076 43326 20132
rect 3332 19964 6412 20020
rect 6468 19964 6478 20020
rect 8866 19964 8876 20020
rect 8932 19964 10556 20020
rect 10612 19964 10622 20020
rect 11442 19964 11452 20020
rect 11508 19964 12348 20020
rect 12404 19964 12796 20020
rect 12852 19964 12862 20020
rect 13682 19964 13692 20020
rect 13748 19964 15148 20020
rect 16706 19964 16716 20020
rect 16772 19964 16782 20020
rect 17388 19908 17444 20076
rect 25442 19964 25452 20020
rect 25508 19964 31724 20020
rect 31780 19964 33180 20020
rect 33236 19964 33246 20020
rect 39218 19964 39228 20020
rect 39284 19964 39788 20020
rect 39844 19964 39854 20020
rect 40226 19964 40236 20020
rect 40292 19964 41356 20020
rect 41412 19964 41422 20020
rect 4162 19852 4172 19908
rect 4228 19852 5628 19908
rect 5684 19852 5694 19908
rect 8372 19852 12012 19908
rect 12068 19852 12078 19908
rect 12226 19852 12236 19908
rect 12292 19852 13580 19908
rect 13636 19852 13646 19908
rect 13794 19852 13804 19908
rect 13860 19852 17444 19908
rect 22530 19852 22540 19908
rect 22596 19852 24556 19908
rect 24612 19852 26124 19908
rect 26180 19852 26190 19908
rect 39890 19852 39900 19908
rect 39956 19852 40572 19908
rect 40628 19852 40638 19908
rect 8372 19796 8428 19852
rect 12236 19796 12292 19852
rect 2034 19740 2044 19796
rect 2100 19740 8428 19796
rect 8754 19740 8764 19796
rect 8820 19740 11116 19796
rect 11172 19740 11182 19796
rect 11330 19740 11340 19796
rect 11396 19740 12292 19796
rect 14242 19740 14252 19796
rect 14308 19740 15708 19796
rect 15764 19740 15774 19796
rect 16706 19740 16716 19796
rect 16772 19740 18172 19796
rect 18228 19740 18238 19796
rect 32498 19740 32508 19796
rect 32564 19740 37436 19796
rect 37492 19740 38668 19796
rect 38724 19740 39564 19796
rect 39620 19740 39630 19796
rect 13570 19628 13580 19684
rect 13636 19628 18620 19684
rect 18676 19628 18686 19684
rect 32162 19628 32172 19684
rect 32228 19628 34076 19684
rect 34132 19628 34142 19684
rect 37538 19628 37548 19684
rect 37604 19628 37884 19684
rect 37940 19628 40348 19684
rect 40404 19628 40908 19684
rect 40964 19628 40974 19684
rect 0 19572 800 19600
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 0 19516 3500 19572
rect 3556 19516 3566 19572
rect 10098 19516 10108 19572
rect 10164 19516 10780 19572
rect 10836 19516 10846 19572
rect 11778 19516 11788 19572
rect 11844 19516 19628 19572
rect 19684 19516 19694 19572
rect 0 19488 800 19516
rect 2930 19404 2940 19460
rect 2996 19404 4508 19460
rect 4564 19404 4574 19460
rect 4834 19404 4844 19460
rect 4900 19404 7196 19460
rect 7252 19404 7262 19460
rect 10658 19404 10668 19460
rect 10724 19404 12796 19460
rect 12852 19404 12862 19460
rect 13458 19404 13468 19460
rect 13524 19404 14476 19460
rect 14532 19404 17612 19460
rect 17668 19404 17678 19460
rect 26852 19404 40460 19460
rect 40516 19404 40526 19460
rect 26852 19348 26908 19404
rect 4610 19292 4620 19348
rect 4676 19292 6076 19348
rect 6132 19292 6142 19348
rect 6738 19292 6748 19348
rect 6804 19292 13692 19348
rect 13748 19292 13758 19348
rect 15698 19292 15708 19348
rect 15764 19292 18508 19348
rect 18564 19292 18574 19348
rect 21746 19292 21756 19348
rect 21812 19292 22764 19348
rect 22820 19292 22830 19348
rect 24770 19292 24780 19348
rect 24836 19292 26908 19348
rect 33506 19292 33516 19348
rect 33572 19292 42140 19348
rect 42196 19292 42206 19348
rect 2258 19180 2268 19236
rect 2324 19180 8428 19236
rect 12674 19180 12684 19236
rect 12740 19180 13804 19236
rect 13860 19180 13870 19236
rect 36082 19180 36092 19236
rect 36148 19180 38220 19236
rect 38276 19180 38286 19236
rect 38882 19180 38892 19236
rect 38948 19180 40236 19236
rect 40292 19180 40302 19236
rect 8372 19124 8428 19180
rect 1922 19068 1932 19124
rect 1988 19068 2604 19124
rect 2660 19068 6636 19124
rect 6692 19068 6702 19124
rect 8372 19068 13356 19124
rect 13412 19068 14028 19124
rect 14084 19068 14094 19124
rect 16706 19068 16716 19124
rect 16772 19068 17948 19124
rect 18004 19068 18014 19124
rect 32386 19068 32396 19124
rect 32452 19068 34412 19124
rect 34468 19068 34478 19124
rect 34738 19068 34748 19124
rect 34804 19068 35420 19124
rect 35476 19068 35868 19124
rect 35924 19068 36988 19124
rect 37044 19068 37054 19124
rect 38434 19068 38444 19124
rect 38500 19068 39900 19124
rect 39956 19068 42588 19124
rect 42644 19068 42654 19124
rect 3826 18956 3836 19012
rect 3892 18956 13580 19012
rect 13636 18956 13646 19012
rect 13794 18956 13804 19012
rect 13860 18956 15372 19012
rect 15428 18956 16380 19012
rect 16436 18956 16828 19012
rect 16884 18956 16894 19012
rect 29362 18956 29372 19012
rect 29428 18956 35532 19012
rect 35588 18956 35756 19012
rect 35812 18956 35822 19012
rect 36530 18956 36540 19012
rect 36596 18956 37100 19012
rect 37156 18956 37166 19012
rect 0 18900 800 18928
rect 0 18844 1820 18900
rect 1876 18844 1886 18900
rect 12338 18844 12348 18900
rect 12404 18844 15932 18900
rect 15988 18844 18956 18900
rect 19012 18844 19022 18900
rect 0 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 2146 18732 2156 18788
rect 2212 18732 4956 18788
rect 5012 18732 5022 18788
rect 13010 18732 13020 18788
rect 13076 18732 15596 18788
rect 15652 18732 18060 18788
rect 18116 18732 18126 18788
rect 12786 18620 12796 18676
rect 12852 18620 14028 18676
rect 14084 18620 14094 18676
rect 15474 18620 15484 18676
rect 15540 18620 16380 18676
rect 16436 18620 16446 18676
rect 21186 18620 21196 18676
rect 21252 18620 23548 18676
rect 23604 18620 23614 18676
rect 35634 18620 35644 18676
rect 35700 18620 37884 18676
rect 37940 18620 38668 18676
rect 38612 18564 38668 18620
rect 1698 18508 1708 18564
rect 1764 18508 2156 18564
rect 2212 18508 2222 18564
rect 12898 18508 12908 18564
rect 12964 18508 12974 18564
rect 17826 18508 17836 18564
rect 17892 18508 18508 18564
rect 18564 18508 18574 18564
rect 19730 18508 19740 18564
rect 19796 18508 22540 18564
rect 22596 18508 22606 18564
rect 24098 18508 24108 18564
rect 24164 18508 31948 18564
rect 32004 18508 33068 18564
rect 33124 18508 33134 18564
rect 38546 18508 38556 18564
rect 38612 18508 41356 18564
rect 41412 18508 41422 18564
rect 12908 18452 12964 18508
rect 3378 18396 3388 18452
rect 3444 18396 4956 18452
rect 5012 18396 5022 18452
rect 8978 18396 8988 18452
rect 9044 18396 10332 18452
rect 10388 18396 10398 18452
rect 12908 18396 13244 18452
rect 13300 18396 13310 18452
rect 14690 18396 14700 18452
rect 14756 18396 18172 18452
rect 18228 18396 18238 18452
rect 23090 18396 23100 18452
rect 23156 18396 23884 18452
rect 23940 18396 24220 18452
rect 24276 18396 24286 18452
rect 32722 18396 32732 18452
rect 32788 18396 34748 18452
rect 34804 18396 34814 18452
rect 34962 18396 34972 18452
rect 35028 18396 35308 18452
rect 35364 18396 35374 18452
rect 36642 18396 36652 18452
rect 36708 18396 39004 18452
rect 39060 18396 39070 18452
rect 39442 18396 39452 18452
rect 39508 18396 40012 18452
rect 40068 18396 43596 18452
rect 43652 18396 43662 18452
rect 44930 18396 44940 18452
rect 44996 18396 45948 18452
rect 46004 18396 46014 18452
rect 2258 18284 2268 18340
rect 2324 18284 6748 18340
rect 6804 18284 6814 18340
rect 12898 18284 12908 18340
rect 12964 18284 15708 18340
rect 15764 18284 15774 18340
rect 17602 18284 17612 18340
rect 17668 18284 19292 18340
rect 19348 18284 20524 18340
rect 20580 18284 20590 18340
rect 25330 18284 25340 18340
rect 25396 18284 26236 18340
rect 26292 18284 26302 18340
rect 31714 18284 31724 18340
rect 31780 18284 33180 18340
rect 33236 18284 33246 18340
rect 34514 18284 34524 18340
rect 34580 18284 37436 18340
rect 37492 18284 37502 18340
rect 38322 18284 38332 18340
rect 38388 18284 38780 18340
rect 38836 18284 38846 18340
rect 0 18228 800 18256
rect 37436 18228 37492 18284
rect 0 18172 1708 18228
rect 1764 18172 1774 18228
rect 5170 18172 5180 18228
rect 5236 18172 6412 18228
rect 6468 18172 6478 18228
rect 7298 18172 7308 18228
rect 7364 18172 15484 18228
rect 15540 18172 16828 18228
rect 16884 18172 17948 18228
rect 18004 18172 35868 18228
rect 35924 18172 35934 18228
rect 37436 18172 38892 18228
rect 38948 18172 39116 18228
rect 39172 18172 39182 18228
rect 0 18144 800 18172
rect 15026 18060 15036 18116
rect 15092 18060 16268 18116
rect 16324 18060 17836 18116
rect 17892 18060 24668 18116
rect 24724 18060 24734 18116
rect 32498 18060 32508 18116
rect 32564 18060 33628 18116
rect 33684 18060 34972 18116
rect 35028 18060 35038 18116
rect 35532 18060 38332 18116
rect 38388 18060 38398 18116
rect 39218 18060 39228 18116
rect 39284 18060 39676 18116
rect 39732 18060 39742 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 9650 17948 9660 18004
rect 9716 17948 10444 18004
rect 10500 17948 11564 18004
rect 11620 17948 29372 18004
rect 29428 17948 29596 18004
rect 29652 17948 29662 18004
rect 35532 17892 35588 18060
rect 2370 17836 2380 17892
rect 2436 17836 4060 17892
rect 4116 17836 4126 17892
rect 8082 17836 8092 17892
rect 8148 17836 10668 17892
rect 10724 17836 10734 17892
rect 20374 17836 20412 17892
rect 20468 17836 20478 17892
rect 35074 17836 35084 17892
rect 35140 17836 35588 17892
rect 35756 17836 39676 17892
rect 39732 17836 39742 17892
rect 35756 17780 35812 17836
rect 1698 17724 1708 17780
rect 1764 17724 4620 17780
rect 4676 17724 4686 17780
rect 16594 17724 16604 17780
rect 16660 17724 22876 17780
rect 22932 17724 22942 17780
rect 30370 17724 30380 17780
rect 30436 17724 31388 17780
rect 31444 17724 35812 17780
rect 36418 17724 36428 17780
rect 36484 17724 37436 17780
rect 37492 17724 42252 17780
rect 42308 17724 42318 17780
rect 1708 17612 3500 17668
rect 3556 17612 6076 17668
rect 6132 17612 6142 17668
rect 11666 17612 11676 17668
rect 11732 17612 12124 17668
rect 12180 17612 12190 17668
rect 13682 17612 13692 17668
rect 13748 17612 15372 17668
rect 15428 17612 15438 17668
rect 18732 17612 23212 17668
rect 23268 17612 25004 17668
rect 25060 17612 25070 17668
rect 31714 17612 31724 17668
rect 31780 17612 33740 17668
rect 33796 17612 34972 17668
rect 35028 17612 35038 17668
rect 1708 17444 1764 17612
rect 18732 17556 18788 17612
rect 3602 17500 3612 17556
rect 3668 17500 9212 17556
rect 9268 17500 9278 17556
rect 12226 17500 12236 17556
rect 12292 17500 12908 17556
rect 12964 17500 13580 17556
rect 13636 17500 18396 17556
rect 18452 17500 18462 17556
rect 18722 17500 18732 17556
rect 18788 17500 18798 17556
rect 19394 17500 19404 17556
rect 19460 17500 20076 17556
rect 20132 17500 21980 17556
rect 22036 17500 23436 17556
rect 23492 17500 23502 17556
rect 28242 17500 28252 17556
rect 28308 17500 29708 17556
rect 29764 17500 29774 17556
rect 35298 17500 35308 17556
rect 35364 17500 35644 17556
rect 35700 17500 35710 17556
rect 36418 17500 36428 17556
rect 36484 17500 36988 17556
rect 37044 17500 37054 17556
rect 1698 17388 1708 17444
rect 1764 17388 1774 17444
rect 2034 17388 2044 17444
rect 2100 17388 2110 17444
rect 2706 17388 2716 17444
rect 2772 17388 11564 17444
rect 11620 17388 11956 17444
rect 15922 17388 15932 17444
rect 15988 17388 17388 17444
rect 17444 17388 17454 17444
rect 2044 17332 2100 17388
rect 2044 17276 11676 17332
rect 11732 17276 11742 17332
rect 4162 17164 4172 17220
rect 4228 17164 5628 17220
rect 5684 17164 5694 17220
rect 6178 17164 6188 17220
rect 6244 17164 8540 17220
rect 8596 17164 9548 17220
rect 9604 17164 9614 17220
rect 5628 17108 5684 17164
rect 5628 17052 8428 17108
rect 8484 17052 8494 17108
rect 0 16884 800 16912
rect 11900 16884 11956 17388
rect 20300 17276 21532 17332
rect 21588 17276 22540 17332
rect 22596 17276 22606 17332
rect 28578 17276 28588 17332
rect 28644 17276 30044 17332
rect 30100 17276 38220 17332
rect 38276 17276 38286 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 20300 17220 20356 17276
rect 20290 17164 20300 17220
rect 20356 17164 20366 17220
rect 39554 17164 39564 17220
rect 39620 17164 42028 17220
rect 42084 17164 44380 17220
rect 44436 17164 44446 17220
rect 13122 17052 13132 17108
rect 13188 17052 16268 17108
rect 16324 17052 16334 17108
rect 18050 17052 18060 17108
rect 18116 17052 18732 17108
rect 18788 17052 18798 17108
rect 24658 17052 24668 17108
rect 24724 17052 26796 17108
rect 26852 17052 26862 17108
rect 28354 17052 28364 17108
rect 28420 17052 28430 17108
rect 37762 17052 37772 17108
rect 37828 17052 38556 17108
rect 38612 17052 38622 17108
rect 28364 16996 28420 17052
rect 12114 16940 12124 16996
rect 12180 16940 12908 16996
rect 12964 16940 12974 16996
rect 28364 16940 30604 16996
rect 30660 16940 30828 16996
rect 30884 16940 36540 16996
rect 36596 16940 36606 16996
rect 38882 16940 38892 16996
rect 38948 16940 39900 16996
rect 39956 16940 43484 16996
rect 43540 16940 43550 16996
rect 0 16828 2380 16884
rect 2436 16828 2446 16884
rect 6066 16828 6076 16884
rect 6132 16828 9100 16884
rect 9156 16828 9166 16884
rect 10658 16828 10668 16884
rect 10724 16828 10734 16884
rect 11900 16828 12684 16884
rect 12740 16828 12750 16884
rect 13906 16828 13916 16884
rect 13972 16828 16380 16884
rect 16436 16828 16446 16884
rect 19506 16828 19516 16884
rect 19572 16828 22652 16884
rect 22708 16828 23884 16884
rect 23940 16828 23950 16884
rect 32274 16828 32284 16884
rect 32340 16828 39452 16884
rect 39508 16828 41244 16884
rect 41300 16828 41310 16884
rect 42354 16828 42364 16884
rect 42420 16828 43372 16884
rect 43428 16828 45052 16884
rect 45108 16828 45118 16884
rect 0 16800 800 16828
rect 10668 16772 10724 16828
rect 8194 16716 8204 16772
rect 8260 16716 8988 16772
rect 9044 16716 9054 16772
rect 9650 16716 9660 16772
rect 9716 16716 10724 16772
rect 11442 16716 11452 16772
rect 11508 16716 19180 16772
rect 19236 16716 19246 16772
rect 20402 16716 20412 16772
rect 20468 16716 20478 16772
rect 21634 16716 21644 16772
rect 21700 16716 23772 16772
rect 23828 16716 23838 16772
rect 27458 16716 27468 16772
rect 27524 16716 29596 16772
rect 29652 16716 29662 16772
rect 30930 16716 30940 16772
rect 30996 16716 33740 16772
rect 33796 16716 33806 16772
rect 34178 16716 34188 16772
rect 34244 16716 36316 16772
rect 36372 16716 36382 16772
rect 11452 16660 11508 16716
rect 20412 16660 20468 16716
rect 9986 16604 9996 16660
rect 10052 16604 11508 16660
rect 12562 16604 12572 16660
rect 12628 16604 15932 16660
rect 15988 16604 15998 16660
rect 16594 16604 16604 16660
rect 16660 16604 17724 16660
rect 17780 16604 20468 16660
rect 21858 16604 21868 16660
rect 21924 16604 21934 16660
rect 25666 16604 25676 16660
rect 25732 16604 26012 16660
rect 26068 16604 26078 16660
rect 32834 16604 32844 16660
rect 32900 16604 32910 16660
rect 33058 16604 33068 16660
rect 33124 16604 35532 16660
rect 35588 16604 35598 16660
rect 16604 16548 16660 16604
rect 21868 16548 21924 16604
rect 12226 16492 12236 16548
rect 12292 16492 16660 16548
rect 18722 16492 18732 16548
rect 18788 16492 19068 16548
rect 19124 16492 19134 16548
rect 19506 16492 19516 16548
rect 19572 16492 21644 16548
rect 21700 16492 21924 16548
rect 32844 16548 32900 16604
rect 32844 16492 34300 16548
rect 34356 16492 34366 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 21410 16380 21420 16436
rect 21476 16380 21868 16436
rect 21924 16380 21934 16436
rect 22652 16380 26908 16436
rect 26964 16380 27244 16436
rect 27300 16380 27310 16436
rect 2146 16268 2156 16324
rect 2212 16268 3500 16324
rect 3556 16268 5516 16324
rect 5572 16268 5582 16324
rect 14354 16268 14364 16324
rect 14420 16268 19404 16324
rect 19460 16268 19470 16324
rect 20514 16268 20524 16324
rect 20580 16268 22428 16324
rect 22484 16268 22494 16324
rect 22652 16212 22708 16380
rect 28018 16268 28028 16324
rect 28084 16268 28364 16324
rect 28420 16268 29260 16324
rect 29316 16268 34412 16324
rect 34468 16268 34478 16324
rect 17490 16156 17500 16212
rect 17556 16156 22708 16212
rect 26562 16156 26572 16212
rect 26628 16156 27580 16212
rect 27636 16156 27646 16212
rect 28466 16156 28476 16212
rect 28532 16156 30044 16212
rect 30100 16156 30110 16212
rect 17378 16044 17388 16100
rect 17444 16044 19796 16100
rect 21858 16044 21868 16100
rect 21924 16044 23100 16100
rect 23156 16044 23166 16100
rect 32162 16044 32172 16100
rect 32228 16044 35756 16100
rect 35812 16044 38668 16100
rect 41906 16044 41916 16100
rect 41972 16044 45276 16100
rect 45332 16044 45342 16100
rect 19740 15988 19796 16044
rect 38612 15988 38668 16044
rect 12674 15932 12684 15988
rect 12740 15932 13580 15988
rect 13636 15932 13646 15988
rect 18610 15932 18620 15988
rect 18676 15932 19516 15988
rect 19572 15932 19582 15988
rect 19740 15932 30268 15988
rect 30324 15932 30334 15988
rect 38612 15932 40124 15988
rect 40180 15932 40190 15988
rect 18162 15820 18172 15876
rect 18228 15820 20524 15876
rect 20580 15820 20590 15876
rect 24322 15820 24332 15876
rect 24388 15820 26572 15876
rect 26628 15820 26638 15876
rect 34962 15820 34972 15876
rect 35028 15820 40796 15876
rect 40852 15820 40862 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 23650 15596 23660 15652
rect 23716 15596 25116 15652
rect 25172 15596 32284 15652
rect 32340 15596 33180 15652
rect 33236 15596 33246 15652
rect 9090 15484 9100 15540
rect 9156 15484 10220 15540
rect 10276 15484 11788 15540
rect 11844 15484 11854 15540
rect 16258 15484 16268 15540
rect 16324 15484 16828 15540
rect 16884 15484 17500 15540
rect 17556 15484 17566 15540
rect 20290 15484 20300 15540
rect 20356 15484 22764 15540
rect 22820 15484 22830 15540
rect 28578 15484 28588 15540
rect 28644 15484 29932 15540
rect 29988 15484 31052 15540
rect 31108 15484 31118 15540
rect 33842 15484 33852 15540
rect 33908 15484 37324 15540
rect 37380 15484 37390 15540
rect 37650 15484 37660 15540
rect 37716 15484 38892 15540
rect 38948 15484 38958 15540
rect 37324 15428 37380 15484
rect 15250 15372 15260 15428
rect 15316 15372 24332 15428
rect 24388 15372 24398 15428
rect 26002 15372 26012 15428
rect 26068 15372 27356 15428
rect 27412 15372 29260 15428
rect 29316 15372 29326 15428
rect 37324 15372 38108 15428
rect 38164 15372 39340 15428
rect 39396 15372 39406 15428
rect 5058 15260 5068 15316
rect 5124 15260 5964 15316
rect 6020 15260 6030 15316
rect 12562 15260 12572 15316
rect 12628 15260 25228 15316
rect 25284 15260 25294 15316
rect 26012 15260 26348 15316
rect 26404 15260 26414 15316
rect 30034 15260 30044 15316
rect 30100 15260 30492 15316
rect 30548 15260 30558 15316
rect 35522 15260 35532 15316
rect 35588 15260 35644 15316
rect 35700 15260 35710 15316
rect 26012 15204 26068 15260
rect 1810 15148 1820 15204
rect 1876 15148 3500 15204
rect 3556 15148 3566 15204
rect 7298 15148 7308 15204
rect 7364 15148 8540 15204
rect 8596 15148 8606 15204
rect 9650 15148 9660 15204
rect 9716 15148 14588 15204
rect 14644 15148 14654 15204
rect 19618 15148 19628 15204
rect 19684 15148 20748 15204
rect 20804 15148 20814 15204
rect 26002 15148 26012 15204
rect 26068 15148 26078 15204
rect 37986 15036 37996 15092
rect 38052 15036 38668 15092
rect 38724 15036 41356 15092
rect 41412 15036 41422 15092
rect 19954 14924 19964 14980
rect 20020 14924 21308 14980
rect 21364 14924 22540 14980
rect 22596 14924 22606 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 24210 14812 24220 14868
rect 24276 14812 24892 14868
rect 24948 14812 31724 14868
rect 31780 14812 31790 14868
rect 9874 14700 9884 14756
rect 9940 14700 12572 14756
rect 12628 14700 12638 14756
rect 16818 14700 16828 14756
rect 16884 14700 23212 14756
rect 23268 14700 25452 14756
rect 25508 14700 25518 14756
rect 32050 14700 32060 14756
rect 32116 14700 33852 14756
rect 33908 14700 33918 14756
rect 10546 14588 10556 14644
rect 10612 14588 11900 14644
rect 11956 14588 11966 14644
rect 18274 14588 18284 14644
rect 18340 14588 24108 14644
rect 24164 14588 25004 14644
rect 25060 14588 25900 14644
rect 25956 14588 29148 14644
rect 29204 14588 29214 14644
rect 32610 14588 32620 14644
rect 32676 14588 33292 14644
rect 33348 14588 34860 14644
rect 34916 14588 34926 14644
rect 4834 14476 4844 14532
rect 4900 14476 7980 14532
rect 8036 14476 9548 14532
rect 9604 14476 9614 14532
rect 24770 14476 24780 14532
rect 24836 14476 25788 14532
rect 25844 14476 25854 14532
rect 28466 14476 28476 14532
rect 28532 14476 29484 14532
rect 29540 14476 29550 14532
rect 30258 14476 30268 14532
rect 30324 14476 33180 14532
rect 33236 14476 35532 14532
rect 35588 14476 35598 14532
rect 39330 14476 39340 14532
rect 39396 14476 41132 14532
rect 41188 14476 41198 14532
rect 32386 14364 32396 14420
rect 32452 14364 32956 14420
rect 33012 14364 38668 14420
rect 38612 14308 38668 14364
rect 5618 14252 5628 14308
rect 5684 14252 7196 14308
rect 7252 14252 7262 14308
rect 19730 14252 19740 14308
rect 19796 14252 20188 14308
rect 20244 14252 20254 14308
rect 31154 14252 31164 14308
rect 31220 14252 32284 14308
rect 32340 14252 37772 14308
rect 37828 14252 37838 14308
rect 38612 14252 43148 14308
rect 43204 14252 43214 14308
rect 27794 14140 27804 14196
rect 27860 14140 29484 14196
rect 29540 14140 36988 14196
rect 37044 14140 37054 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 30492 14028 38220 14084
rect 38276 14028 38286 14084
rect 30492 13972 30548 14028
rect 3714 13916 3724 13972
rect 3780 13916 5292 13972
rect 5348 13916 5358 13972
rect 14914 13916 14924 13972
rect 14980 13916 17612 13972
rect 17668 13916 17678 13972
rect 17826 13916 17836 13972
rect 17892 13916 18732 13972
rect 18788 13916 19852 13972
rect 19908 13916 19918 13972
rect 29698 13916 29708 13972
rect 29764 13916 30492 13972
rect 30548 13916 30558 13972
rect 34962 13916 34972 13972
rect 35028 13916 37380 13972
rect 38770 13916 38780 13972
rect 38836 13916 40348 13972
rect 40404 13916 40414 13972
rect 37324 13860 37380 13916
rect 26338 13804 26348 13860
rect 26404 13804 26796 13860
rect 26852 13804 26862 13860
rect 33618 13804 33628 13860
rect 33684 13804 33964 13860
rect 34020 13804 35420 13860
rect 35476 13804 35486 13860
rect 37314 13804 37324 13860
rect 37380 13804 39228 13860
rect 39284 13804 39294 13860
rect 8306 13692 8316 13748
rect 8372 13692 10332 13748
rect 10388 13692 10398 13748
rect 13234 13692 13244 13748
rect 13300 13692 14812 13748
rect 14868 13692 14878 13748
rect 26002 13692 26012 13748
rect 26068 13692 26684 13748
rect 26740 13692 28140 13748
rect 28196 13692 28206 13748
rect 33618 13692 33628 13748
rect 33684 13692 35308 13748
rect 35364 13692 35374 13748
rect 38434 13692 38444 13748
rect 38500 13692 43708 13748
rect 43764 13692 43774 13748
rect 33628 13524 33684 13692
rect 3602 13468 3612 13524
rect 3668 13468 5068 13524
rect 5124 13468 5134 13524
rect 31388 13468 33684 13524
rect 31388 13412 31444 13468
rect 17602 13356 17612 13412
rect 17668 13356 18284 13412
rect 18340 13356 22204 13412
rect 22260 13356 22270 13412
rect 29810 13356 29820 13412
rect 29876 13356 31164 13412
rect 31220 13356 31444 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 13010 13244 13020 13300
rect 13076 13244 13916 13300
rect 13972 13244 29260 13300
rect 29316 13244 29326 13300
rect 39890 13244 39900 13300
rect 39956 13244 40908 13300
rect 40964 13244 40974 13300
rect 15810 13132 15820 13188
rect 15876 13132 16940 13188
rect 16996 13132 17006 13188
rect 26114 13132 26124 13188
rect 26180 13132 26348 13188
rect 26404 13132 26414 13188
rect 31378 13132 31388 13188
rect 31444 13132 32284 13188
rect 32340 13132 34860 13188
rect 34916 13132 35196 13188
rect 35252 13132 35262 13188
rect 14914 13020 14924 13076
rect 14980 13020 16492 13076
rect 16548 13020 20524 13076
rect 20580 13020 20590 13076
rect 13682 12908 13692 12964
rect 13748 12908 14252 12964
rect 14308 12908 15148 12964
rect 15204 12908 15214 12964
rect 16370 12908 16380 12964
rect 16436 12908 18172 12964
rect 18228 12908 18238 12964
rect 19842 12908 19852 12964
rect 19908 12908 20412 12964
rect 20468 12908 20478 12964
rect 23986 12908 23996 12964
rect 24052 12908 26460 12964
rect 26516 12908 26526 12964
rect 18172 12852 18228 12908
rect 26852 12852 26908 12964
rect 26964 12908 26974 12964
rect 31042 12908 31052 12964
rect 31108 12908 31836 12964
rect 31892 12908 31902 12964
rect 32722 12908 32732 12964
rect 32788 12908 33740 12964
rect 33796 12908 33806 12964
rect 37874 12908 37884 12964
rect 37940 12908 38332 12964
rect 38388 12908 38398 12964
rect 38770 12908 38780 12964
rect 38836 12908 40124 12964
rect 40180 12908 40190 12964
rect 43026 12908 43036 12964
rect 43092 12908 45836 12964
rect 45892 12908 45902 12964
rect 12898 12796 12908 12852
rect 12964 12796 14028 12852
rect 14084 12796 15484 12852
rect 15540 12796 15550 12852
rect 18172 12796 21532 12852
rect 21588 12796 21598 12852
rect 22418 12796 22428 12852
rect 22484 12796 26908 12852
rect 29922 12796 29932 12852
rect 29988 12796 30380 12852
rect 30436 12796 32060 12852
rect 32116 12796 32126 12852
rect 37986 12796 37996 12852
rect 38052 12796 38556 12852
rect 38612 12796 38622 12852
rect 1810 12684 1820 12740
rect 1876 12684 3500 12740
rect 3556 12684 3566 12740
rect 6066 12684 6076 12740
rect 6132 12684 7308 12740
rect 7364 12684 8540 12740
rect 8596 12684 8606 12740
rect 17266 12684 17276 12740
rect 17332 12684 17948 12740
rect 18004 12684 18014 12740
rect 23426 12684 23436 12740
rect 23492 12684 25228 12740
rect 25284 12684 26012 12740
rect 26068 12684 26078 12740
rect 31490 12684 31500 12740
rect 31556 12684 32172 12740
rect 32228 12684 32238 12740
rect 33142 12684 33180 12740
rect 33236 12684 33246 12740
rect 30258 12572 30268 12628
rect 30324 12572 30604 12628
rect 30660 12572 32508 12628
rect 32564 12572 33628 12628
rect 33684 12572 33694 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 15092 12348 17948 12404
rect 18004 12348 18014 12404
rect 18162 12348 18172 12404
rect 18228 12348 19852 12404
rect 19908 12348 19918 12404
rect 22194 12348 22204 12404
rect 22260 12348 26348 12404
rect 26404 12348 26414 12404
rect 28242 12348 28252 12404
rect 28308 12348 30268 12404
rect 30324 12348 30334 12404
rect 32498 12348 32508 12404
rect 32564 12348 34076 12404
rect 34132 12348 34142 12404
rect 37874 12348 37884 12404
rect 37940 12348 41804 12404
rect 41860 12348 41870 12404
rect 15092 12292 15148 12348
rect 11554 12236 11564 12292
rect 11620 12236 13468 12292
rect 13524 12236 15148 12292
rect 17042 12236 17052 12292
rect 17108 12236 19292 12292
rect 19348 12236 19358 12292
rect 19506 12236 19516 12292
rect 19572 12236 19740 12292
rect 19796 12236 23324 12292
rect 23380 12236 23390 12292
rect 28466 12236 28476 12292
rect 28532 12236 30940 12292
rect 30996 12236 34860 12292
rect 34916 12236 34926 12292
rect 36642 12236 36652 12292
rect 36708 12236 36988 12292
rect 37044 12236 37660 12292
rect 37716 12236 38668 12292
rect 38724 12236 38734 12292
rect 4050 12124 4060 12180
rect 4116 12124 8876 12180
rect 8932 12124 8942 12180
rect 12338 12124 12348 12180
rect 12404 12124 24332 12180
rect 24388 12124 27020 12180
rect 27076 12124 27086 12180
rect 32162 12124 32172 12180
rect 32228 12124 32844 12180
rect 32900 12124 32910 12180
rect 33170 12124 33180 12180
rect 33236 12124 33628 12180
rect 33684 12124 33694 12180
rect 33842 12124 33852 12180
rect 33908 12124 35532 12180
rect 35588 12124 35598 12180
rect 36530 12124 36540 12180
rect 36596 12124 38108 12180
rect 38164 12124 38444 12180
rect 38500 12124 41804 12180
rect 41860 12124 42364 12180
rect 42420 12124 42430 12180
rect 14466 12012 14476 12068
rect 14532 12012 15372 12068
rect 15428 12012 15438 12068
rect 24546 12012 24556 12068
rect 24612 12012 25228 12068
rect 25284 12012 25294 12068
rect 30146 12012 30156 12068
rect 30212 12012 34412 12068
rect 34468 12012 34478 12068
rect 37202 12012 37212 12068
rect 37268 12012 38556 12068
rect 38612 12012 42700 12068
rect 42756 12012 42766 12068
rect 3714 11900 3724 11956
rect 3780 11900 5404 11956
rect 5460 11900 5470 11956
rect 7970 11900 7980 11956
rect 8036 11900 9548 11956
rect 9604 11900 9614 11956
rect 14354 11900 14364 11956
rect 14420 11900 15036 11956
rect 15092 11900 15260 11956
rect 15316 11900 18172 11956
rect 18228 11900 18238 11956
rect 29586 11900 29596 11956
rect 29652 11900 33068 11956
rect 33124 11900 33404 11956
rect 33460 11900 33470 11956
rect 15474 11788 15484 11844
rect 15540 11788 16380 11844
rect 16436 11788 16446 11844
rect 17714 11788 17724 11844
rect 17780 11788 17948 11844
rect 18004 11788 18014 11844
rect 18386 11788 18396 11844
rect 18452 11788 20076 11844
rect 20132 11788 20142 11844
rect 30258 11788 30268 11844
rect 30324 11788 31164 11844
rect 31220 11788 31230 11844
rect 31826 11788 31836 11844
rect 31892 11788 34972 11844
rect 35028 11788 35038 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 33740 11732 33796 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 11330 11676 11340 11732
rect 11396 11676 12348 11732
rect 12404 11676 12414 11732
rect 12898 11676 12908 11732
rect 12964 11676 20748 11732
rect 20804 11676 20814 11732
rect 33170 11676 33180 11732
rect 33236 11676 33292 11732
rect 33348 11676 33358 11732
rect 33730 11676 33740 11732
rect 33796 11676 33806 11732
rect 3602 11564 3612 11620
rect 3668 11564 5292 11620
rect 5348 11564 5358 11620
rect 9650 11564 9660 11620
rect 9716 11564 11004 11620
rect 11060 11564 11070 11620
rect 19618 11564 19628 11620
rect 19684 11564 21308 11620
rect 21364 11564 21374 11620
rect 1810 11452 1820 11508
rect 1876 11452 3500 11508
rect 3556 11452 8428 11508
rect 8484 11452 8494 11508
rect 24658 11452 24668 11508
rect 24724 11452 26012 11508
rect 26068 11452 27580 11508
rect 27636 11452 27646 11508
rect 27794 11452 27804 11508
rect 27860 11452 29596 11508
rect 29652 11452 29662 11508
rect 32162 11452 32172 11508
rect 32228 11452 33180 11508
rect 33236 11452 33246 11508
rect 4834 11340 4844 11396
rect 4900 11340 5628 11396
rect 5684 11340 6076 11396
rect 6132 11340 6142 11396
rect 12002 11340 12012 11396
rect 12068 11340 13804 11396
rect 13860 11340 13870 11396
rect 15698 11340 15708 11396
rect 15764 11340 16828 11396
rect 16884 11340 16894 11396
rect 23090 11340 23100 11396
rect 23156 11340 24220 11396
rect 24276 11340 24286 11396
rect 30482 11340 30492 11396
rect 30548 11340 31724 11396
rect 31780 11340 31790 11396
rect 10322 11116 10332 11172
rect 10388 11116 10668 11172
rect 10724 11116 12460 11172
rect 12516 11116 12526 11172
rect 22642 11116 22652 11172
rect 22708 11116 29148 11172
rect 29204 11116 29214 11172
rect 32946 11116 32956 11172
rect 33012 11116 33516 11172
rect 33572 11116 41580 11172
rect 41636 11116 42028 11172
rect 42084 11116 42094 11172
rect 13906 11004 13916 11060
rect 13972 11004 14140 11060
rect 14196 11004 14700 11060
rect 14756 11004 14766 11060
rect 22194 11004 22204 11060
rect 22260 11004 23212 11060
rect 23268 11004 23278 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 12226 10780 12236 10836
rect 12292 10780 13468 10836
rect 13524 10780 16716 10836
rect 16772 10780 16782 10836
rect 26226 10668 26236 10724
rect 26292 10668 27804 10724
rect 27860 10668 27870 10724
rect 6066 10556 6076 10612
rect 6132 10556 6636 10612
rect 6692 10556 8428 10612
rect 8484 10556 8494 10612
rect 9090 10556 9100 10612
rect 9156 10556 9996 10612
rect 10052 10556 10062 10612
rect 13906 10556 13916 10612
rect 13972 10556 14924 10612
rect 14980 10556 16044 10612
rect 16100 10556 17388 10612
rect 17444 10556 17454 10612
rect 19954 10556 19964 10612
rect 20020 10556 22204 10612
rect 22260 10556 22270 10612
rect 33394 10556 33404 10612
rect 33460 10556 34524 10612
rect 34580 10556 34590 10612
rect 18162 10444 18172 10500
rect 18228 10444 18508 10500
rect 18564 10444 18574 10500
rect 29250 10444 29260 10500
rect 29316 10444 29596 10500
rect 29652 10444 29662 10500
rect 3714 10332 3724 10388
rect 3780 10332 5180 10388
rect 5236 10332 6188 10388
rect 6244 10332 6254 10388
rect 9874 10332 9884 10388
rect 9940 10332 13132 10388
rect 13188 10332 13198 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19618 10108 19628 10164
rect 19684 10108 20636 10164
rect 20692 10108 24108 10164
rect 24164 10108 25676 10164
rect 25732 10108 25742 10164
rect 2482 9996 2492 10052
rect 2548 9996 4060 10052
rect 4116 9996 4126 10052
rect 13458 9996 13468 10052
rect 13524 9996 14028 10052
rect 14084 9996 14094 10052
rect 16594 9996 16604 10052
rect 16660 9996 17276 10052
rect 17332 9996 17342 10052
rect 23202 9996 23212 10052
rect 23268 9996 24668 10052
rect 24724 9996 24734 10052
rect 21634 9884 21644 9940
rect 21700 9884 23996 9940
rect 24052 9884 24062 9940
rect 31154 9884 31164 9940
rect 31220 9884 31948 9940
rect 32004 9884 32014 9940
rect 4162 9772 4172 9828
rect 4228 9772 5516 9828
rect 5572 9772 5582 9828
rect 20178 9772 20188 9828
rect 20244 9772 21308 9828
rect 21364 9772 21374 9828
rect 31378 9772 31388 9828
rect 31444 9772 32060 9828
rect 32116 9772 33628 9828
rect 33684 9772 33694 9828
rect 34626 9772 34636 9828
rect 34692 9772 39900 9828
rect 39956 9772 39966 9828
rect 2930 9660 2940 9716
rect 2996 9660 4956 9716
rect 5012 9660 5022 9716
rect 12562 9660 12572 9716
rect 12628 9660 16044 9716
rect 16100 9660 17612 9716
rect 17668 9660 17678 9716
rect 23314 9660 23324 9716
rect 23380 9660 25004 9716
rect 25060 9660 25070 9716
rect 2034 9548 2044 9604
rect 2100 9548 4172 9604
rect 4228 9548 4238 9604
rect 16818 9548 16828 9604
rect 16884 9548 17500 9604
rect 17556 9548 18172 9604
rect 18228 9548 20636 9604
rect 20692 9548 20702 9604
rect 38546 9436 38556 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 30930 9212 30940 9268
rect 30996 9212 31724 9268
rect 31780 9212 32060 9268
rect 32116 9212 37436 9268
rect 37492 9212 37502 9268
rect 38612 9156 38668 9492
rect 41570 9212 41580 9268
rect 41636 9212 43372 9268
rect 43428 9212 43438 9268
rect 16146 9100 16156 9156
rect 16212 9100 18620 9156
rect 18676 9100 18686 9156
rect 37538 9100 37548 9156
rect 37604 9100 37614 9156
rect 37874 9100 37884 9156
rect 37940 9100 41244 9156
rect 41300 9100 41310 9156
rect 1922 8988 1932 9044
rect 1988 8988 4844 9044
rect 4900 8988 5964 9044
rect 6020 8988 6030 9044
rect 19954 8988 19964 9044
rect 20020 8988 20636 9044
rect 20692 8988 25228 9044
rect 25284 8988 25294 9044
rect 37548 8932 37604 9100
rect 14466 8876 14476 8932
rect 14532 8876 15148 8932
rect 22082 8876 22092 8932
rect 22148 8876 23324 8932
rect 23380 8876 23390 8932
rect 24994 8876 25004 8932
rect 25060 8876 25676 8932
rect 25732 8876 25742 8932
rect 37548 8876 38556 8932
rect 38612 8876 41580 8932
rect 41636 8876 41646 8932
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 15092 8484 15148 8876
rect 19618 8764 19628 8820
rect 19684 8764 26908 8820
rect 26964 8764 26974 8820
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 24546 8540 24556 8596
rect 24612 8540 25564 8596
rect 25620 8540 26124 8596
rect 26180 8540 26190 8596
rect 15092 8428 16380 8484
rect 16436 8428 17836 8484
rect 17892 8428 21980 8484
rect 22036 8428 22046 8484
rect 29586 8428 29596 8484
rect 29652 8428 30716 8484
rect 30772 8428 33628 8484
rect 33684 8428 33694 8484
rect 16146 8316 16156 8372
rect 16212 8316 17724 8372
rect 17780 8316 17790 8372
rect 24210 8316 24220 8372
rect 24276 8316 24892 8372
rect 24948 8316 27636 8372
rect 30594 8316 30604 8372
rect 30660 8316 31836 8372
rect 31892 8316 35532 8372
rect 35588 8316 35598 8372
rect 14242 8204 14252 8260
rect 14308 8204 15036 8260
rect 15092 8204 15102 8260
rect 15474 8204 15484 8260
rect 15540 8204 18732 8260
rect 18788 8204 18798 8260
rect 25442 8204 25452 8260
rect 25508 8204 26796 8260
rect 26852 8204 27244 8260
rect 27300 8204 27310 8260
rect 27580 8148 27636 8316
rect 29474 8204 29484 8260
rect 29540 8204 31276 8260
rect 31332 8204 31342 8260
rect 31724 8204 35756 8260
rect 35812 8204 35822 8260
rect 31724 8148 31780 8204
rect 25106 8092 25116 8148
rect 25172 8092 27020 8148
rect 27076 8092 27086 8148
rect 27570 8092 27580 8148
rect 27636 8092 27646 8148
rect 30034 8092 30044 8148
rect 30100 8092 30828 8148
rect 30884 8092 31780 8148
rect 31938 8092 31948 8148
rect 32004 8092 32844 8148
rect 32900 8092 34076 8148
rect 34132 8092 34142 8148
rect 18834 7980 18844 8036
rect 18900 7980 20636 8036
rect 20692 7980 23884 8036
rect 23940 7980 23950 8036
rect 24668 7980 26908 8036
rect 26964 7980 26974 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 24668 7812 24724 7980
rect 20402 7756 20412 7812
rect 20468 7756 21308 7812
rect 21364 7756 24668 7812
rect 24724 7756 24734 7812
rect 22978 7644 22988 7700
rect 23044 7644 26796 7700
rect 26852 7644 26862 7700
rect 21410 7420 21420 7476
rect 21476 7420 22876 7476
rect 22932 7420 22942 7476
rect 28354 7420 28364 7476
rect 28420 7420 29484 7476
rect 29540 7420 29550 7476
rect 33954 7420 33964 7476
rect 34020 7420 36204 7476
rect 36260 7420 36270 7476
rect 21298 7308 21308 7364
rect 21364 7308 21532 7364
rect 21588 7308 23436 7364
rect 23492 7308 23502 7364
rect 30146 7308 30156 7364
rect 30212 7308 34860 7364
rect 34916 7308 35644 7364
rect 35700 7308 35710 7364
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 4274 6860 4284 6916
rect 4340 6860 5852 6916
rect 5908 6860 5918 6916
rect 27570 6748 27580 6804
rect 27636 6748 28364 6804
rect 28420 6748 28430 6804
rect 19170 6636 19180 6692
rect 19236 6636 21644 6692
rect 21700 6636 21710 6692
rect 24434 6636 24444 6692
rect 24500 6636 25340 6692
rect 25396 6636 25406 6692
rect 28578 6636 28588 6692
rect 28644 6636 29148 6692
rect 29204 6636 30156 6692
rect 30212 6636 30222 6692
rect 18274 6412 18284 6468
rect 18340 6412 20524 6468
rect 20580 6412 20590 6468
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 18498 6076 18508 6132
rect 18564 6076 18956 6132
rect 19012 6076 20188 6132
rect 20244 6076 20972 6132
rect 21028 6076 21038 6132
rect 19842 5964 19852 6020
rect 19908 5964 21308 6020
rect 21364 5964 21374 6020
rect 18610 5852 18620 5908
rect 18676 5852 19292 5908
rect 19348 5852 19358 5908
rect 21186 5852 21196 5908
rect 21252 5852 22204 5908
rect 22260 5852 22270 5908
rect 24770 5852 24780 5908
rect 24836 5852 25676 5908
rect 25732 5852 25742 5908
rect 20850 5740 20860 5796
rect 20916 5740 21756 5796
rect 21812 5740 21822 5796
rect 23426 5740 23436 5796
rect 23492 5740 25228 5796
rect 25284 5740 25294 5796
rect 19170 5628 19180 5684
rect 19236 5628 22092 5684
rect 22148 5628 22876 5684
rect 22932 5628 22942 5684
rect 24098 5628 24108 5684
rect 24164 5628 25452 5684
rect 25508 5628 25518 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 20290 5180 20300 5236
rect 20356 5180 21420 5236
rect 21476 5180 21486 5236
rect 19058 5068 19068 5124
rect 19124 5068 21532 5124
rect 21588 5068 21598 5124
rect 21644 4956 22316 5012
rect 22372 4956 23100 5012
rect 23156 4956 23884 5012
rect 23940 4956 23950 5012
rect 1698 4844 1708 4900
rect 1764 4844 1774 4900
rect 0 4788 800 4816
rect 1708 4788 1764 4844
rect 21644 4788 21700 4956
rect 0 4732 1764 4788
rect 21634 4732 21644 4788
rect 21700 4732 21710 4788
rect 0 4704 800 4732
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 16706 4508 16716 4564
rect 16772 4508 19740 4564
rect 19796 4508 19806 4564
rect 18610 4060 18620 4116
rect 18676 4060 19516 4116
rect 19572 4060 21196 4116
rect 21252 4060 21262 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 16268 36988 16324 37044
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 22652 34972 22708 35028
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 22652 34188 22708 34244
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 28588 29708 28644 29764
rect 28588 29036 28644 29092
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 15708 23436 15764 23492
rect 20524 23436 20580 23492
rect 25788 23212 25844 23268
rect 22204 23100 22260 23156
rect 15708 22764 15764 22820
rect 23212 22764 23268 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 25788 22092 25844 22148
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 28588 21532 28644 21588
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 22204 20524 22260 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 16268 18060 16324 18116
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 20412 17836 20468 17892
rect 35644 17500 35700 17556
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 20412 16716 20468 16772
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 20524 15820 20580 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 35644 15260 35700 15316
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 23212 14700 23268 14756
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 33628 13804 33684 13860
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 33180 12684 33236 12740
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 33628 12124 33684 12180
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 33180 11676 33236 11732
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 44716 4768 44748
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 19808 43932 20128 44748
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 16268 37044 16324 37054
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 15708 23492 15764 23502
rect 15708 22820 15764 23436
rect 15708 22754 15764 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 16268 18116 16324 36988
rect 16268 18050 16324 18060
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 35168 44716 35488 44748
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 22652 35028 22708 35038
rect 22652 34244 22708 34972
rect 22652 34178 22708 34188
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 28588 29764 28644 29774
rect 28588 29092 28644 29708
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 17276 20128 18788
rect 20524 23492 20580 23502
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 20412 17892 20468 17902
rect 20412 16772 20468 17836
rect 20412 16706 20468 16716
rect 20524 15876 20580 23436
rect 25788 23268 25844 23278
rect 22204 23156 22260 23166
rect 22204 20580 22260 23100
rect 22204 20514 22260 20524
rect 23212 22820 23268 22830
rect 20524 15810 20580 15820
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 23212 14756 23268 22764
rect 25788 22148 25844 23212
rect 25788 22082 25844 22092
rect 28588 21588 28644 29036
rect 28588 21522 28644 21532
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 23212 14690 23268 14700
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35644 17556 35700 17566
rect 35644 15316 35700 17500
rect 35644 15250 35700 15260
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 33628 13860 33684 13870
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 33180 12740 33236 12750
rect 33180 11732 33236 12684
rect 33628 12180 33684 13804
rect 33628 12114 33684 12124
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 33180 11666 33236 11676
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _243_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18816 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _244_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27440 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _245_
timestamp 1698431365
transform -1 0 22848 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _246_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34608 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _247_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33600 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _248_
timestamp 1698431365
transform -1 0 34832 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _249_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34048 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _250_
timestamp 1698431365
transform 1 0 34160 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _251_
timestamp 1698431365
transform 1 0 41776 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _252_
timestamp 1698431365
transform 1 0 29120 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _253_
timestamp 1698431365
transform 1 0 23184 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _254_
timestamp 1698431365
transform 1 0 24864 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _255_
timestamp 1698431365
transform 1 0 29120 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _256_
timestamp 1698431365
transform 1 0 29120 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _257_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22400 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _258_
timestamp 1698431365
transform 1 0 24192 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _259_
timestamp 1698431365
transform 1 0 31248 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _260_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24864 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _261_
timestamp 1698431365
transform 1 0 30576 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _262_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26768 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _263_
timestamp 1698431365
transform -1 0 19376 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _264_
timestamp 1698431365
transform 1 0 23632 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _265_
timestamp 1698431365
transform 1 0 35168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _266_
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _267_
timestamp 1698431365
transform 1 0 25088 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _268_
timestamp 1698431365
transform 1 0 39760 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _269_
timestamp 1698431365
transform 1 0 28000 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _270_
timestamp 1698431365
transform 1 0 38304 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _271_
timestamp 1698431365
transform 1 0 31920 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _272_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38528 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _273_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _274_
timestamp 1698431365
transform 1 0 17472 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _275_
timestamp 1698431365
transform -1 0 23856 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _276_
timestamp 1698431365
transform -1 0 21952 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _277_
timestamp 1698431365
transform -1 0 22064 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _278_
timestamp 1698431365
transform 1 0 17472 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _279_
timestamp 1698431365
transform 1 0 18816 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _280_
timestamp 1698431365
transform 1 0 23520 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _281_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21952 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _282_
timestamp 1698431365
transform 1 0 22400 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _283_
timestamp 1698431365
transform 1 0 21504 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _284_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22736 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _285_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22400 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _286_
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _287_
timestamp 1698431365
transform 1 0 19824 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _288_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21392 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _289_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20720 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _290_
timestamp 1698431365
transform -1 0 11984 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _291_
timestamp 1698431365
transform 1 0 10528 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _292_
timestamp 1698431365
transform -1 0 12992 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _293_
timestamp 1698431365
transform 1 0 17584 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _294_
timestamp 1698431365
transform 1 0 24080 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _295_
timestamp 1698431365
transform -1 0 24864 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _296_
timestamp 1698431365
transform -1 0 22624 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _297_
timestamp 1698431365
transform -1 0 19152 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _298_
timestamp 1698431365
transform 1 0 15008 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _299_
timestamp 1698431365
transform -1 0 20160 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _300_
timestamp 1698431365
transform -1 0 23744 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _301_
timestamp 1698431365
transform -1 0 20832 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _302_
timestamp 1698431365
transform -1 0 24080 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _303_
timestamp 1698431365
transform -1 0 19936 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _304_
timestamp 1698431365
transform -1 0 24192 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _305_
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _306_
timestamp 1698431365
transform -1 0 28000 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _307_
timestamp 1698431365
transform 1 0 23520 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _308_
timestamp 1698431365
transform 1 0 26656 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _309_
timestamp 1698431365
transform 1 0 23968 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _310_
timestamp 1698431365
transform -1 0 26880 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _311_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _312_
timestamp 1698431365
transform -1 0 26320 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _313_
timestamp 1698431365
transform 1 0 24304 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _314_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26096 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _315_
timestamp 1698431365
transform 1 0 20160 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _316_
timestamp 1698431365
transform -1 0 24304 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _317_
timestamp 1698431365
transform 1 0 23744 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _318_
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _319_
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _320_
timestamp 1698431365
transform 1 0 21840 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _321_
timestamp 1698431365
transform 1 0 26656 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _322_
timestamp 1698431365
transform -1 0 23520 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _323_
timestamp 1698431365
transform 1 0 25312 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _324_
timestamp 1698431365
transform 1 0 22176 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _325_
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _326_
timestamp 1698431365
transform 1 0 19936 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _327_
timestamp 1698431365
transform 1 0 19712 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _328_
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _329_
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _330_
timestamp 1698431365
transform -1 0 20160 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _331_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19376 0 -1 25088
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _332_
timestamp 1698431365
transform 1 0 7504 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _333_
timestamp 1698431365
transform -1 0 7504 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _334_
timestamp 1698431365
transform 1 0 32928 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _335_
timestamp 1698431365
transform -1 0 37408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _336_
timestamp 1698431365
transform 1 0 40320 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _337_
timestamp 1698431365
transform 1 0 34832 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _338_
timestamp 1698431365
transform 1 0 38640 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_2  _339_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _340_
timestamp 1698431365
transform 1 0 38864 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _341_
timestamp 1698431365
transform 1 0 26992 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _342_
timestamp 1698431365
transform 1 0 24752 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _343_
timestamp 1698431365
transform 1 0 25872 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _344_
timestamp 1698431365
transform -1 0 21056 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _345_
timestamp 1698431365
transform -1 0 23072 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _346_
timestamp 1698431365
transform 1 0 21056 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _347_
timestamp 1698431365
transform 1 0 24304 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _348_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25760 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _349_
timestamp 1698431365
transform -1 0 26992 0 -1 25088
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _350_
timestamp 1698431365
transform 1 0 41664 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _351_
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _352_
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _353_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23408 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _354_
timestamp 1698431365
transform -1 0 20720 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _355_
timestamp 1698431365
transform 1 0 23184 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _356_
timestamp 1698431365
transform 1 0 22288 0 -1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _357_
timestamp 1698431365
transform 1 0 23184 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _358_
timestamp 1698431365
transform 1 0 7392 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _359_
timestamp 1698431365
transform 1 0 6160 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _360_
timestamp 1698431365
transform 1 0 21280 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _361_
timestamp 1698431365
transform 1 0 23856 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _362_
timestamp 1698431365
transform -1 0 23968 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _363_
timestamp 1698431365
transform 1 0 30016 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _364_
timestamp 1698431365
transform -1 0 28896 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _365_
timestamp 1698431365
transform 1 0 31808 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _366_
timestamp 1698431365
transform 1 0 29120 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _367_
timestamp 1698431365
transform -1 0 28336 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _368_
timestamp 1698431365
transform 1 0 24864 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _369_
timestamp 1698431365
transform -1 0 27440 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _370_
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _371_
timestamp 1698431365
transform 1 0 14672 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _372_
timestamp 1698431365
transform 1 0 14448 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _373_
timestamp 1698431365
transform -1 0 18928 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _374_
timestamp 1698431365
transform -1 0 17248 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _375_
timestamp 1698431365
transform 1 0 11424 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _376_
timestamp 1698431365
transform -1 0 20944 0 1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _377_
timestamp 1698431365
transform -1 0 20720 0 1 25088
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _378_
timestamp 1698431365
transform -1 0 10304 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _379_
timestamp 1698431365
transform 1 0 5600 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _380_
timestamp 1698431365
transform -1 0 5264 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _381_
timestamp 1698431365
transform 1 0 31584 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _382_
timestamp 1698431365
transform 1 0 33040 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _383_
timestamp 1698431365
transform -1 0 34608 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _384_
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _385_
timestamp 1698431365
transform -1 0 24304 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _386_
timestamp 1698431365
transform 1 0 22736 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _387_
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _388_
timestamp 1698431365
transform 1 0 25200 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _389_
timestamp 1698431365
transform -1 0 26656 0 1 23520
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _390_
timestamp 1698431365
transform 1 0 39648 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _391_
timestamp 1698431365
transform 1 0 32816 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _392_
timestamp 1698431365
transform 1 0 33600 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _393_
timestamp 1698431365
transform 1 0 22400 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _394_
timestamp 1698431365
transform 1 0 22064 0 1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _395_
timestamp 1698431365
transform 1 0 22624 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _396_
timestamp 1698431365
transform 1 0 5712 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _397_
timestamp 1698431365
transform 1 0 4592 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _398_
timestamp 1698431365
transform 1 0 15904 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _399_
timestamp 1698431365
transform 1 0 18368 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _400_
timestamp 1698431365
transform -1 0 20608 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_2  _401_
timestamp 1698431365
transform 1 0 39424 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _402_
timestamp 1698431365
transform -1 0 27664 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _403_
timestamp 1698431365
transform 1 0 25200 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _404_
timestamp 1698431365
transform -1 0 26544 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _405_
timestamp 1698431365
transform 1 0 26096 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _406_
timestamp 1698431365
transform 1 0 20048 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _407_
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _408_
timestamp 1698431365
transform 1 0 22288 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _409_
timestamp 1698431365
transform 1 0 22624 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _410_
timestamp 1698431365
transform -1 0 20272 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _411_
timestamp 1698431365
transform 1 0 19712 0 -1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _412_
timestamp 1698431365
transform 1 0 19040 0 1 23520
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _413_
timestamp 1698431365
transform 1 0 6048 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _414_
timestamp 1698431365
transform -1 0 8736 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _415_
timestamp 1698431365
transform 1 0 35168 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _416_
timestamp 1698431365
transform 1 0 35392 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _417_
timestamp 1698431365
transform 1 0 34832 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _418_
timestamp 1698431365
transform 1 0 27552 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _419_
timestamp 1698431365
transform -1 0 27440 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _420_
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _421_
timestamp 1698431365
transform 1 0 22960 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _422_
timestamp 1698431365
transform 1 0 24864 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _423_
timestamp 1698431365
transform -1 0 26992 0 -1 26656
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _424_
timestamp 1698431365
transform 1 0 40880 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _425_
timestamp 1698431365
transform 1 0 35728 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _426_
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _427_
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _428_
timestamp 1698431365
transform 1 0 19712 0 -1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _429_
timestamp 1698431365
transform 1 0 18144 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _430_
timestamp 1698431365
transform -1 0 9856 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _431_
timestamp 1698431365
transform -1 0 10752 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _432_
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _433_
timestamp 1698431365
transform 1 0 25648 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _434_
timestamp 1698431365
transform -1 0 23632 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _435_
timestamp 1698431365
transform 1 0 29120 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _436_
timestamp 1698431365
transform -1 0 28224 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _437_
timestamp 1698431365
transform 1 0 34944 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _438_
timestamp 1698431365
transform -1 0 27664 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _439_
timestamp 1698431365
transform -1 0 27440 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _440_
timestamp 1698431365
transform 1 0 21728 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _441_
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _442_
timestamp 1698431365
transform 1 0 16016 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _443_
timestamp 1698431365
transform -1 0 19040 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _444_
timestamp 1698431365
transform -1 0 18928 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _445_
timestamp 1698431365
transform -1 0 23744 0 1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _446_
timestamp 1698431365
transform -1 0 23184 0 -1 25088
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _447_
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _448_
timestamp 1698431365
transform -1 0 10080 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _449_
timestamp 1698431365
transform 1 0 9520 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _450_
timestamp 1698431365
transform 1 0 9520 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _451_
timestamp 1698431365
transform 1 0 9296 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _452_
timestamp 1698431365
transform -1 0 9072 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _453_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _454_
timestamp 1698431365
transform -1 0 18368 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _455_
timestamp 1698431365
transform -1 0 18816 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _456_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14000 0 1 18816
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _457_
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _458_
timestamp 1698431365
transform -1 0 17920 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _459_
timestamp 1698431365
transform -1 0 13440 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _460_
timestamp 1698431365
transform -1 0 17024 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _461_
timestamp 1698431365
transform -1 0 15008 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _462_
timestamp 1698431365
transform 1 0 13776 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _463_
timestamp 1698431365
transform -1 0 14000 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _464_
timestamp 1698431365
transform -1 0 14896 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _465_
timestamp 1698431365
transform -1 0 13216 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _466_
timestamp 1698431365
transform 1 0 10192 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _467_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15568 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _468_
timestamp 1698431365
transform 1 0 12432 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _469_
timestamp 1698431365
transform -1 0 16240 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _470_
timestamp 1698431365
transform -1 0 17808 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _471_
timestamp 1698431365
transform -1 0 16576 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _472_
timestamp 1698431365
transform 1 0 12208 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _473_
timestamp 1698431365
transform 1 0 10864 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _474_
timestamp 1698431365
transform 1 0 10080 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _475_
timestamp 1698431365
transform 1 0 11312 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _476_
timestamp 1698431365
transform -1 0 11424 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _477_
timestamp 1698431365
transform 1 0 10864 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _478_
timestamp 1698431365
transform 1 0 8512 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _479_
timestamp 1698431365
transform 1 0 14672 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _480_
timestamp 1698431365
transform 1 0 17024 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _481_
timestamp 1698431365
transform -1 0 13888 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _482_
timestamp 1698431365
transform 1 0 12656 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _483_
timestamp 1698431365
transform -1 0 18704 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _484_
timestamp 1698431365
transform 1 0 13888 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _485_
timestamp 1698431365
transform 1 0 12208 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _486_
timestamp 1698431365
transform -1 0 13552 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _487_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _488_
timestamp 1698431365
transform 1 0 10304 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _489_
timestamp 1698431365
transform -1 0 9072 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _490_
timestamp 1698431365
transform 1 0 10416 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _491_
timestamp 1698431365
transform 1 0 7840 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _492_
timestamp 1698431365
transform 1 0 10752 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _493_
timestamp 1698431365
transform -1 0 10080 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _494_ test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17024 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _495_
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _496_
timestamp 1698431365
transform 1 0 13888 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _497_
timestamp 1698431365
transform 1 0 16240 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _498_
timestamp 1698431365
transform 1 0 15568 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _499_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _500_
timestamp 1698431365
transform -1 0 12880 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _501_
timestamp 1698431365
transform 1 0 10192 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _502_
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _503_
timestamp 1698431365
transform -1 0 17024 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _504_
timestamp 1698431365
transform -1 0 16688 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _505_
timestamp 1698431365
transform 1 0 13888 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _506_
timestamp 1698431365
transform 1 0 9072 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _507_
timestamp 1698431365
transform 1 0 7056 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _508_
timestamp 1698431365
transform 1 0 8064 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _509_
timestamp 1698431365
transform 1 0 7504 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__I test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__I
timestamp 1698431365
transform -1 0 33600 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__I
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__I
timestamp 1698431365
transform 1 0 22960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__I
timestamp 1698431365
transform -1 0 29456 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__I
timestamp 1698431365
transform -1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__S1
timestamp 1698431365
transform -1 0 41216 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__I
timestamp 1698431365
transform 1 0 31696 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__272__S
timestamp 1698431365
transform -1 0 37408 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__I
timestamp 1698431365
transform 1 0 23632 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__I
timestamp 1698431365
transform 1 0 18704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__I
timestamp 1698431365
transform 1 0 18592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__I
timestamp 1698431365
transform -1 0 22736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__288__A2
timestamp 1698431365
transform 1 0 24304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__S0
timestamp 1698431365
transform -1 0 18816 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__S1
timestamp 1698431365
transform -1 0 18256 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__I
timestamp 1698431365
transform 1 0 20384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__I
timestamp 1698431365
transform 1 0 24080 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__323__S
timestamp 1698431365
transform 1 0 26544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__326__A1
timestamp 1698431365
transform 1 0 18144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__S0
timestamp 1698431365
transform 1 0 40096 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__I
timestamp 1698431365
transform 1 0 33936 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__S
timestamp 1698431365
transform -1 0 39760 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__I
timestamp 1698431365
transform 1 0 27888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__S0
timestamp 1698431365
transform 1 0 41888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__A1
timestamp 1698431365
transform 1 0 22624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__S
timestamp 1698431365
transform 1 0 19152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__374__I
timestamp 1698431365
transform -1 0 16352 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__381__S1
timestamp 1698431365
transform -1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__S
timestamp 1698431365
transform -1 0 31808 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__S1
timestamp 1698431365
transform -1 0 39536 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__S
timestamp 1698431365
transform 1 0 34944 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__S0
timestamp 1698431365
transform 1 0 21504 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__S1
timestamp 1698431365
transform 1 0 20608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__S
timestamp 1698431365
transform 1 0 24528 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__415__S0
timestamp 1698431365
transform 1 0 35728 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__S0
timestamp 1698431365
transform 1 0 25312 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__424__S0
timestamp 1698431365
transform 1 0 40992 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__428__A2
timestamp 1698431365
transform 1 0 23968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__442__S0
timestamp 1698431365
transform 1 0 19824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__S
timestamp 1698431365
transform 1 0 19264 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__I1
timestamp 1698431365
transform 1 0 12768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__479__A2
timestamp 1698431365
transform 1 0 14448 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__A2
timestamp 1698431365
transform 1 0 15232 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__483__A2
timestamp 1698431365
transform 1 0 17920 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__CLK
timestamp 1698431365
transform 1 0 13664 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__497__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__CLK
timestamp 1698431365
transform 1 0 15344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__499__CLK
timestamp 1698431365
transform 1 0 18032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.and3_2_inst_A3
timestamp 1698431365
transform 1 0 26432 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_1_inst_A4
timestamp 1698431365
transform -1 0 31136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.and4_4_inst_A3
timestamp 1698431365
transform 1 0 21952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi22_1_inst_B2
timestamp 1698431365
transform -1 0 29120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_4_inst_B2
timestamp 1698431365
transform 1 0 24976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.aoi221_4_inst_C
timestamp 1698431365
transform -1 0 24752 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_3_inst_EN
timestamp 1698431365
transform -1 0 16800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.bufz_3_inst_I
timestamp 1698431365
transform 1 0 16464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.dffnrsnq_2_inst_SETN
timestamp 1698431365
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtn_1_inst_TE
timestamp 1698431365
transform 1 0 19600 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_2_inst_TE
timestamp 1698431365
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.icgtp_4_inst_TE
timestamp 1698431365
transform 1 0 15904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_1_inst_A2
timestamp 1698431365
transform -1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.nand3_1_inst_A3
timestamp 1698431365
transform -1 0 28336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai22_2_inst_B2
timestamp 1698431365
transform 1 0 24080 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai31_4_inst_B
timestamp 1698431365
transform 1 0 22176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_B1
timestamp 1698431365
transform 1 0 25312 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_B2
timestamp 1698431365
transform 1 0 24304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_1_inst_B3
timestamp 1698431365
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.oai33_2_inst_B2
timestamp 1698431365
transform 1 0 33936 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrnq_2_inst_SI
timestamp 1698431365
transform -1 0 18592 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SETN
timestamp 1698431365
transform -1 0 34832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_1_inst_SI
timestamp 1698431365
transform -1 0 27776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SETN
timestamp 1698431365
transform 1 0 22064 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffrsnq_4_inst_SI
timestamp 1698431365
transform 1 0 21728 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_cm_inst.cc_inst.sdffsnq_2_inst_SI
timestamp 1698431365
transform -1 0 27216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout17_I
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout18_I
timestamp 1698431365
transform 1 0 36736 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout19_I
timestamp 1698431365
transform 1 0 36400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout21_I
timestamp 1698431365
transform 1 0 39536 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout22_I
timestamp 1698431365
transform 1 0 35840 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout24_I
timestamp 1698431365
transform 1 0 17360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout25_I
timestamp 1698431365
transform -1 0 19152 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout28_I
timestamp 1698431365
transform -1 0 31024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout29_I
timestamp 1698431365
transform 1 0 35616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout30_I
timestamp 1698431365
transform 1 0 37520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout31_I
timestamp 1698431365
transform 1 0 40320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout32_I
timestamp 1698431365
transform 1 0 32592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout33_I
timestamp 1698431365
transform -1 0 36512 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout34_I
timestamp 1698431365
transform 1 0 42336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout35_I
timestamp 1698431365
transform 1 0 40992 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout36_I
timestamp 1698431365
transform 1 0 35504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout39_I
timestamp 1698431365
transform 1 0 17584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout40_I
timestamp 1698431365
transform -1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout41_I
timestamp 1698431365
transform -1 0 14224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout51_I
timestamp 1698431365
transform -1 0 31808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout58_I
timestamp 1698431365
transform -1 0 15680 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout59_I
timestamp 1698431365
transform 1 0 39648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout60_I
timestamp 1698431365
transform 1 0 41552 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout68_I
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout78_I
timestamp 1698431365
transform -1 0 11872 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout79_I
timestamp 1698431365
transform 1 0 27216 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout80_I
timestamp 1698431365
transform -1 0 10752 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout81_I
timestamp 1698431365
transform -1 0 11760 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout98_I
timestamp 1698431365
transform 1 0 28336 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout101_I
timestamp 1698431365
transform -1 0 13888 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout110_I
timestamp 1698431365
transform -1 0 17696 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout113_I
timestamp 1698431365
transform -1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout116_I
timestamp 1698431365
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout117_I
timestamp 1698431365
transform 1 0 36960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout126_I
timestamp 1698431365
transform 1 0 34272 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout163_I
timestamp 1698431365
transform -1 0 13776 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout181_I
timestamp 1698431365
transform 1 0 16800 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout184_I
timestamp 1698431365
transform -1 0 27552 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout187_I
timestamp 1698431365
transform 1 0 40208 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout188_I
timestamp 1698431365
transform 1 0 44912 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout198_I
timestamp 1698431365
transform 1 0 33600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout199_I
timestamp 1698431365
transform -1 0 14560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout223_I
timestamp 1698431365
transform -1 0 9744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout245_I
timestamp 1698431365
transform -1 0 29456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout246_I
timestamp 1698431365
transform -1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout267_I
timestamp 1698431365
transform -1 0 11424 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout283_I
timestamp 1698431365
transform -1 0 27888 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout284_I
timestamp 1698431365
transform -1 0 28000 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout289_I
timestamp 1698431365
transform 1 0 39872 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout291_I
timestamp 1698431365
transform 1 0 33824 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout292_I
timestamp 1698431365
transform 1 0 11536 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout304_I
timestamp 1698431365
transform -1 0 8176 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout312_I
timestamp 1698431365
transform 1 0 3584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout313_I
timestamp 1698431365
transform -1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 1792 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 4592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 2688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 6384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 2240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 6608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 3360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cells7_316 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cells7_317
timestamp 1698431365
transform -1 0 2016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cells7_318
timestamp 1698431365
transform 1 0 45920 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cells7_319
timestamp 1698431365
transform -1 0 2016 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__addf_1  cm_inst.cc_inst.addf_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42000 0 -1 23520
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__addf_2  cm_inst.cc_inst.addf_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30688 0 1 17248
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__addf_4  cm_inst.cc_inst.addf_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37184 0 1 28224
box -86 -86 5014 870
use gf180mcu_fd_sc_mcu7t5v0__addh_1  cm_inst.cc_inst.addh_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__addh_2  cm_inst.cc_inst.addh_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38192 0 1 23520
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__addh_4  cm_inst.cc_inst.addh_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27440 0 -1 17248
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  cm_inst.cc_inst.and2_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25984 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  cm_inst.cc_inst.and2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22848 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  cm_inst.cc_inst.and2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22848 0 1 29792
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  cm_inst.cc_inst.and3_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  cm_inst.cc_inst.and3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25984 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_4  cm_inst.cc_inst.and3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24416 0 1 7840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  cm_inst.cc_inst.and4_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29456 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  cm_inst.cc_inst.and4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15568 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and4_4  cm_inst.cc_inst.and4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22176 0 -1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  cm_inst.cc_inst.aoi21_1_inst
timestamp 1698431365
transform -1 0 43680 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  cm_inst.cc_inst.aoi21_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  cm_inst.cc_inst.aoi21_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35168 0 -1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  cm_inst.cc_inst.aoi22_1_inst
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  cm_inst.cc_inst.aoi22_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39648 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  cm_inst.cc_inst.aoi22_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  cm_inst.cc_inst.aoi211_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  cm_inst.cc_inst.aoi211_2_inst
timestamp 1698431365
transform -1 0 28224 0 1 12544
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  cm_inst.cc_inst.aoi211_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 44464 0 1 37632
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  cm_inst.cc_inst.aoi221_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31696 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  cm_inst.cc_inst.aoi221_2_inst
timestamp 1698431365
transform 1 0 34384 0 -1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  cm_inst.cc_inst.aoi221_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25760 0 -1 15680
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  cm_inst.cc_inst.aoi222_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  cm_inst.cc_inst.aoi222_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 36624 0 1 18816
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  cm_inst.cc_inst.aoi222_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39200 0 1 29792
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  cm_inst.cc_inst.buf_1_inst
timestamp 1698431365
transform -1 0 29344 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  cm_inst.cc_inst.buf_2_inst
timestamp 1698431365
transform -1 0 28112 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  cm_inst.cc_inst.buf_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30128 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  cm_inst.cc_inst.buf_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  cm_inst.cc_inst.buf_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29344 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  cm_inst.cc_inst.buf_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26544 0 -1 6272
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__buf_16  cm_inst.cc_inst.buf_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_20  cm_inst.cc_inst.buf_20_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7030 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_1  cm_inst.cc_inst.bufz_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_2  cm_inst.cc_inst.bufz_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14112 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_3  cm_inst.cc_inst.bufz_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14112 0 -1 39200
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_4  cm_inst.cc_inst.bufz_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43344 0 -1 17248
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_8  cm_inst.cc_inst.bufz_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42560 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_12  cm_inst.cc_inst.bufz_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41216 0 -1 15680
box -86 -86 5238 870
use gf180mcu_fd_sc_mcu7t5v0__bufz_16  cm_inst.cc_inst.bufz_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 6582 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  cm_inst.cc_inst.clkbuf_1_inst
timestamp 1698431365
transform -1 0 41440 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  cm_inst.cc_inst.clkbuf_2_inst
timestamp 1698431365
transform 1 0 31136 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  cm_inst.cc_inst.clkbuf_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42896 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  cm_inst.cc_inst.clkbuf_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  cm_inst.cc_inst.clkbuf_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_12  cm_inst.cc_inst.clkbuf_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19040 0 -1 14112
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  cm_inst.cc_inst.clkbuf_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22064 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_20  cm_inst.cc_inst.clkbuf_20_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 7030 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  cm_inst.cc_inst.clkinv_1_inst
timestamp 1698431365
transform -1 0 24752 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  cm_inst.cc_inst.clkinv_2_inst
timestamp 1698431365
transform -1 0 19600 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  cm_inst.cc_inst.clkinv_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19824 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  cm_inst.cc_inst.clkinv_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_8  cm_inst.cc_inst.clkinv_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22288 0 -1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_12  cm_inst.cc_inst.clkinv_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22736 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_16  cm_inst.cc_inst.clkinv_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23072 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_20  cm_inst.cc_inst.clkinv_20_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9856 0 -1 31360
box -86 -86 4790 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  cm_inst.cc_inst.dffnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_2  cm_inst.cc_inst.dffnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37632 0 1 7840
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_4  cm_inst.cc_inst.dffnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25648 0 -1 42336
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  cm_inst.cc_inst.dffnrnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34944 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2  cm_inst.cc_inst.dffnrnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10528 0 -1 37632
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4  cm_inst.cc_inst.dffnrnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31136 0 1 7840
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1  cm_inst.cc_inst.dffnrsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19488 0 -1 42336
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2  cm_inst.cc_inst.dffnrsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 5126 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4  cm_inst.cc_inst.dffnrsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 5574 870
use gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1  cm_inst.cc_inst.dffnsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34608 0 -1 9408
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2  cm_inst.cc_inst.dffnsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22624 0 1 42336
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4  cm_inst.cc_inst.dffnsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31696 0 1 37632
box -86 -86 4790 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  cm_inst.cc_inst.dffq_1_inst
timestamp 1698431365
transform 1 0 9856 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  cm_inst.cc_inst.dffq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29232 0 -1 7840
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  cm_inst.cc_inst.dffq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18928 0 -1 43904
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  cm_inst.cc_inst.dffrnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31808 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  cm_inst.cc_inst.dffrnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10752 0 -1 34496
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_4  cm_inst.cc_inst.dffrnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35616 0 -1 7840
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1  cm_inst.cc_inst.dffrsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23408 0 1 40768
box -86 -86 4454 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2  cm_inst.cc_inst.dffrsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 4678 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4  cm_inst.cc_inst.dffrsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9968 0 -1 36064
box -86 -86 5126 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  cm_inst.cc_inst.dffsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_2  cm_inst.cc_inst.dffsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19152 0 -1 40768
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_4  cm_inst.cc_inst.dffsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31808 0 1 31360
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_1  cm_inst.cc_inst.dlya_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38528 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  cm_inst.cc_inst.dlya_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27328 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_4  cm_inst.cc_inst.dlya_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42336 0 1 20384
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  cm_inst.cc_inst.dlyb_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12320 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_2  cm_inst.cc_inst.dlyb_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37856 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_4  cm_inst.cc_inst.dlyb_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27216 0 -1 39200
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  cm_inst.cc_inst.dlyc_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38080 0 1 32928
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_2  cm_inst.cc_inst.dlyc_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11088 0 -1 39200
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_4  cm_inst.cc_inst.dlyc_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37072 0 -1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dlyd_1  cm_inst.cc_inst.dlyd_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26208 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dlyd_2  cm_inst.cc_inst.dlyd_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38864 0 1 17248
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dlyd_4  cm_inst.cc_inst.dlyd_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8624 0 1 39200
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__hold  cm_inst.cc_inst.hold_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__icgtn_1  cm_inst.cc_inst.icgtn_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19824 0 -1 20384
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__icgtn_2  cm_inst.cc_inst.icgtn_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14448 0 1 29792
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__icgtn_4  cm_inst.cc_inst.icgtn_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14448 0 1 28224
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__icgtp_1  cm_inst.cc_inst.icgtp_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13664 0 -1 28224
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__icgtp_2  cm_inst.cc_inst.icgtp_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__icgtp_4  cm_inst.cc_inst.icgtp_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  cm_inst.cc_inst.inv_1_inst
timestamp 1698431365
transform -1 0 28000 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  cm_inst.cc_inst.inv_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26656 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_3  cm_inst.cc_inst.inv_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26656 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_4  cm_inst.cc_inst.inv_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  cm_inst.cc_inst.inv_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29120 0 1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_12  cm_inst.cc_inst.inv_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_16  cm_inst.cc_inst.inv_16_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27776 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__inv_20  cm_inst.cc_inst.inv_20_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14000 0 1 6272
box -86 -86 4790 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  cm_inst.cc_inst.invz_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 -1 42336
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  cm_inst.cc_inst.invz_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43344 0 -1 36064
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  cm_inst.cc_inst.invz_3_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42896 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_4  cm_inst.cc_inst.invz_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41776 0 1 34496
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__invz_8  cm_inst.cc_inst.invz_8_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12656 0 -1 42336
box -86 -86 4454 870
use gf180mcu_fd_sc_mcu7t5v0__invz_12  cm_inst.cc_inst.invz_12_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 6134 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  cm_inst.cc_inst.latq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28896 0 -1 20384
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_2  cm_inst.cc_inst.latq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30240 0 -1 15680
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latq_4  cm_inst.cc_inst.latq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37408 0 -1 29792
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  cm_inst.cc_inst.latrnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33712 0 -1 29792
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_2  cm_inst.cc_inst.latrnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31696 0 1 21952
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_4  cm_inst.cc_inst.latrnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__latrsnq_1  cm_inst.cc_inst.latrsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27664 0 -1 43904
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__latrsnq_2  cm_inst.cc_inst.latrsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__latrsnq_4  cm_inst.cc_inst.latrsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14672 0 1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__latsnq_1  cm_inst.cc_inst.latsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33264 0 -1 7840
box -86 -86 2438 870
use gf180mcu_fd_sc_mcu7t5v0__latsnq_2  cm_inst.cc_inst.latsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__latsnq_4  cm_inst.cc_inst.latsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39984 0 1 31360
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_1  cm_inst.cc_inst.mux2_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39088 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  cm_inst.cc_inst.mux2_2_inst
timestamp 1698431365
transform 1 0 34944 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_4  cm_inst.cc_inst.mux2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29232 0 -1 23520
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  cm_inst.cc_inst.mux4_1_inst
timestamp 1698431365
transform 1 0 33040 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_2  cm_inst.cc_inst.mux4_2_inst
timestamp 1698431365
transform 1 0 40656 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_4  cm_inst.cc_inst.mux4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39648 0 1 21952
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  cm_inst.cc_inst.nand2_1_inst
timestamp 1698431365
transform 1 0 24304 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  cm_inst.cc_inst.nand2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24976 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  cm_inst.cc_inst.nand2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20384 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  cm_inst.cc_inst.nand3_1_inst
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  cm_inst.cc_inst.nand3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26656 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  cm_inst.cc_inst.nand3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32704 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  cm_inst.cc_inst.nand4_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  cm_inst.cc_inst.nand4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23072 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  cm_inst.cc_inst.nand4_4_inst
timestamp 1698431365
transform 1 0 23184 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  cm_inst.cc_inst.nor2_1_inst
timestamp 1698431365
transform -1 0 26656 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  cm_inst.cc_inst.nor2_2_inst
timestamp 1698431365
transform -1 0 20608 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  cm_inst.cc_inst.nor2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22736 0 -1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  cm_inst.cc_inst.nor3_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  cm_inst.cc_inst.nor3_2_inst
timestamp 1698431365
transform 1 0 30800 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  cm_inst.cc_inst.nor3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14112 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  cm_inst.cc_inst.nor4_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22624 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  cm_inst.cc_inst.nor4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22848 0 -1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  cm_inst.cc_inst.nor4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23296 0 1 36064
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  cm_inst.cc_inst.oai21_1_inst
timestamp 1698431365
transform -1 0 24864 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  cm_inst.cc_inst.oai21_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38864 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  cm_inst.cc_inst.oai21_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32144 0 -1 10976
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  cm_inst.cc_inst.oai22_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34048 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  cm_inst.cc_inst.oai22_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26656 0 1 15680
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  cm_inst.cc_inst.oai22_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 36624 0 1 36064
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  cm_inst.cc_inst.oai31_1_inst
timestamp 1698431365
transform -1 0 34944 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  cm_inst.cc_inst.oai31_2_inst
timestamp 1698431365
transform 1 0 42224 0 1 28224
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  cm_inst.cc_inst.oai31_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23296 0 1 10976
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  cm_inst.cc_inst.oai32_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  cm_inst.cc_inst.oai32_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29120 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  cm_inst.cc_inst.oai32_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31248 0 1 10976
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_1  cm_inst.cc_inst.oai33_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26992 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_2  cm_inst.cc_inst.oai33_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34832 0 -1 37632
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_4  cm_inst.cc_inst.oai33_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33040 0 -1 18816
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  cm_inst.cc_inst.oai211_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  cm_inst.cc_inst.oai211_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44352 0 -1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  cm_inst.cc_inst.oai211_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42224 0 -1 21952
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  cm_inst.cc_inst.oai221_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33600 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  cm_inst.cc_inst.oai221_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 36176 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  cm_inst.cc_inst.oai221_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40880 0 -1 28224
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_1  cm_inst.cc_inst.oai222_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37072 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  cm_inst.cc_inst.oai222_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31696 0 1 21952
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_4  cm_inst.cc_inst.oai222_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33824 0 -1 23520
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  cm_inst.cc_inst.or2_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16576 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  cm_inst.cc_inst.or2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  cm_inst.cc_inst.or2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  cm_inst.cc_inst.or3_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  cm_inst.cc_inst.or3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13664 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_4  cm_inst.cc_inst.or3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18480 0 1 36064
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  cm_inst.cc_inst.or4_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  cm_inst.cc_inst.or4_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21504 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or4_4  cm_inst.cc_inst.or4_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12880 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__sdffq_1  cm_inst.cc_inst.sdffq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12432 0 -1 32928
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__sdffq_2  cm_inst.cc_inst.sdffq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41664 0 -1 12544
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__sdffq_4  cm_inst.cc_inst.sdffq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 5014 870
use gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1  cm_inst.cc_inst.sdffrnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41216 0 -1 18816
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2  cm_inst.cc_inst.sdffrnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 5126 870
use gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4  cm_inst.cc_inst.sdffrnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38304 0 1 14112
box -86 -86 5574 870
use gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1  cm_inst.cc_inst.sdffrsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 5462 870
use gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2  cm_inst.cc_inst.sdffrsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4  cm_inst.cc_inst.sdffrsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14896 0 1 39200
box -86 -86 6134 870
use gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1  cm_inst.cc_inst.sdffsnq_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37632 0 1 10976
box -86 -86 5126 870
use gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2  cm_inst.cc_inst.sdffsnq_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26992 0 -1 36064
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4  cm_inst.cc_inst.sdffsnq_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38528 0 1 18816
box -86 -86 6022 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  cm_inst.cc_inst.tieh_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 33376 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  cm_inst.cc_inst.tiel_inst
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  cm_inst.cc_inst.xnor2_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20608 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  cm_inst.cc_inst.xnor2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19040 0 1 6272
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_4  cm_inst.cc_inst.xnor2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28224 0 -1 29792
box -86 -86 2438 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  cm_inst.cc_inst.xnor3_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  cm_inst.cc_inst.xnor3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19152 0 -1 37632
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_4  cm_inst.cc_inst.xnor3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17696 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  cm_inst.cc_inst.xor2_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22736 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  cm_inst.cc_inst.xor2_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13888 0 1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  cm_inst.cc_inst.xor2_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19600 0 -1 31360
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  cm_inst.cc_inst.xor3_1_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19264 0 -1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  cm_inst.cc_inst.xor3_2_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43008 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_4  cm_inst.cc_inst.xor3_4_inst test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25424 0 -1 10976
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout17
timestamp 1698431365
transform -1 0 15680 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout18
timestamp 1698431365
transform -1 0 35840 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout19
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout20
timestamp 1698431365
transform 1 0 36512 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout21
timestamp 1698431365
transform -1 0 38640 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout22
timestamp 1698431365
transform 1 0 35504 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout23
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout24
timestamp 1698431365
transform 1 0 15680 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout25
timestamp 1698431365
transform 1 0 19152 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout26
timestamp 1698431365
transform -1 0 31920 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout27
timestamp 1698431365
transform 1 0 32032 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout28
timestamp 1698431365
transform -1 0 31920 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout29
timestamp 1698431365
transform -1 0 33824 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout30
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout31
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout32
timestamp 1698431365
transform -1 0 32592 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout33
timestamp 1698431365
transform 1 0 35728 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout34
timestamp 1698431365
transform 1 0 42560 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout35
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout36
timestamp 1698431365
transform -1 0 33488 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout37
timestamp 1698431365
transform -1 0 13104 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout38
timestamp 1698431365
transform 1 0 21840 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout39
timestamp 1698431365
transform -1 0 18480 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout40
timestamp 1698431365
transform 1 0 13664 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout41
timestamp 1698431365
transform -1 0 15232 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout42
timestamp 1698431365
transform 1 0 34608 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout43
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout44
timestamp 1698431365
transform -1 0 33600 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout45
timestamp 1698431365
transform -1 0 37744 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout46
timestamp 1698431365
transform -1 0 32704 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout47
timestamp 1698431365
transform -1 0 38640 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout48
timestamp 1698431365
transform 1 0 39424 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout49
timestamp 1698431365
transform -1 0 39312 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout50
timestamp 1698431365
transform 1 0 34720 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout51
timestamp 1698431365
transform 1 0 33040 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout52
timestamp 1698431365
transform 1 0 16128 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout53
timestamp 1698431365
transform -1 0 18144 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout54
timestamp 1698431365
transform -1 0 16464 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout55
timestamp 1698431365
transform -1 0 22736 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout56
timestamp 1698431365
transform 1 0 21952 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout57
timestamp 1698431365
transform -1 0 17024 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout58
timestamp 1698431365
transform -1 0 16352 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout59
timestamp 1698431365
transform 1 0 38528 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout60
timestamp 1698431365
transform 1 0 41776 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout61
timestamp 1698431365
transform 1 0 32144 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout62
timestamp 1698431365
transform 1 0 31024 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout63
timestamp 1698431365
transform -1 0 31024 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout64
timestamp 1698431365
transform -1 0 40544 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout65
timestamp 1698431365
transform -1 0 45360 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout66
timestamp 1698431365
transform 1 0 39312 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout67
timestamp 1698431365
transform 1 0 31920 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout68
timestamp 1698431365
transform 1 0 31360 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout69
timestamp 1698431365
transform 1 0 16352 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout70
timestamp 1698431365
transform 1 0 15456 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout71
timestamp 1698431365
transform 1 0 13216 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout72
timestamp 1698431365
transform 1 0 11088 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout73
timestamp 1698431365
transform 1 0 22736 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout74
timestamp 1698431365
transform 1 0 22848 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout75
timestamp 1698431365
transform 1 0 20272 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout76
timestamp 1698431365
transform -1 0 21840 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout77
timestamp 1698431365
transform -1 0 24640 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout78
timestamp 1698431365
transform 1 0 11872 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout79
timestamp 1698431365
transform 1 0 26656 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout80
timestamp 1698431365
transform 1 0 10752 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout81
timestamp 1698431365
transform -1 0 12432 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout82
timestamp 1698431365
transform -1 0 30688 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout83
timestamp 1698431365
transform -1 0 32256 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout84
timestamp 1698431365
transform 1 0 30912 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout85
timestamp 1698431365
transform -1 0 32592 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout86
timestamp 1698431365
transform 1 0 37408 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout87
timestamp 1698431365
transform 1 0 37632 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout88
timestamp 1698431365
transform 1 0 30688 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout89
timestamp 1698431365
transform 1 0 29232 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout90
timestamp 1698431365
transform 1 0 34944 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout91
timestamp 1698431365
transform -1 0 35616 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout92
timestamp 1698431365
transform -1 0 39648 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout93
timestamp 1698431365
transform -1 0 43904 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout94
timestamp 1698431365
transform -1 0 38640 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout95
timestamp 1698431365
transform -1 0 46256 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout96
timestamp 1698431365
transform 1 0 37520 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout97
timestamp 1698431365
transform 1 0 27440 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout98
timestamp 1698431365
transform 1 0 28560 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout99
timestamp 1698431365
transform -1 0 12096 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout100
timestamp 1698431365
transform -1 0 15232 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout101
timestamp 1698431365
transform 1 0 12992 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout102
timestamp 1698431365
transform -1 0 15680 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout103
timestamp 1698431365
transform -1 0 14448 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout104
timestamp 1698431365
transform 1 0 12768 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout105
timestamp 1698431365
transform -1 0 20048 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout106
timestamp 1698431365
transform -1 0 25984 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout107
timestamp 1698431365
transform 1 0 21728 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout108
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout109
timestamp 1698431365
transform -1 0 15232 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout110
timestamp 1698431365
transform -1 0 17920 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout111
timestamp 1698431365
transform 1 0 28224 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout112
timestamp 1698431365
transform 1 0 34272 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout113
timestamp 1698431365
transform 1 0 27440 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout114
timestamp 1698431365
transform -1 0 37856 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout115
timestamp 1698431365
transform -1 0 46032 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout116
timestamp 1698431365
transform 1 0 37632 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout117
timestamp 1698431365
transform 1 0 37856 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout118
timestamp 1698431365
transform -1 0 34272 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout119
timestamp 1698431365
transform -1 0 30800 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout120
timestamp 1698431365
transform -1 0 34944 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout121
timestamp 1698431365
transform -1 0 38752 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout122
timestamp 1698431365
transform -1 0 39648 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout123
timestamp 1698431365
transform 1 0 38416 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout124
timestamp 1698431365
transform 1 0 38416 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout125
timestamp 1698431365
transform 1 0 34160 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout126
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout127
timestamp 1698431365
transform 1 0 15904 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout128
timestamp 1698431365
transform -1 0 12768 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout129
timestamp 1698431365
transform -1 0 16016 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout130
timestamp 1698431365
transform 1 0 15344 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout131
timestamp 1698431365
transform 1 0 12432 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout132
timestamp 1698431365
transform -1 0 13104 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout133
timestamp 1698431365
transform -1 0 20048 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout134
timestamp 1698431365
transform -1 0 20832 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout135
timestamp 1698431365
transform -1 0 24864 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout136
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout137
timestamp 1698431365
transform 1 0 19488 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout138
timestamp 1698431365
transform -1 0 24416 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout139
timestamp 1698431365
transform 1 0 20608 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout140
timestamp 1698431365
transform 1 0 12432 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout141
timestamp 1698431365
transform -1 0 12768 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout142
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout143
timestamp 1698431365
transform -1 0 13216 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout144
timestamp 1698431365
transform -1 0 31136 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout145
timestamp 1698431365
transform 1 0 35616 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout146
timestamp 1698431365
transform 1 0 29904 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout147
timestamp 1698431365
transform -1 0 34720 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout148
timestamp 1698431365
transform 1 0 29344 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout149
timestamp 1698431365
transform -1 0 38528 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout150
timestamp 1698431365
transform 1 0 30016 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout151
timestamp 1698431365
transform -1 0 30800 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout152
timestamp 1698431365
transform -1 0 36848 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout153
timestamp 1698431365
transform 1 0 28224 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout154
timestamp 1698431365
transform -1 0 36512 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout155
timestamp 1698431365
transform -1 0 31472 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout156
timestamp 1698431365
transform -1 0 39648 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout157
timestamp 1698431365
transform -1 0 40544 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout158
timestamp 1698431365
transform -1 0 38528 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout159
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout160
timestamp 1698431365
transform 1 0 39536 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout161
timestamp 1698431365
transform 1 0 29904 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout162
timestamp 1698431365
transform 1 0 29120 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout163
timestamp 1698431365
transform -1 0 14448 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout164
timestamp 1698431365
transform -1 0 17024 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout165
timestamp 1698431365
transform -1 0 15904 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout166
timestamp 1698431365
transform -1 0 14448 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout167
timestamp 1698431365
transform 1 0 23968 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout168
timestamp 1698431365
transform 1 0 24976 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout169
timestamp 1698431365
transform -1 0 20944 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout170
timestamp 1698431365
transform 1 0 22064 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout171
timestamp 1698431365
transform -1 0 14784 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout172
timestamp 1698431365
transform -1 0 16016 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout173
timestamp 1698431365
transform 1 0 11648 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout174
timestamp 1698431365
transform 1 0 18480 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout175
timestamp 1698431365
transform -1 0 19376 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout176
timestamp 1698431365
transform -1 0 20944 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout177
timestamp 1698431365
transform -1 0 20272 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout178
timestamp 1698431365
transform 1 0 23632 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout179
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout180
timestamp 1698431365
transform 1 0 15568 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout181
timestamp 1698431365
transform -1 0 15232 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout182
timestamp 1698431365
transform 1 0 29680 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout183
timestamp 1698431365
transform -1 0 32480 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout184
timestamp 1698431365
transform 1 0 28112 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout185
timestamp 1698431365
transform 1 0 38752 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout186
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout187
timestamp 1698431365
transform 1 0 39312 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout188
timestamp 1698431365
transform -1 0 45360 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout189
timestamp 1698431365
transform -1 0 28112 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout190
timestamp 1698431365
transform -1 0 31136 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout191
timestamp 1698431365
transform 1 0 32032 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout192
timestamp 1698431365
transform -1 0 29904 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout193
timestamp 1698431365
transform -1 0 37744 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout194
timestamp 1698431365
transform 1 0 39648 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout195
timestamp 1698431365
transform 1 0 37520 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout196
timestamp 1698431365
transform -1 0 39984 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout197
timestamp 1698431365
transform -1 0 30576 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout198
timestamp 1698431365
transform -1 0 33600 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout199
timestamp 1698431365
transform 1 0 15232 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout200
timestamp 1698431365
transform 1 0 14672 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout201
timestamp 1698431365
transform 1 0 13216 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout202
timestamp 1698431365
transform 1 0 11760 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout203
timestamp 1698431365
transform -1 0 14672 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  fanout204
timestamp 1698431365
transform -1 0 17024 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout205
timestamp 1698431365
transform -1 0 19488 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout206
timestamp 1698431365
transform 1 0 18592 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout207
timestamp 1698431365
transform 1 0 24752 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout208
timestamp 1698431365
transform 1 0 23744 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout209
timestamp 1698431365
transform 1 0 20160 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout210
timestamp 1698431365
transform -1 0 19264 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout211
timestamp 1698431365
transform -1 0 21504 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout212
timestamp 1698431365
transform 1 0 22400 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout213
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout214
timestamp 1698431365
transform 1 0 22400 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout215
timestamp 1698431365
transform 1 0 19488 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout216
timestamp 1698431365
transform -1 0 20832 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout217
timestamp 1698431365
transform 1 0 14448 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  fanout218
timestamp 1698431365
transform -1 0 19488 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout219
timestamp 1698431365
transform -1 0 18256 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout220
timestamp 1698431365
transform -1 0 19824 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout221
timestamp 1698431365
transform 1 0 19040 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout222
timestamp 1698431365
transform 1 0 9520 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout223
timestamp 1698431365
transform 1 0 10192 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout224
timestamp 1698431365
transform -1 0 28784 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout225
timestamp 1698431365
transform -1 0 29680 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout226
timestamp 1698431365
transform -1 0 33824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout227
timestamp 1698431365
transform -1 0 30912 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout228
timestamp 1698431365
transform -1 0 30128 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout229
timestamp 1698431365
transform -1 0 37520 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout230
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout231
timestamp 1698431365
transform 1 0 27328 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout232
timestamp 1698431365
transform 1 0 27888 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout233
timestamp 1698431365
transform -1 0 29904 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout234
timestamp 1698431365
transform 1 0 28112 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout235
timestamp 1698431365
transform -1 0 36512 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout236
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout237
timestamp 1698431365
transform -1 0 37856 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout238
timestamp 1698431365
transform -1 0 39424 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout239
timestamp 1698431365
transform 1 0 38416 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout240
timestamp 1698431365
transform -1 0 43008 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout241
timestamp 1698431365
transform -1 0 37968 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout242
timestamp 1698431365
transform 1 0 40992 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout243
timestamp 1698431365
transform 1 0 38080 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout244
timestamp 1698431365
transform 1 0 29232 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout245
timestamp 1698431365
transform -1 0 30128 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout246
timestamp 1698431365
transform -1 0 12096 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout247
timestamp 1698431365
transform -1 0 13104 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout248
timestamp 1698431365
transform -1 0 12992 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout249
timestamp 1698431365
transform -1 0 14224 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout250
timestamp 1698431365
transform -1 0 24864 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout251
timestamp 1698431365
transform -1 0 26208 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout252
timestamp 1698431365
transform 1 0 24080 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout253
timestamp 1698431365
transform 1 0 19824 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout254
timestamp 1698431365
transform 1 0 20720 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout255
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout256
timestamp 1698431365
transform 1 0 12432 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout257
timestamp 1698431365
transform -1 0 14000 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout258
timestamp 1698431365
transform 1 0 9184 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout259
timestamp 1698431365
transform 1 0 10976 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout260
timestamp 1698431365
transform -1 0 24752 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout261
timestamp 1698431365
transform 1 0 24752 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout262
timestamp 1698431365
transform -1 0 20160 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout263
timestamp 1698431365
transform -1 0 20944 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout264
timestamp 1698431365
transform 1 0 22736 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout265
timestamp 1698431365
transform 1 0 20832 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout266
timestamp 1698431365
transform -1 0 11648 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout267
timestamp 1698431365
transform 1 0 11424 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  fanout268
timestamp 1698431365
transform 1 0 29120 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout269
timestamp 1698431365
transform 1 0 28336 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout270
timestamp 1698431365
transform 1 0 27552 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  fanout271
timestamp 1698431365
transform -1 0 28784 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout272
timestamp 1698431365
transform -1 0 30800 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout273
timestamp 1698431365
transform 1 0 33040 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout274
timestamp 1698431365
transform -1 0 28784 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout275
timestamp 1698431365
transform 1 0 34496 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout276
timestamp 1698431365
transform 1 0 43680 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout277
timestamp 1698431365
transform 1 0 45360 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout278
timestamp 1698431365
transform 1 0 37184 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout279
timestamp 1698431365
transform 1 0 38528 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout280
timestamp 1698431365
transform -1 0 29680 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout281
timestamp 1698431365
transform -1 0 28448 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout282
timestamp 1698431365
transform 1 0 27776 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout283
timestamp 1698431365
transform -1 0 28784 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout284
timestamp 1698431365
transform -1 0 28672 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout285
timestamp 1698431365
transform 1 0 40768 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout286
timestamp 1698431365
transform -1 0 41216 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout287
timestamp 1698431365
transform -1 0 39648 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout288
timestamp 1698431365
transform -1 0 41664 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout289
timestamp 1698431365
transform 1 0 39984 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout290
timestamp 1698431365
transform -1 0 28896 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout291
timestamp 1698431365
transform -1 0 32704 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout292
timestamp 1698431365
transform 1 0 11760 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout293
timestamp 1698431365
transform 1 0 9744 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout294
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout295
timestamp 1698431365
transform -1 0 5152 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout296
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout297
timestamp 1698431365
transform 1 0 7840 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout298
timestamp 1698431365
transform 1 0 4144 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout299
timestamp 1698431365
transform -1 0 6384 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout300
timestamp 1698431365
transform -1 0 5264 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout301
timestamp 1698431365
transform -1 0 7168 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout302
timestamp 1698431365
transform -1 0 6496 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout303
timestamp 1698431365
transform 1 0 12992 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout304
timestamp 1698431365
transform -1 0 8064 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout305
timestamp 1698431365
transform -1 0 7168 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout306
timestamp 1698431365
transform -1 0 5152 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout307
timestamp 1698431365
transform -1 0 6160 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout308
timestamp 1698431365
transform -1 0 6384 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout309
timestamp 1698431365
transform -1 0 5264 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout310
timestamp 1698431365
transform 1 0 3920 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout311
timestamp 1698431365
transform -1 0 10864 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout312
timestamp 1698431365
transform 1 0 3248 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout313
timestamp 1698431365
transform -1 0 6160 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout314
timestamp 1698431365
transform 1 0 6160 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_138 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_154 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18592 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_158 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_160 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19264 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_167
timestamp 1698431365
transform 1 0 20048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698431365
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_392 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45248 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_400
timestamp 1698431365
transform 1 0 46144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_186
timestamp 1698431365
transform 1 0 22176 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_190
timestamp 1698431365
transform 1 0 22624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_384
timestamp 1698431365
transform 1 0 44352 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_400
timestamp 1698431365
transform 1 0 46144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_6
timestamp 1698431365
transform 1 0 2016 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_22
timestamp 1698431365
transform 1 0 3808 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_30
timestamp 1698431365
transform 1 0 4704 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_227
timestamp 1698431365
transform 1 0 26768 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_395
timestamp 1698431365
transform 1 0 45584 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_399
timestamp 1698431365
transform 1 0 46032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_401
timestamp 1698431365
transform 1 0 46256 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_6
timestamp 1698431365
transform 1 0 2016 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_41
timestamp 1698431365
transform 1 0 5936 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_57
timestamp 1698431365
transform 1 0 7728 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_65
timestamp 1698431365
transform 1 0 8624 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_69
timestamp 1698431365
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_104
timestamp 1698431365
transform 1 0 12992 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_120
timestamp 1698431365
transform 1 0 14784 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_124
timestamp 1698431365
transform 1 0 15232 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_126
timestamp 1698431365
transform 1 0 15456 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_220
timestamp 1698431365
transform 1 0 25984 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_224
timestamp 1698431365
transform 1 0 26432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_263
timestamp 1698431365
transform 1 0 30800 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_384
timestamp 1698431365
transform 1 0 44352 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_400
timestamp 1698431365
transform 1 0 46144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_111
timestamp 1698431365
transform 1 0 13776 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_155
timestamp 1698431365
transform 1 0 18704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_157
timestamp 1698431365
transform 1 0 18928 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_217
timestamp 1698431365
transform 1 0 25648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_253
timestamp 1698431365
transform 1 0 29680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_291
timestamp 1698431365
transform 1 0 33936 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_307
timestamp 1698431365
transform 1 0 35728 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_395
timestamp 1698431365
transform 1 0 45584 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_399
timestamp 1698431365
transform 1 0 46032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_401
timestamp 1698431365
transform 1 0 46256 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_38
timestamp 1698431365
transform 1 0 5600 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_150
timestamp 1698431365
transform 1 0 18144 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_199
timestamp 1698431365
transform 1 0 23632 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_201
timestamp 1698431365
transform 1 0 23856 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_284
timestamp 1698431365
transform 1 0 33152 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_384
timestamp 1698431365
transform 1 0 44352 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_400
timestamp 1698431365
transform 1 0 46144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_131
timestamp 1698431365
transform 1 0 16016 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_147
timestamp 1698431365
transform 1 0 17808 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_151
timestamp 1698431365
transform 1 0 18256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_153
timestamp 1698431365
transform 1 0 18480 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_183
timestamp 1698431365
transform 1 0 21840 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_199
timestamp 1698431365
transform 1 0 23632 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_239
timestamp 1698431365
transform 1 0 28112 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_243
timestamp 1698431365
transform 1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_259
timestamp 1698431365
transform 1 0 30352 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_312
timestamp 1698431365
transform 1 0 36288 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_314
timestamp 1698431365
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_321
timestamp 1698431365
transform 1 0 37296 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_323
timestamp 1698431365
transform 1 0 37520 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_357
timestamp 1698431365
transform 1 0 41328 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_373
timestamp 1698431365
transform 1 0 43120 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698431365
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_395
timestamp 1698431365
transform 1 0 45584 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_399
timestamp 1698431365
transform 1 0 46032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_401
timestamp 1698431365
transform 1 0 46256 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_10
timestamp 1698431365
transform 1 0 2464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_48
timestamp 1698431365
transform 1 0 6720 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_64
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_68
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_74
timestamp 1698431365
transform 1 0 9632 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_79
timestamp 1698431365
transform 1 0 10192 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_95
timestamp 1698431365
transform 1 0 11984 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_129
timestamp 1698431365
transform 1 0 15792 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_137
timestamp 1698431365
transform 1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_146
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_148
timestamp 1698431365
transform 1 0 17920 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_174
timestamp 1698431365
transform 1 0 20832 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_190
timestamp 1698431365
transform 1 0 22624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_226
timestamp 1698431365
transform 1 0 26656 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_242
timestamp 1698431365
transform 1 0 28448 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_250
timestamp 1698431365
transform 1 0 29344 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_257
timestamp 1698431365
transform 1 0 30128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_261
timestamp 1698431365
transform 1 0 30576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_288
timestamp 1698431365
transform 1 0 33600 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_296
timestamp 1698431365
transform 1 0 34496 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_333
timestamp 1698431365
transform 1 0 38640 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_349
timestamp 1698431365
transform 1 0 40432 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_383
timestamp 1698431365
transform 1 0 44240 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_399
timestamp 1698431365
transform 1 0 46032 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_401
timestamp 1698431365
transform 1 0 46256 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_18
timestamp 1698431365
transform 1 0 3360 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_22
timestamp 1698431365
transform 1 0 3808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_28
timestamp 1698431365
transform 1 0 4480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_39
timestamp 1698431365
transform 1 0 5712 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_44
timestamp 1698431365
transform 1 0 6272 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_52
timestamp 1698431365
transform 1 0 7168 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_56
timestamp 1698431365
transform 1 0 7616 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_91
timestamp 1698431365
transform 1 0 11536 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_109
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_170
timestamp 1698431365
transform 1 0 20384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_191
timestamp 1698431365
transform 1 0 22736 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_233
timestamp 1698431365
transform 1 0 27440 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_249
timestamp 1698431365
transform 1 0 29232 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_276
timestamp 1698431365
transform 1 0 32256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_278
timestamp 1698431365
transform 1 0 32480 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_313
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_329
timestamp 1698431365
transform 1 0 38192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_362
timestamp 1698431365
transform 1 0 41888 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_378
timestamp 1698431365
transform 1 0 43680 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_382
timestamp 1698431365
transform 1 0 44128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1698431365
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_395
timestamp 1698431365
transform 1 0 45584 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_399
timestamp 1698431365
transform 1 0 46032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_401
timestamp 1698431365
transform 1 0 46256 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_184
timestamp 1698431365
transform 1 0 21952 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_186
timestamp 1698431365
transform 1 0 22176 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_214
timestamp 1698431365
transform 1 0 25312 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_275
timestamp 1698431365
transform 1 0 32144 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_292
timestamp 1698431365
transform 1 0 34048 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_324
timestamp 1698431365
transform 1 0 37632 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_340
timestamp 1698431365
transform 1 0 39424 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_348
timestamp 1698431365
transform 1 0 40320 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_384
timestamp 1698431365
transform 1 0 44352 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_400
timestamp 1698431365
transform 1 0 46144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_18
timestamp 1698431365
transform 1 0 3360 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_27
timestamp 1698431365
transform 1 0 4368 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_45
timestamp 1698431365
transform 1 0 6384 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_111
timestamp 1698431365
transform 1 0 13776 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_172
timestamp 1698431365
transform 1 0 20608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_187
timestamp 1698431365
transform 1 0 22288 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_239
timestamp 1698431365
transform 1 0 28112 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_243
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_263
timestamp 1698431365
transform 1 0 30800 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_310
timestamp 1698431365
transform 1 0 36064 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_314
timestamp 1698431365
transform 1 0 36512 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_323
timestamp 1698431365
transform 1 0 37520 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_369
timestamp 1698431365
transform 1 0 42672 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_395
timestamp 1698431365
transform 1 0 45584 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_399
timestamp 1698431365
transform 1 0 46032 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_401
timestamp 1698431365
transform 1 0 46256 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_80
timestamp 1698431365
transform 1 0 10304 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_88
timestamp 1698431365
transform 1 0 11200 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_144
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_154
timestamp 1698431365
transform 1 0 18592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_156
timestamp 1698431365
transform 1 0 18816 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_178
timestamp 1698431365
transform 1 0 21280 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_182
timestamp 1698431365
transform 1 0 21728 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_244
timestamp 1698431365
transform 1 0 28672 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_318
timestamp 1698431365
transform 1 0 36960 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_356
timestamp 1698431365
transform 1 0 41216 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_400
timestamp 1698431365
transform 1 0 46144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_22
timestamp 1698431365
transform 1 0 3808 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_30
timestamp 1698431365
transform 1 0 4704 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_53
timestamp 1698431365
transform 1 0 7280 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_61
timestamp 1698431365
transform 1 0 8176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_67
timestamp 1698431365
transform 1 0 8848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_131
timestamp 1698431365
transform 1 0 16016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_135
timestamp 1698431365
transform 1 0 16464 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_168
timestamp 1698431365
transform 1 0 20160 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_172
timestamp 1698431365
transform 1 0 20608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_193
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_203
timestamp 1698431365
transform 1 0 24080 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_210
timestamp 1698431365
transform 1 0 24864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_218
timestamp 1698431365
transform 1 0 25760 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_222
timestamp 1698431365
transform 1 0 26208 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_240
timestamp 1698431365
transform 1 0 28224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_282
timestamp 1698431365
transform 1 0 32928 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_319
timestamp 1698431365
transform 1 0 37072 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_330
timestamp 1698431365
transform 1 0 38304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_375
timestamp 1698431365
transform 1 0 43344 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_383
timestamp 1698431365
transform 1 0 44240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_395
timestamp 1698431365
transform 1 0 45584 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_399
timestamp 1698431365
transform 1 0 46032 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_401
timestamp 1698431365
transform 1 0 46256 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_76
timestamp 1698431365
transform 1 0 9856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_78
timestamp 1698431365
transform 1 0 10080 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_108
timestamp 1698431365
transform 1 0 13440 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_112
timestamp 1698431365
transform 1 0 13888 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_131
timestamp 1698431365
transform 1 0 16016 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_144
timestamp 1698431365
transform 1 0 17472 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_153
timestamp 1698431365
transform 1 0 18480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_157
timestamp 1698431365
transform 1 0 18928 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_196
timestamp 1698431365
transform 1 0 23296 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_200
timestamp 1698431365
transform 1 0 23744 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_202
timestamp 1698431365
transform 1 0 23968 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_205
timestamp 1698431365
transform 1 0 24304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_228
timestamp 1698431365
transform 1 0 26880 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_244
timestamp 1698431365
transform 1 0 28672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_262
timestamp 1698431365
transform 1 0 30688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_264
timestamp 1698431365
transform 1 0 30912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_298
timestamp 1698431365
transform 1 0 34720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_347
timestamp 1698431365
transform 1 0 40208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_358
timestamp 1698431365
transform 1 0 41440 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_366
timestamp 1698431365
transform 1 0 42336 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_26
timestamp 1698431365
transform 1 0 4256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_45
timestamp 1698431365
transform 1 0 6384 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_49
timestamp 1698431365
transform 1 0 6832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_55
timestamp 1698431365
transform 1 0 7504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_57
timestamp 1698431365
transform 1 0 7728 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_64
timestamp 1698431365
transform 1 0 8512 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_72
timestamp 1698431365
transform 1 0 9408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_103
timestamp 1698431365
transform 1 0 12880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_140
timestamp 1698431365
transform 1 0 17024 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_148
timestamp 1698431365
transform 1 0 17920 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_183
timestamp 1698431365
transform 1 0 21840 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_201
timestamp 1698431365
transform 1 0 23856 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_205
timestamp 1698431365
transform 1 0 24304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_209
timestamp 1698431365
transform 1 0 24752 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_268
timestamp 1698431365
transform 1 0 31360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_270
timestamp 1698431365
transform 1 0 31584 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_287
timestamp 1698431365
transform 1 0 33488 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_303
timestamp 1698431365
transform 1 0 35280 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_307
timestamp 1698431365
transform 1 0 35728 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_323
timestamp 1698431365
transform 1 0 37520 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_379
timestamp 1698431365
transform 1 0 43792 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_383
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_395
timestamp 1698431365
transform 1 0 45584 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_399
timestamp 1698431365
transform 1 0 46032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_401
timestamp 1698431365
transform 1 0 46256 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_22
timestamp 1698431365
transform 1 0 3808 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_24
timestamp 1698431365
transform 1 0 4032 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_65
timestamp 1698431365
transform 1 0 8624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_67
timestamp 1698431365
transform 1 0 8848 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_108
timestamp 1698431365
transform 1 0 13440 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_110
timestamp 1698431365
transform 1 0 13664 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_117
timestamp 1698431365
transform 1 0 14448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_133
timestamp 1698431365
transform 1 0 16240 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_192
timestamp 1698431365
transform 1 0 22848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_194
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_201
timestamp 1698431365
transform 1 0 23856 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_311
timestamp 1698431365
transform 1 0 36176 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_319
timestamp 1698431365
transform 1 0 37072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_6
timestamp 1698431365
transform 1 0 2016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_10
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_14
timestamp 1698431365
transform 1 0 2912 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_22
timestamp 1698431365
transform 1 0 3808 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_30
timestamp 1698431365
transform 1 0 4704 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_39
timestamp 1698431365
transform 1 0 5712 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_44
timestamp 1698431365
transform 1 0 6272 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_122
timestamp 1698431365
transform 1 0 15008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_126
timestamp 1698431365
transform 1 0 15456 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698431365
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_203
timestamp 1698431365
transform 1 0 24080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_234
timestamp 1698431365
transform 1 0 27552 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_236
timestamp 1698431365
transform 1 0 27776 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_269
timestamp 1698431365
transform 1 0 31472 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_310
timestamp 1698431365
transform 1 0 36064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_325
timestamp 1698431365
transform 1 0 37744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_327
timestamp 1698431365
transform 1 0 37968 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_380
timestamp 1698431365
transform 1 0 43904 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_384
timestamp 1698431365
transform 1 0 44352 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_395
timestamp 1698431365
transform 1 0 45584 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_399
timestamp 1698431365
transform 1 0 46032 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_401
timestamp 1698431365
transform 1 0 46256 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_106
timestamp 1698431365
transform 1 0 13216 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698431365
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698431365
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_204
timestamp 1698431365
transform 1 0 24192 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_229
timestamp 1698431365
transform 1 0 26992 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_273
timestamp 1698431365
transform 1 0 31920 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_317
timestamp 1698431365
transform 1 0 36848 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_321
timestamp 1698431365
transform 1 0 37296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_325
timestamp 1698431365
transform 1 0 37744 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_329
timestamp 1698431365
transform 1 0 38192 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_337
timestamp 1698431365
transform 1 0 39088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_347
timestamp 1698431365
transform 1 0 40208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_368
timestamp 1698431365
transform 1 0 42560 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_372
timestamp 1698431365
transform 1 0 43008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_374
timestamp 1698431365
transform 1 0 43232 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_397
timestamp 1698431365
transform 1 0 45808 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_401
timestamp 1698431365
transform 1 0 46256 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_14
timestamp 1698431365
transform 1 0 2912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_22
timestamp 1698431365
transform 1 0 3808 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_27
timestamp 1698431365
transform 1 0 4368 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_71
timestamp 1698431365
transform 1 0 9296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_96
timestamp 1698431365
transform 1 0 12096 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_141
timestamp 1698431365
transform 1 0 17136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_145
timestamp 1698431365
transform 1 0 17584 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_147
timestamp 1698431365
transform 1 0 17808 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_150
timestamp 1698431365
transform 1 0 18144 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_228
timestamp 1698431365
transform 1 0 26880 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_236
timestamp 1698431365
transform 1 0 27776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_238
timestamp 1698431365
transform 1 0 28000 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_257
timestamp 1698431365
transform 1 0 30128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_261
timestamp 1698431365
transform 1 0 30576 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_306
timestamp 1698431365
transform 1 0 35616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_310
timestamp 1698431365
transform 1 0 36064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_312
timestamp 1698431365
transform 1 0 36288 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_333
timestamp 1698431365
transform 1 0 38640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_371
timestamp 1698431365
transform 1 0 42896 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_379
timestamp 1698431365
transform 1 0 43792 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_383
timestamp 1698431365
transform 1 0 44240 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_395
timestamp 1698431365
transform 1 0 45584 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_399
timestamp 1698431365
transform 1 0 46032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_401
timestamp 1698431365
transform 1 0 46256 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_10
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_46
timestamp 1698431365
transform 1 0 6496 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_54
timestamp 1698431365
transform 1 0 7392 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_109
timestamp 1698431365
transform 1 0 13552 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_111
timestamp 1698431365
transform 1 0 13776 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_136
timestamp 1698431365
transform 1 0 16576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_155
timestamp 1698431365
transform 1 0 18704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_157
timestamp 1698431365
transform 1 0 18928 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_166
timestamp 1698431365
transform 1 0 19936 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_168
timestamp 1698431365
transform 1 0 20160 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_187
timestamp 1698431365
transform 1 0 22288 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_191
timestamp 1698431365
transform 1 0 22736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_216
timestamp 1698431365
transform 1 0 25536 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_248
timestamp 1698431365
transform 1 0 29120 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_261
timestamp 1698431365
transform 1 0 30576 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_269
timestamp 1698431365
transform 1 0 31472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_342
timestamp 1698431365
transform 1 0 39648 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_399
timestamp 1698431365
transform 1 0 46032 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_401
timestamp 1698431365
transform 1 0 46256 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_24
timestamp 1698431365
transform 1 0 4032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_26
timestamp 1698431365
transform 1 0 4256 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_45
timestamp 1698431365
transform 1 0 6384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_49
timestamp 1698431365
transform 1 0 6832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_95
timestamp 1698431365
transform 1 0 11984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_169
timestamp 1698431365
transform 1 0 20272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_179
timestamp 1698431365
transform 1 0 21392 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_184
timestamp 1698431365
transform 1 0 21952 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_235
timestamp 1698431365
transform 1 0 27664 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698431365
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_255
timestamp 1698431365
transform 1 0 29904 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_271
timestamp 1698431365
transform 1 0 31696 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_273
timestamp 1698431365
transform 1 0 31920 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_331
timestamp 1698431365
transform 1 0 38416 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_395
timestamp 1698431365
transform 1 0 45584 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_399
timestamp 1698431365
transform 1 0 46032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_401
timestamp 1698431365
transform 1 0 46256 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_8
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_43
timestamp 1698431365
transform 1 0 6160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_47
timestamp 1698431365
transform 1 0 6608 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_78
timestamp 1698431365
transform 1 0 10080 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_100
timestamp 1698431365
transform 1 0 12544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_104
timestamp 1698431365
transform 1 0 12992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_106
timestamp 1698431365
transform 1 0 13216 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_156
timestamp 1698431365
transform 1 0 18816 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_160
timestamp 1698431365
transform 1 0 19264 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_162
timestamp 1698431365
transform 1 0 19488 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_196
timestamp 1698431365
transform 1 0 23296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_198
timestamp 1698431365
transform 1 0 23520 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_228
timestamp 1698431365
transform 1 0 26880 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_236
timestamp 1698431365
transform 1 0 27776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_266
timestamp 1698431365
transform 1 0 31136 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698431365
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_392
timestamp 1698431365
transform 1 0 45248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_400
timestamp 1698431365
transform 1 0 46144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_28
timestamp 1698431365
transform 1 0 4480 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_39
timestamp 1698431365
transform 1 0 5712 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_52
timestamp 1698431365
transform 1 0 7168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_54
timestamp 1698431365
transform 1 0 7392 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_148
timestamp 1698431365
transform 1 0 17920 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_164
timestamp 1698431365
transform 1 0 19712 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_166
timestamp 1698431365
transform 1 0 19936 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_185
timestamp 1698431365
transform 1 0 22064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_187
timestamp 1698431365
transform 1 0 22288 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_203
timestamp 1698431365
transform 1 0 24080 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_207
timestamp 1698431365
transform 1 0 24528 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_223
timestamp 1698431365
transform 1 0 26320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_227
timestamp 1698431365
transform 1 0 26768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_372
timestamp 1698431365
transform 1 0 43008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_380
timestamp 1698431365
transform 1 0 43904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1698431365
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_395
timestamp 1698431365
transform 1 0 45584 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_399
timestamp 1698431365
transform 1 0 46032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_401
timestamp 1698431365
transform 1 0 46256 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_4
timestamp 1698431365
transform 1 0 1792 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_39
timestamp 1698431365
transform 1 0 5712 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_41
timestamp 1698431365
transform 1 0 5936 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_57
timestamp 1698431365
transform 1 0 7728 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_61
timestamp 1698431365
transform 1 0 8176 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_80
timestamp 1698431365
transform 1 0 10304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_102
timestamp 1698431365
transform 1 0 12768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_147
timestamp 1698431365
transform 1 0 17808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_151
timestamp 1698431365
transform 1 0 18256 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_159
timestamp 1698431365
transform 1 0 19152 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_176
timestamp 1698431365
transform 1 0 21056 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_180
timestamp 1698431365
transform 1 0 21504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_216
timestamp 1698431365
transform 1 0 25536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_218
timestamp 1698431365
transform 1 0 25760 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_233
timestamp 1698431365
transform 1 0 27440 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_246
timestamp 1698431365
transform 1 0 28896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_314
timestamp 1698431365
transform 1 0 36512 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_318
timestamp 1698431365
transform 1 0 36960 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698431365
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_329
timestamp 1698431365
transform 1 0 38192 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_345
timestamp 1698431365
transform 1 0 39984 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_360
timestamp 1698431365
transform 1 0 41664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_364
timestamp 1698431365
transform 1 0 42112 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_398
timestamp 1698431365
transform 1 0 45920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_28
timestamp 1698431365
transform 1 0 4480 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_66
timestamp 1698431365
transform 1 0 8736 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_70
timestamp 1698431365
transform 1 0 9184 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_86
timestamp 1698431365
transform 1 0 10976 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_90
timestamp 1698431365
transform 1 0 11424 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_99
timestamp 1698431365
transform 1 0 12432 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_113
timestamp 1698431365
transform 1 0 14000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_115
timestamp 1698431365
transform 1 0 14224 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_162
timestamp 1698431365
transform 1 0 19488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_164
timestamp 1698431365
transform 1 0 19712 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698431365
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_208
timestamp 1698431365
transform 1 0 24640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_216
timestamp 1698431365
transform 1 0 25536 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_223
timestamp 1698431365
transform 1 0 26320 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_304
timestamp 1698431365
transform 1 0 35392 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_308
timestamp 1698431365
transform 1 0 35840 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698431365
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_332
timestamp 1698431365
transform 1 0 38528 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_340
timestamp 1698431365
transform 1 0 39424 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_380
timestamp 1698431365
transform 1 0 43904 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_384
timestamp 1698431365
transform 1 0 44352 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_395
timestamp 1698431365
transform 1 0 45584 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_399
timestamp 1698431365
transform 1 0 46032 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_401
timestamp 1698431365
transform 1 0 46256 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_53
timestamp 1698431365
transform 1 0 7280 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_105
timestamp 1698431365
transform 1 0 13104 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_115
timestamp 1698431365
transform 1 0 14224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_124
timestamp 1698431365
transform 1 0 15232 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698431365
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_171
timestamp 1698431365
transform 1 0 20496 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_235
timestamp 1698431365
transform 1 0 27664 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_239
timestamp 1698431365
transform 1 0 28112 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_274
timestamp 1698431365
transform 1 0 32032 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_341
timestamp 1698431365
transform 1 0 39536 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_349
timestamp 1698431365
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_360
timestamp 1698431365
transform 1 0 41664 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_362
timestamp 1698431365
transform 1 0 41888 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_396
timestamp 1698431365
transform 1 0 45696 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_400
timestamp 1698431365
transform 1 0 46144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_28
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_67
timestamp 1698431365
transform 1 0 8848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_71
timestamp 1698431365
transform 1 0 9296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_111
timestamp 1698431365
transform 1 0 13776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_121
timestamp 1698431365
transform 1 0 14896 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_156
timestamp 1698431365
transform 1 0 18816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_202
timestamp 1698431365
transform 1 0 23968 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_238
timestamp 1698431365
transform 1 0 28000 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698431365
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_262
timestamp 1698431365
transform 1 0 30688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_266
timestamp 1698431365
transform 1 0 31136 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_281
timestamp 1698431365
transform 1 0 32816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_327
timestamp 1698431365
transform 1 0 37968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_401
timestamp 1698431365
transform 1 0 46256 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_41
timestamp 1698431365
transform 1 0 5936 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_80
timestamp 1698431365
transform 1 0 10304 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_109
timestamp 1698431365
transform 1 0 13552 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_125
timestamp 1698431365
transform 1 0 15344 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_133
timestamp 1698431365
transform 1 0 16240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_135
timestamp 1698431365
transform 1 0 16464 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_144
timestamp 1698431365
transform 1 0 17472 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_235
timestamp 1698431365
transform 1 0 27664 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_286
timestamp 1698431365
transform 1 0 33376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_290
timestamp 1698431365
transform 1 0 33824 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_332
timestamp 1698431365
transform 1 0 38528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_334
timestamp 1698431365
transform 1 0 38752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_109
timestamp 1698431365
transform 1 0 13552 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_141
timestamp 1698431365
transform 1 0 17136 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_143
timestamp 1698431365
transform 1 0 17360 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698431365
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_297
timestamp 1698431365
transform 1 0 34608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_301
timestamp 1698431365
transform 1 0 35056 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_309
timestamp 1698431365
transform 1 0 35952 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_339
timestamp 1698431365
transform 1 0 39312 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_343
timestamp 1698431365
transform 1 0 39760 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_345
timestamp 1698431365
transform 1 0 39984 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_380
timestamp 1698431365
transform 1 0 43904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_395
timestamp 1698431365
transform 1 0 45584 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_399
timestamp 1698431365
transform 1 0 46032 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_401
timestamp 1698431365
transform 1 0 46256 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_52
timestamp 1698431365
transform 1 0 7168 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_95
timestamp 1698431365
transform 1 0 11984 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_127
timestamp 1698431365
transform 1 0 15568 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_135
timestamp 1698431365
transform 1 0 16464 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698431365
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_229
timestamp 1698431365
transform 1 0 26992 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_231
timestamp 1698431365
transform 1 0 27216 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_294
timestamp 1698431365
transform 1 0 34272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_296
timestamp 1698431365
transform 1 0 34496 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_305
timestamp 1698431365
transform 1 0 35504 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_309
timestamp 1698431365
transform 1 0 35952 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_311
timestamp 1698431365
transform 1 0 36176 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_322
timestamp 1698431365
transform 1 0 37408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_340
timestamp 1698431365
transform 1 0 39424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_344
timestamp 1698431365
transform 1 0 39872 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_368
timestamp 1698431365
transform 1 0 42560 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_376
timestamp 1698431365
transform 1 0 43456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_384
timestamp 1698431365
transform 1 0 44352 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_400
timestamp 1698431365
transform 1 0 46144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698431365
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_53
timestamp 1698431365
transform 1 0 7280 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_94
timestamp 1698431365
transform 1 0 11872 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_102
timestamp 1698431365
transform 1 0 12768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_109
timestamp 1698431365
transform 1 0 13552 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_112
timestamp 1698431365
transform 1 0 13888 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_128
timestamp 1698431365
transform 1 0 15680 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_200
timestamp 1698431365
transform 1 0 23744 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_226
timestamp 1698431365
transform 1 0 26656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_230
timestamp 1698431365
transform 1 0 27104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_232
timestamp 1698431365
transform 1 0 27328 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_374
timestamp 1698431365
transform 1 0 43232 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_382
timestamp 1698431365
transform 1 0 44128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_384
timestamp 1698431365
transform 1 0 44352 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_395
timestamp 1698431365
transform 1 0 45584 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_399
timestamp 1698431365
transform 1 0 46032 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_401
timestamp 1698431365
transform 1 0 46256 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_36
timestamp 1698431365
transform 1 0 5376 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_44
timestamp 1698431365
transform 1 0 6272 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_84
timestamp 1698431365
transform 1 0 10752 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_100
timestamp 1698431365
transform 1 0 12544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698431365
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_163
timestamp 1698431365
transform 1 0 19600 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_187
timestamp 1698431365
transform 1 0 22288 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_189
timestamp 1698431365
transform 1 0 22512 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_217
timestamp 1698431365
transform 1 0 25648 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_224
timestamp 1698431365
transform 1 0 26432 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_233
timestamp 1698431365
transform 1 0 27440 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_247
timestamp 1698431365
transform 1 0 29008 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_288
timestamp 1698431365
transform 1 0 33600 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_292
timestamp 1698431365
transform 1 0 34048 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_334
timestamp 1698431365
transform 1 0 38752 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_336
timestamp 1698431365
transform 1 0 38976 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_396
timestamp 1698431365
transform 1 0 45696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_400
timestamp 1698431365
transform 1 0 46144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_41
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_80
timestamp 1698431365
transform 1 0 10304 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_88
timestamp 1698431365
transform 1 0 11200 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_169
timestamp 1698431365
transform 1 0 20272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_173
timestamp 1698431365
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_182
timestamp 1698431365
transform 1 0 21728 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_188
timestamp 1698431365
transform 1 0 22400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_192
timestamp 1698431365
transform 1 0 22848 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_216
timestamp 1698431365
transform 1 0 25536 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_232
timestamp 1698431365
transform 1 0 27328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_234
timestamp 1698431365
transform 1 0 27552 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_306
timestamp 1698431365
transform 1 0 35616 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_319
timestamp 1698431365
transform 1 0 37072 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_364
timestamp 1698431365
transform 1 0 42112 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_384
timestamp 1698431365
transform 1 0 44352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_397
timestamp 1698431365
transform 1 0 45808 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_401
timestamp 1698431365
transform 1 0 46256 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_43
timestamp 1698431365
transform 1 0 6160 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_59
timestamp 1698431365
transform 1 0 7952 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_67
timestamp 1698431365
transform 1 0 8848 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_69
timestamp 1698431365
transform 1 0 9072 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_148
timestamp 1698431365
transform 1 0 17920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_179
timestamp 1698431365
transform 1 0 21392 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_183
timestamp 1698431365
transform 1 0 21840 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_186
timestamp 1698431365
transform 1 0 22176 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_190
timestamp 1698431365
transform 1 0 22624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_192
timestamp 1698431365
transform 1 0 22848 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_201
timestamp 1698431365
transform 1 0 23856 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_224
timestamp 1698431365
transform 1 0 26432 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_238
timestamp 1698431365
transform 1 0 28000 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_261
timestamp 1698431365
transform 1 0 30576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_277
timestamp 1698431365
transform 1 0 32368 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_311
timestamp 1698431365
transform 1 0 36176 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_313
timestamp 1698431365
transform 1 0 36400 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_360
timestamp 1698431365
transform 1 0 41664 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_401
timestamp 1698431365
transform 1 0 46256 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_18
timestamp 1698431365
transform 1 0 3360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_24
timestamp 1698431365
transform 1 0 4032 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_32
timestamp 1698431365
transform 1 0 4928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_69
timestamp 1698431365
transform 1 0 9072 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_85
timestamp 1698431365
transform 1 0 10864 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_89
timestamp 1698431365
transform 1 0 11312 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_115
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_150
timestamp 1698431365
transform 1 0 18144 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_154
timestamp 1698431365
transform 1 0 18592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_156
timestamp 1698431365
transform 1 0 18816 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_173
timestamp 1698431365
transform 1 0 20720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_263
timestamp 1698431365
transform 1 0 30800 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_279
timestamp 1698431365
transform 1 0 32592 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_283
timestamp 1698431365
transform 1 0 33040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_285
timestamp 1698431365
transform 1 0 33264 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_399
timestamp 1698431365
transform 1 0 46032 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_401
timestamp 1698431365
transform 1 0 46256 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_38
timestamp 1698431365
transform 1 0 5600 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_54
timestamp 1698431365
transform 1 0 7392 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_58
timestamp 1698431365
transform 1 0 7840 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_64
timestamp 1698431365
transform 1 0 8512 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_68
timestamp 1698431365
transform 1 0 8960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_146
timestamp 1698431365
transform 1 0 17696 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_150
timestamp 1698431365
transform 1 0 18144 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_159
timestamp 1698431365
transform 1 0 19152 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_185
timestamp 1698431365
transform 1 0 22064 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_290
timestamp 1698431365
transform 1 0 33824 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_347
timestamp 1698431365
transform 1 0 40208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_356
timestamp 1698431365
transform 1 0 41216 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_358
timestamp 1698431365
transform 1 0 41440 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_367
timestamp 1698431365
transform 1 0 42448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_371
timestamp 1698431365
transform 1 0 42896 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_401
timestamp 1698431365
transform 1 0 46256 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_18
timestamp 1698431365
transform 1 0 3360 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_20
timestamp 1698431365
transform 1 0 3584 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_25
timestamp 1698431365
transform 1 0 4144 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_33
timestamp 1698431365
transform 1 0 5040 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_45
timestamp 1698431365
transform 1 0 6384 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_47
timestamp 1698431365
transform 1 0 6608 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_82
timestamp 1698431365
transform 1 0 10528 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_86
timestamp 1698431365
transform 1 0 10976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_113
timestamp 1698431365
transform 1 0 14000 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_115
timestamp 1698431365
transform 1 0 14224 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_130
timestamp 1698431365
transform 1 0 15904 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_163
timestamp 1698431365
transform 1 0 19600 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_167
timestamp 1698431365
transform 1 0 20048 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_209
timestamp 1698431365
transform 1 0 24752 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_266
timestamp 1698431365
transform 1 0 31136 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_270
timestamp 1698431365
transform 1 0 31584 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_345
timestamp 1698431365
transform 1 0 39984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_349
timestamp 1698431365
transform 1 0 40432 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_381
timestamp 1698431365
transform 1 0 44016 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_391
timestamp 1698431365
transform 1 0 45136 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_399
timestamp 1698431365
transform 1 0 46032 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_401
timestamp 1698431365
transform 1 0 46256 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_37
timestamp 1698431365
transform 1 0 5488 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_53
timestamp 1698431365
transform 1 0 7280 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_61
timestamp 1698431365
transform 1 0 8176 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_67
timestamp 1698431365
transform 1 0 8848 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_88
timestamp 1698431365
transform 1 0 11200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_90
timestamp 1698431365
transform 1 0 11424 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_137
timestamp 1698431365
transform 1 0 16688 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_139
timestamp 1698431365
transform 1 0 16912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_209
timestamp 1698431365
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_222
timestamp 1698431365
transform 1 0 26208 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_226
timestamp 1698431365
transform 1 0 26656 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_266
timestamp 1698431365
transform 1 0 31136 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_274
timestamp 1698431365
transform 1 0 32032 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_339
timestamp 1698431365
transform 1 0 39312 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_343
timestamp 1698431365
transform 1 0 39760 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_347
timestamp 1698431365
transform 1 0 40208 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_349
timestamp 1698431365
transform 1 0 40432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_356
timestamp 1698431365
transform 1 0 41216 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_394
timestamp 1698431365
transform 1 0 45472 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_18
timestamp 1698431365
transform 1 0 3360 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_28
timestamp 1698431365
transform 1 0 4480 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_85
timestamp 1698431365
transform 1 0 10864 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_156
timestamp 1698431365
transform 1 0 18816 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_172
timestamp 1698431365
transform 1 0 20608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_195
timestamp 1698431365
transform 1 0 23184 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_217
timestamp 1698431365
transform 1 0 25648 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_233
timestamp 1698431365
transform 1 0 27440 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_237
timestamp 1698431365
transform 1 0 27888 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_254
timestamp 1698431365
transform 1 0 29792 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_270
timestamp 1698431365
transform 1 0 31584 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_306
timestamp 1698431365
transform 1 0 35616 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698431365
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_326
timestamp 1698431365
transform 1 0 37856 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_395
timestamp 1698431365
transform 1 0 45584 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_399
timestamp 1698431365
transform 1 0 46032 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_401
timestamp 1698431365
transform 1 0 46256 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_76
timestamp 1698431365
transform 1 0 9856 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_120
timestamp 1698431365
transform 1 0 14784 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_124
timestamp 1698431365
transform 1 0 15232 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_158
timestamp 1698431365
transform 1 0 19040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_162
timestamp 1698431365
transform 1 0 19488 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_178
timestamp 1698431365
transform 1 0 21280 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_182
timestamp 1698431365
transform 1 0 21728 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_218
timestamp 1698431365
transform 1 0 25760 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_256
timestamp 1698431365
transform 1 0 30016 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_272
timestamp 1698431365
transform 1 0 31808 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_314
timestamp 1698431365
transform 1 0 36512 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_332
timestamp 1698431365
transform 1 0 38528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_8
timestamp 1698431365
transform 1 0 2240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_12
timestamp 1698431365
transform 1 0 2688 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_71
timestamp 1698431365
transform 1 0 9296 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_79
timestamp 1698431365
transform 1 0 10192 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_83
timestamp 1698431365
transform 1 0 10640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_85
timestamp 1698431365
transform 1 0 10864 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_92
timestamp 1698431365
transform 1 0 11648 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_100
timestamp 1698431365
transform 1 0 12544 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698431365
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_115
timestamp 1698431365
transform 1 0 14224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_149
timestamp 1698431365
transform 1 0 18032 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_165
timestamp 1698431365
transform 1 0 19824 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_181
timestamp 1698431365
transform 1 0 21616 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_223
timestamp 1698431365
transform 1 0 26320 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_227
timestamp 1698431365
transform 1 0 26768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_231
timestamp 1698431365
transform 1 0 27216 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_291
timestamp 1698431365
transform 1 0 33936 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_307
timestamp 1698431365
transform 1 0 35728 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_351
timestamp 1698431365
transform 1 0 40656 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_360
timestamp 1698431365
transform 1 0 41664 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_393
timestamp 1698431365
transform 1 0 45360 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_401
timestamp 1698431365
transform 1 0 46256 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_18
timestamp 1698431365
transform 1 0 3360 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_60
timestamp 1698431365
transform 1 0 8064 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_68
timestamp 1698431365
transform 1 0 8960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_76
timestamp 1698431365
transform 1 0 9856 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_122
timestamp 1698431365
transform 1 0 15008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_124
timestamp 1698431365
transform 1 0 15232 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_131
timestamp 1698431365
transform 1 0 16016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_133
timestamp 1698431365
transform 1 0 16240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_157
timestamp 1698431365
transform 1 0 18928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_161
timestamp 1698431365
transform 1 0 19376 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_208
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_290
timestamp 1698431365
transform 1 0 33824 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_300
timestamp 1698431365
transform 1 0 34944 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_342
timestamp 1698431365
transform 1 0 39648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_360
timestamp 1698431365
transform 1 0 41664 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_364
timestamp 1698431365
transform 1 0 42112 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_374
timestamp 1698431365
transform 1 0 43232 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_392
timestamp 1698431365
transform 1 0 45248 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_400
timestamp 1698431365
transform 1 0 46144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_18
timestamp 1698431365
transform 1 0 3360 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_26
timestamp 1698431365
transform 1 0 4256 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_30
timestamp 1698431365
transform 1 0 4704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_32
timestamp 1698431365
transform 1 0 4928 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_53
timestamp 1698431365
transform 1 0 7280 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_69
timestamp 1698431365
transform 1 0 9072 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_117
timestamp 1698431365
transform 1 0 14448 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_150
timestamp 1698431365
transform 1 0 18144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_152
timestamp 1698431365
transform 1 0 18368 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_179
timestamp 1698431365
transform 1 0 21392 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_194
timestamp 1698431365
transform 1 0 23072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_233
timestamp 1698431365
transform 1 0 27440 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_279
timestamp 1698431365
transform 1 0 32592 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_325
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_348
timestamp 1698431365
transform 1 0 40320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_356
timestamp 1698431365
transform 1 0 41216 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_364
timestamp 1698431365
transform 1 0 42112 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_368
timestamp 1698431365
transform 1 0 42560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_378
timestamp 1698431365
transform 1 0 43680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_382
timestamp 1698431365
transform 1 0 44128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_384
timestamp 1698431365
transform 1 0 44352 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_395
timestamp 1698431365
transform 1 0 45584 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_399
timestamp 1698431365
transform 1 0 46032 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_401
timestamp 1698431365
transform 1 0 46256 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_44
timestamp 1698431365
transform 1 0 6272 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_60
timestamp 1698431365
transform 1 0 8064 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_68
timestamp 1698431365
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_80
timestamp 1698431365
transform 1 0 10304 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_124
timestamp 1698431365
transform 1 0 15232 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_126
timestamp 1698431365
transform 1 0 15456 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_133
timestamp 1698431365
transform 1 0 16240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_137
timestamp 1698431365
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_150
timestamp 1698431365
transform 1 0 18144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_152
timestamp 1698431365
transform 1 0 18368 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_187
timestamp 1698431365
transform 1 0 22288 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_226
timestamp 1698431365
transform 1 0 26656 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_234
timestamp 1698431365
transform 1 0 27552 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_238
timestamp 1698431365
transform 1 0 28000 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_246
timestamp 1698431365
transform 1 0 28896 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_261
timestamp 1698431365
transform 1 0 30576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_290
timestamp 1698431365
transform 1 0 33824 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_334
timestamp 1698431365
transform 1 0 38752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_386
timestamp 1698431365
transform 1 0 44576 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_113
timestamp 1698431365
transform 1 0 14000 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_117
timestamp 1698431365
transform 1 0 14448 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_151
timestamp 1698431365
transform 1 0 18256 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_215
timestamp 1698431365
transform 1 0 25424 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_231
timestamp 1698431365
transform 1 0 27216 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_239
timestamp 1698431365
transform 1 0 28112 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_243
timestamp 1698431365
transform 1 0 28560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_263
timestamp 1698431365
transform 1 0 30800 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_313
timestamp 1698431365
transform 1 0 36400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_395
timestamp 1698431365
transform 1 0 45584 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_399
timestamp 1698431365
transform 1 0 46032 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_401
timestamp 1698431365
transform 1 0 46256 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_37
timestamp 1698431365
transform 1 0 5488 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698431365
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_80
timestamp 1698431365
transform 1 0 10304 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_84
timestamp 1698431365
transform 1 0 10752 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_86
timestamp 1698431365
transform 1 0 10976 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_134
timestamp 1698431365
transform 1 0 16352 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_138
timestamp 1698431365
transform 1 0 16800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_180
timestamp 1698431365
transform 1 0 21504 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_205
timestamp 1698431365
transform 1 0 24304 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_209
timestamp 1698431365
transform 1 0 24752 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_228
timestamp 1698431365
transform 1 0 26880 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_230
timestamp 1698431365
transform 1 0 27104 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_253
timestamp 1698431365
transform 1 0 29680 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_269
timestamp 1698431365
transform 1 0 31472 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_273
timestamp 1698431365
transform 1 0 31920 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_345
timestamp 1698431365
transform 1 0 39984 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_349
timestamp 1698431365
transform 1 0 40432 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_364
timestamp 1698431365
transform 1 0 42112 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_396
timestamp 1698431365
transform 1 0 45696 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_400
timestamp 1698431365
transform 1 0 46144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_53
timestamp 1698431365
transform 1 0 7280 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_61
timestamp 1698431365
transform 1 0 8176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_183
timestamp 1698431365
transform 1 0 21840 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_219
timestamp 1698431365
transform 1 0 25872 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_227
timestamp 1698431365
transform 1 0 26768 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_231
timestamp 1698431365
transform 1 0 27216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_233
timestamp 1698431365
transform 1 0 27440 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_242
timestamp 1698431365
transform 1 0 28448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_295
timestamp 1698431365
transform 1 0 34384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_299
timestamp 1698431365
transform 1 0 34832 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_342
timestamp 1698431365
transform 1 0 39648 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_374
timestamp 1698431365
transform 1 0 43232 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_382
timestamp 1698431365
transform 1 0 44128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_395
timestamp 1698431365
transform 1 0 45584 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_399
timestamp 1698431365
transform 1 0 46032 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_401
timestamp 1698431365
transform 1 0 46256 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_80
timestamp 1698431365
transform 1 0 10304 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_84
timestamp 1698431365
transform 1 0 10752 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_135
timestamp 1698431365
transform 1 0 16464 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_139
timestamp 1698431365
transform 1 0 16912 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_156
timestamp 1698431365
transform 1 0 18816 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_158
timestamp 1698431365
transform 1 0 19040 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_197
timestamp 1698431365
transform 1 0 23408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_205
timestamp 1698431365
transform 1 0 24304 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_220
timestamp 1698431365
transform 1 0 25984 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_224
timestamp 1698431365
transform 1 0 26432 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_274
timestamp 1698431365
transform 1 0 32032 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_278
timestamp 1698431365
transform 1 0 32480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_298
timestamp 1698431365
transform 1 0 34720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_334
timestamp 1698431365
transform 1 0 38752 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_384
timestamp 1698431365
transform 1 0 44352 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_400
timestamp 1698431365
transform 1 0 46144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_69
timestamp 1698431365
transform 1 0 9072 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_85
timestamp 1698431365
transform 1 0 10864 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_93
timestamp 1698431365
transform 1 0 11760 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_97
timestamp 1698431365
transform 1 0 12208 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_152
timestamp 1698431365
transform 1 0 18368 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_156
timestamp 1698431365
transform 1 0 18816 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_165
timestamp 1698431365
transform 1 0 19824 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_173
timestamp 1698431365
transform 1 0 20720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_185
timestamp 1698431365
transform 1 0 22064 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_189
timestamp 1698431365
transform 1 0 22512 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_242
timestamp 1698431365
transform 1 0 28448 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_244
timestamp 1698431365
transform 1 0 28672 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_279
timestamp 1698431365
transform 1 0 32592 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698431365
transform 1 0 44016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_395
timestamp 1698431365
transform 1 0 45584 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_399
timestamp 1698431365
transform 1 0 46032 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_401
timestamp 1698431365
transform 1 0 46256 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698431365
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_88
timestamp 1698431365
transform 1 0 11200 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_96
timestamp 1698431365
transform 1 0 12096 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_100
timestamp 1698431365
transform 1 0 12544 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_150
timestamp 1698431365
transform 1 0 18144 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_154
timestamp 1698431365
transform 1 0 18592 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_205
timestamp 1698431365
transform 1 0 24304 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_209
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_216
timestamp 1698431365
transform 1 0 25536 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_291
timestamp 1698431365
transform 1 0 33936 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_323
timestamp 1698431365
transform 1 0 37520 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_339
timestamp 1698431365
transform 1 0 39312 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_347
timestamp 1698431365
transform 1 0 40208 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_349
timestamp 1698431365
transform 1 0 40432 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_384
timestamp 1698431365
transform 1 0 44352 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_400
timestamp 1698431365
transform 1 0 46144 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_6
timestamp 1698431365
transform 1 0 2016 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_22
timestamp 1698431365
transform 1 0 3808 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_30
timestamp 1698431365
transform 1 0 4704 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_101
timestamp 1698431365
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_161
timestamp 1698431365
transform 1 0 19376 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_181
timestamp 1698431365
transform 1 0 21616 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_228
timestamp 1698431365
transform 1 0 26880 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_305
timestamp 1698431365
transform 1 0 35504 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_313
timestamp 1698431365
transform 1 0 36400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698431365
transform 1 0 44016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_395
timestamp 1698431365
transform 1 0 45584 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_397
timestamp 1698431365
transform 1 0 45808 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_6
timestamp 1698431365
transform 1 0 2016 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_88
timestamp 1698431365
transform 1 0 11200 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_96
timestamp 1698431365
transform 1 0 12096 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_100
timestamp 1698431365
transform 1 0 12544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_108
timestamp 1698431365
transform 1 0 13440 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_150
timestamp 1698431365
transform 1 0 18144 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_154
timestamp 1698431365
transform 1 0 18592 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_156
timestamp 1698431365
transform 1 0 18816 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_193
timestamp 1698431365
transform 1 0 22960 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_234
timestamp 1698431365
transform 1 0 27552 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_265
timestamp 1698431365
transform 1 0 31024 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_273
timestamp 1698431365
transform 1 0 31920 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_277
timestamp 1698431365
transform 1 0 32368 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1698431365
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_346
timestamp 1698431365
transform 1 0 40096 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_384
timestamp 1698431365
transform 1 0 44352 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_400
timestamp 1698431365
transform 1 0 46144 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_36
timestamp 1698431365
transform 1 0 5376 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_70
timestamp 1698431365
transform 1 0 9184 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_104
timestamp 1698431365
transform 1 0 12992 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_138
timestamp 1698431365
transform 1 0 16800 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_172
timestamp 1698431365
transform 1 0 20608 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_206
timestamp 1698431365
transform 1 0 24416 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_240
timestamp 1698431365
transform 1 0 28224 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_274
timestamp 1698431365
transform 1 0 32032 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_308
timestamp 1698431365
transform 1 0 35840 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_342
timestamp 1698431365
transform 1 0 39648 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_376
timestamp 1698431365
transform 1 0 43456 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_392
timestamp 1698431365
transform 1 0 45248 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_400
timestamp 1698431365
transform 1 0 46144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 2240 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input6
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input7
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input8
timestamp 1698431365
transform 1 0 3360 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698431365
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698431365
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698431365
transform -1 0 8400 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698431365
transform -1 0 4480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698431365
transform -1 0 4480 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698431365
transform -1 0 4480 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698431365
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_53 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 46592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 46592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 46592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 46592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 46592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 46592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 46592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 46592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 46592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 46592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 46592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 46592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 46592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 46592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 46592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 46592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 46592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 46592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 46592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 46592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 46592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 46592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 46592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 46592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 46592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 46592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 46592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 46592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 46592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 46592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 46592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 46592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 46592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 46592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 46592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 46592 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 46592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 46592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 46592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 46592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 46592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 46592 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 46592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 46592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 46592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 46592 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 46592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 46592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 46592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 46592 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 46592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 46592 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 46592 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ro_inst.clock_gate_315
timestamp 1698431365
transform -1 0 8176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__icgtp_1  ro_inst.clock_gate
timestamp 1698431365
transform 1 0 7728 0 1 26656
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.clock_gate_inv
timestamp 1698431365
transform -1 0 4928 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[1\].div_flop_inv
timestamp 1698431365
transform -1 0 4928 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[1\].div_flop
timestamp 1698431365
transform 1 0 2464 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[2\].div_flop
timestamp 1698431365
transform 1 0 2128 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[2\].div_flop_inv
timestamp 1698431365
transform 1 0 1680 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[3\].div_flop_inv
timestamp 1698431365
transform -1 0 8848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[3\].div_flop
timestamp 1698431365
transform 1 0 1792 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[4\].div_flop
timestamp 1698431365
transform 1 0 1904 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[4\].div_flop_inv
timestamp 1698431365
transform -1 0 4368 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[5\].div_flop
timestamp 1698431365
transform 1 0 2352 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[5\].div_flop_inv
timestamp 1698431365
transform -1 0 4816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[6\].div_flop
timestamp 1698431365
transform 1 0 2688 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[6\].div_flop_inv
timestamp 1698431365
transform -1 0 5264 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[7\].div_flop
timestamp 1698431365
transform 1 0 5376 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[7\].div_flop_inv
timestamp 1698431365
transform -1 0 6272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[8\].div_flop
timestamp 1698431365
transform 1 0 4816 0 -1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[8\].div_flop_inv
timestamp 1698431365
transform -1 0 7504 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[9\].div_flop
timestamp 1698431365
transform 1 0 5376 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[9\].div_flop_inv
timestamp 1698431365
transform -1 0 8848 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[10\].div_flop_inv
timestamp 1698431365
transform -1 0 9856 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[10\].div_flop
timestamp 1698431365
transform 1 0 7280 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[11\].div_flop_inv
timestamp 1698431365
transform -1 0 10304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[11\].div_flop
timestamp 1698431365
transform 1 0 7728 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[12\].div_flop
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[12\].div_flop_inv
timestamp 1698431365
transform -1 0 10192 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[13\].div_flop
timestamp 1698431365
transform -1 0 9184 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[13\].div_flop_inv
timestamp 1698431365
transform 1 0 5824 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[14\].div_flop_inv
timestamp 1698431365
transform -1 0 5152 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[14\].div_flop
timestamp 1698431365
transform -1 0 6720 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[15\].div_flop_inv
timestamp 1698431365
transform -1 0 4480 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[15\].div_flop
timestamp 1698431365
transform 1 0 2128 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[16\].div_flop_inv
timestamp 1698431365
transform -1 0 4368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[16\].div_flop
timestamp 1698431365
transform 1 0 1792 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[17\].div_flop
timestamp 1698431365
transform -1 0 9184 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[17\].div_flop_inv
timestamp 1698431365
transform -1 0 3920 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[18\].div_flop_inv
timestamp 1698431365
transform -1 0 3808 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[18\].div_flop
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[19\].div_flop_inv
timestamp 1698431365
transform -1 0 3808 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[19\].div_flop
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[20\].div_flop_inv
timestamp 1698431365
transform -1 0 3808 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[20\].div_flop
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[21\].div_flop
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[21\].div_flop_inv
timestamp 1698431365
transform -1 0 3808 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[22\].div_flop_inv
timestamp 1698431365
transform -1 0 5264 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[22\].div_flop
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[23\].div_flop_inv
timestamp 1698431365
transform -1 0 5936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[23\].div_flop
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[24\].div_flop
timestamp 1698431365
transform 1 0 1680 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[24\].div_flop_inv
timestamp 1698431365
transform -1 0 4032 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[25\].div_flop_inv
timestamp 1698431365
transform -1 0 4144 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[25\].div_flop
timestamp 1698431365
transform 1 0 1792 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[26\].div_flop_inv
timestamp 1698431365
transform -1 0 4032 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[26\].div_flop
timestamp 1698431365
transform 1 0 1680 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[27\].div_flop
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[27\].div_flop_inv
timestamp 1698431365
transform -1 0 4480 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[28\].div_flop
timestamp 1698431365
transform 1 0 1680 0 -1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[28\].div_flop_inv
timestamp 1698431365
transform -1 0 3248 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[29\].div_flop
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[29\].div_flop_inv
timestamp 1698431365
transform -1 0 5152 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[30\].div_flop_inv
timestamp 1698431365
transform -1 0 7280 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[30\].div_flop
timestamp 1698431365
transform 1 0 3808 0 -1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[31\].div_flop_inv
timestamp 1698431365
transform -1 0 8064 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[31\].div_flop
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[32\].div_flop_inv
timestamp 1698431365
transform -1 0 9856 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[32\].div_flop
timestamp 1698431365
transform 1 0 5376 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[33\].div_flop
timestamp 1698431365
transform 1 0 6384 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[33\].div_flop_inv
timestamp 1698431365
transform -1 0 8848 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  ro_inst.gcount\[34\].div_flop
timestamp 1698431365
transform 1 0 6720 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.gcount\[34\].div_flop_inv
timestamp 1698431365
transform -1 0 8512 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  ro_inst.ring_osc_0
timestamp 1698431365
transform 1 0 10864 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.ring_osc_1
timestamp 1698431365
transform -1 0 11872 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.ring_osc_2
timestamp 1698431365
transform -1 0 10304 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  ro_inst.sig_cmp
timestamp 1698431365
transform -1 0 9072 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  ro_inst.sig_latch
timestamp 1698431365
transform 1 0 6944 0 -1 28224
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ro_inst.slow_clock_inv
timestamp 1698431365
transform 1 0 6496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_106 test/tapeout/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_108
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_109
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_117
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_118
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_119
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_120
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_121
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_122
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_123
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_124
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_125
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_126
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_127
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_128
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_129
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_130
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_131
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_132
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_133
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_134
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_135
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_136
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_137
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_138
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_139
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_140
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_141
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_142
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_143
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_144
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_145
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_146
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_147
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_148
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_149
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_150
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_151
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_152
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_153
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_154
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_155
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_156
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_157
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_158
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_159
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_160
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_161
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_162
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_163
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_164
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_165
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_166
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_167
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_168
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_169
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_170
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_171
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_172
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_173
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_174
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_175
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_176
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_177
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_178
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_179
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_180
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_181
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_183
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_184
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_185
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_186
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_187
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_188
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_189
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_190
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_191
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_192
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_193
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_194
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_195
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_196
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_197
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_198
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_199
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_200
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_201
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_202
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_203
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_204
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_205
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_206
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_207
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_208
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_209
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_210
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_211
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_212
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_213
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_214
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_215
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_216
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_217
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_218
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_219
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_220
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_221
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_222
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_223
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_224
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_225
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_226
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_227
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_228
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_229
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_230
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_231
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_232
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_233
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_234
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_235
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_236
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_237
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_238
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_239
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_240
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_241
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_242
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_243
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_244
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_245
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_246
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_247
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_248
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_249
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_250
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_251
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_252
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_253
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_254
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_255
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_256
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_257
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_258
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_259
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_260
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_261
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_262
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_263
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_264
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_265
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_266
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_267
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_268
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_269
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_270
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_271
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_272
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_273
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_274
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_275
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_276
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_277
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_278
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_279
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_280
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_281
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_282
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_283
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_284
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_285
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_286
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_287
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_288
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_289
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_290
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_291
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_292
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_293
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_294
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_295
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_296
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_297
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_298
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_299
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_300
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_301
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_302
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_303
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_304
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_305
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_306
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_307
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_308
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_309
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_310
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_311
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_312
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_313
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_314
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_315
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_316
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_317
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_318
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_319
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_320
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_321
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_322
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_323
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_324
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_325
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_326
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_327
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_328
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_329
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_330
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_331
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_332
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_333
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_334
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_335
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_336
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_337
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_338
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_339
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_340
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_341
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_342
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_343
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_344
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_345
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_346
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_347
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_348
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_349
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_350
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_351
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_352
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_353
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_354
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_355
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_356
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_357
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_358
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_359
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_360
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_361
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_362
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_363
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_364
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_365
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_366
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_367
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_368
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_369
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_370
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_371
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_372
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_373
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_374
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_375
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_376
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_377
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_378
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_379
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_380
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_381
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_382
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_383
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_384
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_385
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_386
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_387
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_388
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_389
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_390
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_391
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_392
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_393
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_394
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_395
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_396
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_397
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_398
timestamp 1698431365
transform 1 0 8960 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_399
timestamp 1698431365
transform 1 0 12768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_400
timestamp 1698431365
transform 1 0 16576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_401
timestamp 1698431365
transform 1 0 20384 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_402
timestamp 1698431365
transform 1 0 24192 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_403
timestamp 1698431365
transform 1 0 28000 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_404
timestamp 1698431365
transform 1 0 31808 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_405
timestamp 1698431365
transform 1 0 35616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_406
timestamp 1698431365
transform 1 0 39424 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_407
timestamp 1698431365
transform 1 0 43232 0 1 43904
box -86 -86 310 870
<< labels >>
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 34272 800 34384 0 FreeSans 448 0 0 0 in[0]
port 1 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 in[10]
port 2 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 in[11]
port 3 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 in[12]
port 4 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 in[13]
port 5 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 in[14]
port 6 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 in[15]
port 7 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 in[16]
port 8 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 in[17]
port 9 nsew signal input
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 in[1]
port 10 nsew signal input
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 in[2]
port 11 nsew signal input
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 in[3]
port 12 nsew signal input
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 in[4]
port 13 nsew signal input
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 in[5]
port 14 nsew signal input
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 in[6]
port 15 nsew signal input
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 in[7]
port 16 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 in[8]
port 17 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 in[9]
port 18 nsew signal input
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 out[0]
port 19 nsew signal tristate
flabel metal3 s 47200 42336 48000 42448 0 FreeSans 448 0 0 0 out[10]
port 20 nsew signal tristate
flabel metal3 s 0 43008 800 43120 0 FreeSans 448 0 0 0 out[11]
port 21 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 out[1]
port 22 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 out[2]
port 23 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 out[3]
port 24 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 out[4]
port 25 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 out[5]
port 26 nsew signal tristate
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 out[6]
port 27 nsew signal tristate
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 out[7]
port 28 nsew signal tristate
flabel metal3 s 0 42336 800 42448 0 FreeSans 448 0 0 0 out[8]
port 29 nsew signal tristate
flabel metal3 s 0 4704 800 4816 0 FreeSans 448 0 0 0 out[9]
port 30 nsew signal tristate
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 rst_n
port 31 nsew signal input
flabel metal4 s 4448 3076 4768 44748 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 35168 3076 35488 44748 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 19808 3076 20128 44748 0 FreeSans 1280 90 0 0 vss
port 33 nsew ground bidirectional
rlabel metal1 23968 44688 23968 44688 0 vdd
rlabel metal1 23968 43904 23968 43904 0 vss
rlabel metal3 17360 19096 17360 19096 0 _000_
rlabel metal2 14728 15008 14728 15008 0 _001_
rlabel metal2 14616 24696 14616 24696 0 _002_
rlabel metal2 15064 21840 15064 21840 0 _003_
rlabel metal3 16128 22456 16128 22456 0 _004_
rlabel metal2 16072 21896 16072 21896 0 _005_
rlabel metal3 11256 14616 11256 14616 0 _006_
rlabel metal2 11144 14616 11144 14616 0 _007_
rlabel metal3 9688 18424 9688 18424 0 _008_
rlabel metal3 16688 20664 16688 20664 0 _009_
rlabel metal2 15736 17640 15736 17640 0 _010_
rlabel metal2 14840 17808 14840 17808 0 _011_
rlabel metal3 11648 24696 11648 24696 0 _012_
rlabel metal2 8008 19712 8008 19712 0 _013_
rlabel metal2 8232 16856 8232 16856 0 _014_
rlabel metal2 9576 20440 9576 20440 0 _015_
rlabel metal2 17640 21896 17640 21896 0 _016_
rlabel metal2 25704 24304 25704 24304 0 _017_
rlabel metal2 22736 18424 22736 18424 0 _018_
rlabel metal2 40040 27104 40040 27104 0 _019_
rlabel metal2 38808 32424 38808 32424 0 _020_
rlabel metal2 35672 25088 35672 25088 0 _021_
rlabel metal2 35224 25312 35224 25312 0 _022_
rlabel metal2 43624 29456 43624 29456 0 _023_
rlabel metal2 42952 29064 42952 29064 0 _024_
rlabel metal2 29736 23912 29736 23912 0 _025_
rlabel metal3 22568 34216 22568 34216 0 _026_
rlabel metal2 26376 30240 26376 30240 0 _027_
rlabel metal3 30520 27160 30520 27160 0 _028_
rlabel metal2 30408 26488 30408 26488 0 _029_
rlabel metal2 24024 24920 24024 24920 0 _030_
rlabel metal2 24696 21112 24696 21112 0 _031_
rlabel metal3 37576 25144 37576 25144 0 _032_
rlabel metal2 19376 26488 19376 26488 0 _033_
rlabel metal2 26600 26320 26600 26320 0 _034_
rlabel metal2 21224 23688 21224 23688 0 _035_
rlabel metal3 16912 24696 16912 24696 0 _036_
rlabel metal2 24136 17808 24136 17808 0 _037_
rlabel metal2 40208 12936 40208 12936 0 _038_
rlabel metal3 24360 12712 24360 12712 0 _039_
rlabel metal2 41384 12600 41384 12600 0 _040_
rlabel metal2 40936 13048 40936 13048 0 _041_
rlabel metal2 34888 11368 34888 11368 0 _042_
rlabel metal2 39480 11592 39480 11592 0 _043_
rlabel metal2 39704 25032 39704 25032 0 _044_
rlabel metal3 39592 13944 39592 13944 0 _045_
rlabel metal2 22568 26096 22568 26096 0 _046_
rlabel metal2 21336 25424 21336 25424 0 _047_
rlabel metal3 19768 17528 19768 17528 0 _048_
rlabel metal2 21784 32648 21784 32648 0 _049_
rlabel metal2 19208 24248 19208 24248 0 _050_
rlabel metal3 17136 8232 17136 8232 0 _051_
rlabel metal3 23688 18424 23688 18424 0 _052_
rlabel metal3 22736 16744 22736 16744 0 _053_
rlabel metal2 22568 17360 22568 17360 0 _054_
rlabel metal2 22904 17640 22904 17640 0 _055_
rlabel metal2 22008 15792 22008 15792 0 _056_
rlabel metal2 22232 17304 22232 17304 0 _057_
rlabel metal2 22120 23912 22120 23912 0 _058_
rlabel metal2 17864 23520 17864 23520 0 _059_
rlabel metal2 23464 22344 23464 22344 0 _060_
rlabel metal2 21560 23352 21560 23352 0 _061_
rlabel metal2 12824 23744 12824 23744 0 _062_
rlabel metal2 8456 23968 8456 23968 0 _063_
rlabel metal2 10808 25088 10808 25088 0 _064_
rlabel metal2 18200 24136 18200 24136 0 _065_
rlabel metal2 24640 25480 24640 25480 0 _066_
rlabel metal2 22120 21616 22120 21616 0 _067_
rlabel metal2 17640 32704 17640 32704 0 _068_
rlabel metal3 19376 15848 19376 15848 0 _069_
rlabel metal2 16184 9352 16184 9352 0 _070_
rlabel metal2 18984 11144 18984 11144 0 _071_
rlabel metal2 22904 5768 22904 5768 0 _072_
rlabel metal2 19656 6048 19656 6048 0 _073_
rlabel metal2 23128 10752 23128 10752 0 _074_
rlabel metal2 20328 21336 20328 21336 0 _075_
rlabel metal2 14504 24416 14504 24416 0 _076_
rlabel metal3 41944 24136 41944 24136 0 _077_
rlabel metal3 26712 23688 26712 23688 0 _078_
rlabel metal2 24584 26040 24584 26040 0 _079_
rlabel metal2 26152 21280 26152 21280 0 _080_
rlabel metal2 24696 15148 24696 15148 0 _081_
rlabel metal2 25480 8960 25480 8960 0 _082_
rlabel metal3 26432 22008 26432 22008 0 _083_
rlabel metal2 25928 22792 25928 22792 0 _084_
rlabel via2 26376 25592 26376 25592 0 _085_
rlabel metal2 21000 21616 21000 21616 0 _086_
rlabel metal3 19992 21784 19992 21784 0 _087_
rlabel metal3 22680 26264 22680 26264 0 _088_
rlabel metal2 25592 30912 25592 30912 0 _089_
rlabel metal2 24136 39144 24136 39144 0 _090_
rlabel metal2 26712 36008 26712 36008 0 _091_
rlabel metal2 27160 40768 27160 40768 0 _092_
rlabel metal2 25928 36792 25928 36792 0 _093_
rlabel metal2 19320 33936 19320 33936 0 _094_
rlabel metal3 25256 25368 25256 25368 0 _095_
rlabel metal2 22456 15904 22456 15904 0 _096_
rlabel metal2 20944 16408 20944 16408 0 _097_
rlabel metal2 20216 17024 20216 17024 0 _098_
rlabel metal3 22008 25480 22008 25480 0 _099_
rlabel metal2 21336 26208 21336 26208 0 _100_
rlabel metal2 21000 24976 21000 24976 0 _101_
rlabel metal3 19824 23912 19824 23912 0 _102_
rlabel metal2 11928 24248 11928 24248 0 _103_
rlabel metal2 7560 24696 7560 24696 0 _104_
rlabel metal2 41104 32760 41104 32760 0 _105_
rlabel metal3 43288 20160 43288 20160 0 _106_
rlabel metal2 40264 25032 40264 25032 0 _107_
rlabel metal2 41272 37296 41272 37296 0 _108_
rlabel metal2 42784 33320 42784 33320 0 _109_
rlabel metal2 43736 27944 43736 27944 0 _110_
rlabel metal2 26824 24640 26824 24640 0 _111_
rlabel metal2 27552 23352 27552 23352 0 _112_
rlabel metal2 26040 28952 26040 28952 0 _113_
rlabel metal2 26152 27328 26152 27328 0 _114_
rlabel metal2 14952 36176 14952 36176 0 _115_
rlabel metal3 17808 38248 17808 38248 0 _116_
rlabel metal2 24416 26376 24416 26376 0 _117_
rlabel metal3 25312 26488 25312 26488 0 _118_
rlabel metal2 26040 25760 26040 25760 0 _119_
rlabel metal3 25200 24696 25200 24696 0 _120_
rlabel metal2 38248 21168 38248 21168 0 _121_
rlabel metal2 37520 22568 37520 22568 0 _122_
rlabel metal2 24584 23296 24584 23296 0 _123_
rlabel metal2 20552 28224 20552 28224 0 _124_
rlabel metal2 22680 23016 22680 23016 0 _125_
rlabel metal2 23464 19880 23464 19880 0 _126_
rlabel metal2 24024 23968 24024 23968 0 _127_
rlabel metal2 8792 23520 8792 23520 0 _128_
rlabel metal3 7056 23352 7056 23352 0 _129_
rlabel metal2 22456 6160 22456 6160 0 _130_
rlabel metal3 24192 9688 24192 9688 0 _131_
rlabel metal3 22400 18648 22400 18648 0 _132_
rlabel metal2 31192 21000 31192 21000 0 _133_
rlabel metal2 27048 21504 27048 21504 0 _134_
rlabel metal2 32536 18200 32536 18200 0 _135_
rlabel metal2 28168 17892 28168 17892 0 _136_
rlabel metal2 27832 21280 27832 21280 0 _137_
rlabel metal2 26712 22680 26712 22680 0 _138_
rlabel metal2 27160 21336 27160 21336 0 _139_
rlabel metal2 20608 25480 20608 25480 0 _140_
rlabel metal2 15848 37296 15848 37296 0 _141_
rlabel metal2 15624 35112 15624 35112 0 _142_
rlabel metal2 18872 31192 18872 31192 0 _143_
rlabel metal2 12712 27888 12712 27888 0 _144_
rlabel metal2 11816 27832 11816 27832 0 _145_
rlabel metal2 19096 26152 19096 26152 0 _146_
rlabel metal2 7000 23352 7000 23352 0 _147_
rlabel metal2 6888 23184 6888 23184 0 _148_
rlabel metal3 5432 23352 5432 23352 0 _149_
rlabel metal2 32760 16184 32760 16184 0 _150_
rlabel metal2 34048 16632 34048 16632 0 _151_
rlabel metal3 26684 23912 26684 23912 0 _152_
rlabel metal3 25200 26040 25200 26040 0 _153_
rlabel metal3 24696 25480 24696 25480 0 _154_
rlabel metal2 25256 28112 25256 28112 0 _155_
rlabel metal2 25368 25760 25368 25760 0 _156_
rlabel metal2 25032 24024 25032 24024 0 _157_
rlabel metal2 23128 21840 23128 21840 0 _158_
rlabel metal3 37912 15848 37912 15848 0 _159_
rlabel metal2 34048 9688 34048 9688 0 _160_
rlabel metal3 25620 22232 25620 22232 0 _161_
rlabel metal2 22736 21000 22736 21000 0 _162_
rlabel metal2 23240 21784 23240 21784 0 _163_
rlabel metal2 12824 22680 12824 22680 0 _164_
rlabel metal3 5376 22344 5376 22344 0 _165_
rlabel metal2 17080 11760 17080 11760 0 _166_
rlabel metal2 19544 10976 19544 10976 0 _167_
rlabel metal2 20384 17416 20384 17416 0 _168_
rlabel metal2 40712 26096 40712 26096 0 _169_
rlabel metal2 26488 23408 26488 23408 0 _170_
rlabel metal2 26432 21336 26432 21336 0 _171_
rlabel metal2 26320 21784 26320 21784 0 _172_
rlabel metal2 20888 21000 20888 21000 0 _173_
rlabel metal3 19992 20888 19992 20888 0 _174_
rlabel metal2 24024 39928 24024 39928 0 _175_
rlabel metal2 23240 39088 23240 39088 0 _176_
rlabel metal2 22904 38024 22904 38024 0 _177_
rlabel metal2 20888 28112 20888 28112 0 _178_
rlabel metal2 21000 25368 21000 25368 0 _179_
rlabel metal2 11984 23128 11984 23128 0 _180_
rlabel metal2 6384 21784 6384 21784 0 _181_
rlabel metal2 36288 26936 36288 26936 0 _182_
rlabel metal2 35504 27272 35504 27272 0 _183_
rlabel metal2 26824 26544 26824 26544 0 _184_
rlabel metal2 27272 29960 27272 29960 0 _185_
rlabel metal2 26936 27440 26936 27440 0 _186_
rlabel metal2 23128 28896 23128 28896 0 _187_
rlabel metal2 24920 27720 24920 27720 0 _188_
rlabel metal2 25256 26544 25256 26544 0 _189_
rlabel metal2 18648 26208 18648 26208 0 _190_
rlabel metal2 42056 32032 42056 32032 0 _191_
rlabel metal2 37464 30632 37464 30632 0 _192_
rlabel metal3 23016 26376 23016 26376 0 _193_
rlabel metal2 20832 26264 20832 26264 0 _194_
rlabel metal2 19768 26320 19768 26320 0 _195_
rlabel metal2 9688 23352 9688 23352 0 _196_
rlabel metal2 10472 28112 10472 28112 0 _197_
rlabel metal2 22344 7336 22344 7336 0 _198_
rlabel metal3 24920 7672 24920 7672 0 _199_
rlabel metal2 22008 17304 22008 17304 0 _200_
rlabel metal3 29176 21672 29176 21672 0 _201_
rlabel metal2 27720 21672 27720 21672 0 _202_
rlabel metal3 33152 20104 33152 20104 0 _203_
rlabel metal2 27440 20888 27440 20888 0 _204_
rlabel metal2 27160 21952 27160 21952 0 _205_
rlabel metal2 22512 24696 22512 24696 0 _206_
rlabel metal2 18480 38920 18480 38920 0 _207_
rlabel metal2 17192 32760 17192 32760 0 _208_
rlabel metal2 21448 27496 21448 27496 0 _209_
rlabel metal2 22232 27328 22232 27328 0 _210_
rlabel metal2 22232 25704 22232 25704 0 _211_
rlabel metal3 10640 23128 10640 23128 0 _212_
rlabel metal2 9744 26488 9744 26488 0 _213_
rlabel metal2 10584 22960 10584 22960 0 _214_
rlabel metal2 9912 22904 9912 22904 0 _215_
rlabel metal2 9464 22568 9464 22568 0 _216_
rlabel metal2 14952 21280 14952 21280 0 _217_
rlabel metal2 13048 18704 13048 18704 0 _218_
rlabel metal2 14280 19208 14280 19208 0 _219_
rlabel metal2 14504 19376 14504 19376 0 _220_
rlabel metal2 16856 19040 16856 19040 0 _221_
rlabel metal3 13888 23912 13888 23912 0 _222_
rlabel metal2 13160 16296 13160 16296 0 _223_
rlabel metal2 14112 15288 14112 15288 0 _224_
rlabel metal2 13720 23128 13720 23128 0 _225_
rlabel metal3 11088 20104 11088 20104 0 _226_
rlabel metal2 14840 21168 14840 21168 0 _227_
rlabel metal2 14952 23408 14952 23408 0 _228_
rlabel metal3 16856 21560 16856 21560 0 _229_
rlabel metal2 12936 17584 12936 17584 0 _230_
rlabel metal2 10360 15960 10360 15960 0 _231_
rlabel metal2 11256 15624 11256 15624 0 _232_
rlabel metal2 8792 19096 8792 19096 0 _233_
rlabel metal2 14952 22344 14952 22344 0 _234_
rlabel metal2 13384 18032 13384 18032 0 _235_
rlabel metal3 16464 18424 16464 18424 0 _236_
rlabel metal2 13384 24864 13384 24864 0 _237_
rlabel metal2 12152 20468 12152 20468 0 _238_
rlabel metal2 10584 19712 10584 19712 0 _239_
rlabel metal2 8120 18144 8120 18144 0 _240_
rlabel metal3 10472 20552 10472 20552 0 _241_
rlabel metal2 9800 16072 9800 16072 0 cm_inst.cc_inst.in\[0\]
rlabel metal2 13272 13664 13272 13664 0 cm_inst.cc_inst.in\[1\]
rlabel metal2 12544 21560 12544 21560 0 cm_inst.cc_inst.in\[2\]
rlabel metal2 13944 22008 13944 22008 0 cm_inst.cc_inst.in\[3\]
rlabel metal2 13608 17024 13608 17024 0 cm_inst.cc_inst.in\[4\]
rlabel metal2 16968 18088 16968 18088 0 cm_inst.cc_inst.in\[5\]
rlabel metal2 33096 25312 33096 25312 0 cm_inst.cc_inst.out_notouch_\[0\]
rlabel metal2 34888 15624 34888 15624 0 cm_inst.cc_inst.out_notouch_\[100\]
rlabel metal2 42840 27384 42840 27384 0 cm_inst.cc_inst.out_notouch_\[101\]
rlabel metal2 38360 27552 38360 27552 0 cm_inst.cc_inst.out_notouch_\[102\]
rlabel metal2 32424 22064 32424 22064 0 cm_inst.cc_inst.out_notouch_\[103\]
rlabel metal2 36344 23800 36344 23800 0 cm_inst.cc_inst.out_notouch_\[104\]
rlabel metal2 42952 23912 42952 23912 0 cm_inst.cc_inst.out_notouch_\[105\]
rlabel metal2 42056 24416 42056 24416 0 cm_inst.cc_inst.out_notouch_\[106\]
rlabel metal2 32424 19936 32424 19936 0 cm_inst.cc_inst.out_notouch_\[107\]
rlabel metal2 33768 16408 33768 16408 0 cm_inst.cc_inst.out_notouch_\[108\]
rlabel metal2 41832 27720 41832 27720 0 cm_inst.cc_inst.out_notouch_\[109\]
rlabel metal3 27440 30184 27440 30184 0 cm_inst.cc_inst.out_notouch_\[10\]
rlabel metal2 37464 28112 37464 28112 0 cm_inst.cc_inst.out_notouch_\[110\]
rlabel metal3 32256 21560 32256 21560 0 cm_inst.cc_inst.out_notouch_\[111\]
rlabel metal2 34720 21784 34720 21784 0 cm_inst.cc_inst.out_notouch_\[112\]
rlabel metal2 40936 24360 40936 24360 0 cm_inst.cc_inst.out_notouch_\[113\]
rlabel metal2 40488 24640 40488 24640 0 cm_inst.cc_inst.out_notouch_\[114\]
rlabel metal2 30296 17752 30296 17752 0 cm_inst.cc_inst.out_notouch_\[115\]
rlabel metal2 31752 16408 31752 16408 0 cm_inst.cc_inst.out_notouch_\[116\]
rlabel metal2 39536 27160 39536 27160 0 cm_inst.cc_inst.out_notouch_\[117\]
rlabel metal2 35224 27944 35224 27944 0 cm_inst.cc_inst.out_notouch_\[118\]
rlabel metal2 29288 21840 29288 21840 0 cm_inst.cc_inst.out_notouch_\[119\]
rlabel metal2 26152 9464 26152 9464 0 cm_inst.cc_inst.out_notouch_\[11\]
rlabel metal2 34216 23968 34216 23968 0 cm_inst.cc_inst.out_notouch_\[120\]
rlabel metal2 41888 24024 41888 24024 0 cm_inst.cc_inst.out_notouch_\[121\]
rlabel metal2 41384 23968 41384 23968 0 cm_inst.cc_inst.out_notouch_\[122\]
rlabel metal2 30856 20496 30856 20496 0 cm_inst.cc_inst.out_notouch_\[123\]
rlabel metal2 32424 15792 32424 15792 0 cm_inst.cc_inst.out_notouch_\[124\]
rlabel metal2 40320 27048 40320 27048 0 cm_inst.cc_inst.out_notouch_\[125\]
rlabel metal2 36120 28504 36120 28504 0 cm_inst.cc_inst.out_notouch_\[126\]
rlabel metal2 30072 21952 30072 21952 0 cm_inst.cc_inst.out_notouch_\[127\]
rlabel metal2 41608 9520 41608 9520 0 cm_inst.cc_inst.out_notouch_\[128\]
rlabel metal2 30016 40376 30016 40376 0 cm_inst.cc_inst.out_notouch_\[129\]
rlabel metal2 27384 30296 27384 30296 0 cm_inst.cc_inst.out_notouch_\[12\]
rlabel metal2 40040 38752 40040 38752 0 cm_inst.cc_inst.out_notouch_\[130\]
rlabel metal2 17752 35728 17752 35728 0 cm_inst.cc_inst.out_notouch_\[131\]
rlabel metal2 36008 8736 36008 8736 0 cm_inst.cc_inst.out_notouch_\[132\]
rlabel metal2 25592 40488 25592 40488 0 cm_inst.cc_inst.out_notouch_\[133\]
rlabel metal2 39032 31304 39032 31304 0 cm_inst.cc_inst.out_notouch_\[134\]
rlabel metal2 19320 32088 19320 32088 0 cm_inst.cc_inst.out_notouch_\[135\]
rlabel metal2 40936 8316 40936 8316 0 cm_inst.cc_inst.out_notouch_\[136\]
rlabel metal2 28952 41104 28952 41104 0 cm_inst.cc_inst.out_notouch_\[137\]
rlabel metal2 39032 39088 39032 39088 0 cm_inst.cc_inst.out_notouch_\[138\]
rlabel metal2 14392 36568 14392 36568 0 cm_inst.cc_inst.out_notouch_\[139\]
rlabel metal2 20776 10864 20776 10864 0 cm_inst.cc_inst.out_notouch_\[13\]
rlabel metal2 35112 9072 35112 9072 0 cm_inst.cc_inst.out_notouch_\[140\]
rlabel metal2 24472 40656 24472 40656 0 cm_inst.cc_inst.out_notouch_\[141\]
rlabel metal2 37856 30968 37856 30968 0 cm_inst.cc_inst.out_notouch_\[142\]
rlabel metal2 18144 31752 18144 31752 0 cm_inst.cc_inst.out_notouch_\[143\]
rlabel metal2 38528 9240 38528 9240 0 cm_inst.cc_inst.out_notouch_\[144\]
rlabel metal2 26768 40488 26768 40488 0 cm_inst.cc_inst.out_notouch_\[145\]
rlabel metal3 36568 37912 36568 37912 0 cm_inst.cc_inst.out_notouch_\[146\]
rlabel metal2 14560 34888 14560 34888 0 cm_inst.cc_inst.out_notouch_\[147\]
rlabel metal2 32480 7672 32480 7672 0 cm_inst.cc_inst.out_notouch_\[148\]
rlabel metal2 22400 39704 22400 39704 0 cm_inst.cc_inst.out_notouch_\[149\]
rlabel metal2 29848 32256 29848 32256 0 cm_inst.cc_inst.out_notouch_\[14\]
rlabel metal2 35896 32088 35896 32088 0 cm_inst.cc_inst.out_notouch_\[150\]
rlabel metal2 14504 33376 14504 33376 0 cm_inst.cc_inst.out_notouch_\[151\]
rlabel metal2 39368 8512 39368 8512 0 cm_inst.cc_inst.out_notouch_\[152\]
rlabel metal2 27608 40712 27608 40712 0 cm_inst.cc_inst.out_notouch_\[153\]
rlabel metal2 37240 38472 37240 38472 0 cm_inst.cc_inst.out_notouch_\[154\]
rlabel metal2 14616 35280 14616 35280 0 cm_inst.cc_inst.out_notouch_\[155\]
rlabel metal2 33768 8344 33768 8344 0 cm_inst.cc_inst.out_notouch_\[156\]
rlabel metal2 23240 39872 23240 39872 0 cm_inst.cc_inst.out_notouch_\[157\]
rlabel metal2 36680 31304 36680 31304 0 cm_inst.cc_inst.out_notouch_\[158\]
rlabel metal2 16856 31752 16856 31752 0 cm_inst.cc_inst.out_notouch_\[159\]
rlabel metal2 28056 7168 28056 7168 0 cm_inst.cc_inst.out_notouch_\[15\]
rlabel metal2 45864 12656 45864 12656 0 cm_inst.cc_inst.out_notouch_\[160\]
rlabel metal2 32312 35784 32312 35784 0 cm_inst.cc_inst.out_notouch_\[161\]
rlabel metal3 45472 18424 45472 18424 0 cm_inst.cc_inst.out_notouch_\[162\]
rlabel metal2 18088 39788 18088 39788 0 cm_inst.cc_inst.out_notouch_\[163\]
rlabel metal2 43064 14924 43064 14924 0 cm_inst.cc_inst.out_notouch_\[164\]
rlabel metal3 33264 39816 33264 39816 0 cm_inst.cc_inst.out_notouch_\[165\]
rlabel metal2 44184 33600 44184 33600 0 cm_inst.cc_inst.out_notouch_\[166\]
rlabel metal2 20552 39088 20552 39088 0 cm_inst.cc_inst.out_notouch_\[167\]
rlabel metal2 42168 12264 42168 12264 0 cm_inst.cc_inst.out_notouch_\[168\]
rlabel metal2 31416 36176 31416 36176 0 cm_inst.cc_inst.out_notouch_\[169\]
rlabel metal2 29288 25480 29288 25480 0 cm_inst.cc_inst.out_notouch_\[16\]
rlabel metal2 44072 19712 44072 19712 0 cm_inst.cc_inst.out_notouch_\[170\]
rlabel metal3 16576 38808 16576 38808 0 cm_inst.cc_inst.out_notouch_\[171\]
rlabel metal2 45360 15064 45360 15064 0 cm_inst.cc_inst.out_notouch_\[172\]
rlabel metal2 31752 42000 31752 42000 0 cm_inst.cc_inst.out_notouch_\[173\]
rlabel metal2 43960 33544 43960 33544 0 cm_inst.cc_inst.out_notouch_\[174\]
rlabel metal2 17976 41664 17976 41664 0 cm_inst.cc_inst.out_notouch_\[175\]
rlabel metal2 39816 12824 39816 12824 0 cm_inst.cc_inst.out_notouch_\[176\]
rlabel metal2 28504 35728 28504 35728 0 cm_inst.cc_inst.out_notouch_\[177\]
rlabel metal2 41832 20496 41832 20496 0 cm_inst.cc_inst.out_notouch_\[178\]
rlabel metal2 14840 38640 14840 38640 0 cm_inst.cc_inst.out_notouch_\[179\]
rlabel metal2 20608 4424 20608 4424 0 cm_inst.cc_inst.out_notouch_\[17\]
rlabel metal2 39760 15400 39760 15400 0 cm_inst.cc_inst.out_notouch_\[180\]
rlabel metal2 29344 39032 29344 39032 0 cm_inst.cc_inst.out_notouch_\[181\]
rlabel metal2 40936 33208 40936 33208 0 cm_inst.cc_inst.out_notouch_\[182\]
rlabel metal3 15624 38696 15624 38696 0 cm_inst.cc_inst.out_notouch_\[183\]
rlabel metal2 40320 12376 40320 12376 0 cm_inst.cc_inst.out_notouch_\[184\]
rlabel metal2 29960 35392 29960 35392 0 cm_inst.cc_inst.out_notouch_\[185\]
rlabel metal2 42672 17864 42672 17864 0 cm_inst.cc_inst.out_notouch_\[186\]
rlabel metal2 12824 38696 12824 38696 0 cm_inst.cc_inst.out_notouch_\[187\]
rlabel metal2 40936 14532 40936 14532 0 cm_inst.cc_inst.out_notouch_\[188\]
rlabel metal2 31864 40768 31864 40768 0 cm_inst.cc_inst.out_notouch_\[189\]
rlabel metal2 25200 29624 25200 29624 0 cm_inst.cc_inst.out_notouch_\[18\]
rlabel metal2 41832 32872 41832 32872 0 cm_inst.cc_inst.out_notouch_\[190\]
rlabel metal2 18312 39536 18312 39536 0 cm_inst.cc_inst.out_notouch_\[191\]
rlabel metal2 23688 16408 23688 16408 0 cm_inst.cc_inst.out_notouch_\[192\]
rlabel metal2 22344 14504 22344 14504 0 cm_inst.cc_inst.out_notouch_\[193\]
rlabel metal2 24584 18816 24584 18816 0 cm_inst.cc_inst.out_notouch_\[194\]
rlabel metal2 12824 28896 12824 28896 0 cm_inst.cc_inst.out_notouch_\[195\]
rlabel metal2 23800 20496 23800 20496 0 cm_inst.cc_inst.out_notouch_\[196\]
rlabel metal2 19096 28224 19096 28224 0 cm_inst.cc_inst.out_notouch_\[197\]
rlabel metal2 19544 29736 19544 29736 0 cm_inst.cc_inst.out_notouch_\[198\]
rlabel metal2 17640 27552 17640 27552 0 cm_inst.cc_inst.out_notouch_\[199\]
rlabel metal2 23800 9688 23800 9688 0 cm_inst.cc_inst.out_notouch_\[19\]
rlabel metal2 17528 5152 17528 5152 0 cm_inst.cc_inst.out_notouch_\[1\]
rlabel metal2 21728 15400 21728 15400 0 cm_inst.cc_inst.out_notouch_\[200\]
rlabel metal2 21560 15876 21560 15876 0 cm_inst.cc_inst.out_notouch_\[201\]
rlabel metal2 23800 18032 23800 18032 0 cm_inst.cc_inst.out_notouch_\[202\]
rlabel metal2 12040 29848 12040 29848 0 cm_inst.cc_inst.out_notouch_\[203\]
rlabel metal2 23072 20216 23072 20216 0 cm_inst.cc_inst.out_notouch_\[204\]
rlabel metal2 19656 29400 19656 29400 0 cm_inst.cc_inst.out_notouch_\[205\]
rlabel metal2 18480 28728 18480 28728 0 cm_inst.cc_inst.out_notouch_\[206\]
rlabel metal3 17472 27608 17472 27608 0 cm_inst.cc_inst.out_notouch_\[207\]
rlabel metal3 21560 15512 21560 15512 0 cm_inst.cc_inst.out_notouch_\[208\]
rlabel metal2 19880 16072 19880 16072 0 cm_inst.cc_inst.out_notouch_\[209\]
rlabel metal2 24360 30520 24360 30520 0 cm_inst.cc_inst.out_notouch_\[20\]
rlabel metal3 18368 10472 18368 10472 0 cm_inst.cc_inst.out_notouch_\[21\]
rlabel metal2 26936 32088 26936 32088 0 cm_inst.cc_inst.out_notouch_\[22\]
rlabel metal2 25816 7784 25816 7784 0 cm_inst.cc_inst.out_notouch_\[23\]
rlabel metal2 30408 24136 30408 24136 0 cm_inst.cc_inst.out_notouch_\[24\]
rlabel metal2 19768 4424 19768 4424 0 cm_inst.cc_inst.out_notouch_\[25\]
rlabel metal3 25200 30184 25200 30184 0 cm_inst.cc_inst.out_notouch_\[26\]
rlabel metal2 24808 11256 24808 11256 0 cm_inst.cc_inst.out_notouch_\[27\]
rlabel metal2 26152 31248 26152 31248 0 cm_inst.cc_inst.out_notouch_\[28\]
rlabel metal2 19320 10248 19320 10248 0 cm_inst.cc_inst.out_notouch_\[29\]
rlabel metal3 28448 31080 28448 31080 0 cm_inst.cc_inst.out_notouch_\[2\]
rlabel metal2 28616 32984 28616 32984 0 cm_inst.cc_inst.out_notouch_\[30\]
rlabel metal2 26712 7784 26712 7784 0 cm_inst.cc_inst.out_notouch_\[31\]
rlabel metal2 32312 28672 32312 28672 0 cm_inst.cc_inst.out_notouch_\[32\]
rlabel metal2 18312 10864 18312 10864 0 cm_inst.cc_inst.out_notouch_\[33\]
rlabel metal2 24360 36344 24360 36344 0 cm_inst.cc_inst.out_notouch_\[34\]
rlabel metal2 24584 5544 24584 5544 0 cm_inst.cc_inst.out_notouch_\[35\]
rlabel metal2 26096 34888 26096 34888 0 cm_inst.cc_inst.out_notouch_\[36\]
rlabel metal2 19432 11368 19432 11368 0 cm_inst.cc_inst.out_notouch_\[37\]
rlabel metal2 24248 31752 24248 31752 0 cm_inst.cc_inst.out_notouch_\[38\]
rlabel metal2 25368 6384 25368 6384 0 cm_inst.cc_inst.out_notouch_\[39\]
rlabel metal2 27160 10528 27160 10528 0 cm_inst.cc_inst.out_notouch_\[3\]
rlabel metal2 31304 28896 31304 28896 0 cm_inst.cc_inst.out_notouch_\[40\]
rlabel metal2 17304 9912 17304 9912 0 cm_inst.cc_inst.out_notouch_\[41\]
rlabel metal2 23352 35000 23352 35000 0 cm_inst.cc_inst.out_notouch_\[42\]
rlabel metal2 23688 5208 23688 5208 0 cm_inst.cc_inst.out_notouch_\[43\]
rlabel metal2 24920 35560 24920 35560 0 cm_inst.cc_inst.out_notouch_\[44\]
rlabel metal2 18088 12040 18088 12040 0 cm_inst.cc_inst.out_notouch_\[45\]
rlabel metal2 23352 32424 23352 32424 0 cm_inst.cc_inst.out_notouch_\[46\]
rlabel metal2 23016 5936 23016 5936 0 cm_inst.cc_inst.out_notouch_\[47\]
rlabel metal3 28504 28616 28504 28616 0 cm_inst.cc_inst.out_notouch_\[48\]
rlabel metal2 15008 9688 15008 9688 0 cm_inst.cc_inst.out_notouch_\[49\]
rlabel metal3 28784 30184 28784 30184 0 cm_inst.cc_inst.out_notouch_\[4\]
rlabel metal2 21224 36064 21224 36064 0 cm_inst.cc_inst.out_notouch_\[50\]
rlabel metal2 22120 4760 22120 4760 0 cm_inst.cc_inst.out_notouch_\[51\]
rlabel metal2 22848 35000 22848 35000 0 cm_inst.cc_inst.out_notouch_\[52\]
rlabel metal2 15736 9128 15736 9128 0 cm_inst.cc_inst.out_notouch_\[53\]
rlabel metal2 21336 32088 21336 32088 0 cm_inst.cc_inst.out_notouch_\[54\]
rlabel metal2 21000 6552 21000 6552 0 cm_inst.cc_inst.out_notouch_\[55\]
rlabel metal2 30184 28896 30184 28896 0 cm_inst.cc_inst.out_notouch_\[56\]
rlabel metal2 15960 9072 15960 9072 0 cm_inst.cc_inst.out_notouch_\[57\]
rlabel metal2 22008 36400 22008 36400 0 cm_inst.cc_inst.out_notouch_\[58\]
rlabel metal3 21728 5880 21728 5880 0 cm_inst.cc_inst.out_notouch_\[59\]
rlabel metal2 21840 10024 21840 10024 0 cm_inst.cc_inst.out_notouch_\[5\]
rlabel metal2 23800 36400 23800 36400 0 cm_inst.cc_inst.out_notouch_\[60\]
rlabel metal2 15736 11312 15736 11312 0 cm_inst.cc_inst.out_notouch_\[61\]
rlabel metal2 21672 31360 21672 31360 0 cm_inst.cc_inst.out_notouch_\[62\]
rlabel metal2 21952 6664 21952 6664 0 cm_inst.cc_inst.out_notouch_\[63\]
rlabel metal2 44968 30128 44968 30128 0 cm_inst.cc_inst.out_notouch_\[64\]
rlabel metal2 28280 11424 28280 11424 0 cm_inst.cc_inst.out_notouch_\[65\]
rlabel metal3 44184 37128 44184 37128 0 cm_inst.cc_inst.out_notouch_\[66\]
rlabel metal2 32424 12264 32424 12264 0 cm_inst.cc_inst.out_notouch_\[67\]
rlabel metal2 36344 13272 36344 13272 0 cm_inst.cc_inst.out_notouch_\[68\]
rlabel metal3 29008 14504 29008 14504 0 cm_inst.cc_inst.out_notouch_\[69\]
rlabel metal2 30744 31696 30744 31696 0 cm_inst.cc_inst.out_notouch_\[6\]
rlabel metal2 38584 35952 38584 35952 0 cm_inst.cc_inst.out_notouch_\[70\]
rlabel metal2 38136 20272 38136 20272 0 cm_inst.cc_inst.out_notouch_\[71\]
rlabel metal2 43960 28952 43960 28952 0 cm_inst.cc_inst.out_notouch_\[72\]
rlabel metal2 27496 12432 27496 12432 0 cm_inst.cc_inst.out_notouch_\[73\]
rlabel metal2 43176 37688 43176 37688 0 cm_inst.cc_inst.out_notouch_\[74\]
rlabel metal2 31528 12432 31528 12432 0 cm_inst.cc_inst.out_notouch_\[75\]
rlabel metal2 35616 12936 35616 12936 0 cm_inst.cc_inst.out_notouch_\[76\]
rlabel metal2 27664 14504 27664 14504 0 cm_inst.cc_inst.out_notouch_\[77\]
rlabel metal2 37800 35168 37800 35168 0 cm_inst.cc_inst.out_notouch_\[78\]
rlabel metal3 36848 18984 36848 18984 0 cm_inst.cc_inst.out_notouch_\[79\]
rlabel metal2 28840 6608 28840 6608 0 cm_inst.cc_inst.out_notouch_\[7\]
rlabel metal2 41944 29736 41944 29736 0 cm_inst.cc_inst.out_notouch_\[80\]
rlabel metal2 24584 11424 24584 11424 0 cm_inst.cc_inst.out_notouch_\[81\]
rlabel metal2 40656 37352 40656 37352 0 cm_inst.cc_inst.out_notouch_\[82\]
rlabel metal2 29288 11256 29288 11256 0 cm_inst.cc_inst.out_notouch_\[83\]
rlabel metal2 33320 11256 33320 11256 0 cm_inst.cc_inst.out_notouch_\[84\]
rlabel metal2 25368 15288 25368 15288 0 cm_inst.cc_inst.out_notouch_\[85\]
rlabel metal2 35560 36232 35560 36232 0 cm_inst.cc_inst.out_notouch_\[86\]
rlabel metal2 34888 19992 34888 19992 0 cm_inst.cc_inst.out_notouch_\[87\]
rlabel metal2 42728 29064 42728 29064 0 cm_inst.cc_inst.out_notouch_\[88\]
rlabel metal2 26152 11816 26152 11816 0 cm_inst.cc_inst.out_notouch_\[89\]
rlabel metal2 31304 25928 31304 25928 0 cm_inst.cc_inst.out_notouch_\[8\]
rlabel metal2 41720 38080 41720 38080 0 cm_inst.cc_inst.out_notouch_\[90\]
rlabel metal2 30072 12656 30072 12656 0 cm_inst.cc_inst.out_notouch_\[91\]
rlabel metal2 33992 12208 33992 12208 0 cm_inst.cc_inst.out_notouch_\[92\]
rlabel metal2 26208 16632 26208 16632 0 cm_inst.cc_inst.out_notouch_\[93\]
rlabel metal2 36456 36008 36456 36008 0 cm_inst.cc_inst.out_notouch_\[94\]
rlabel metal2 36008 19152 36008 19152 0 cm_inst.cc_inst.out_notouch_\[95\]
rlabel metal2 37240 24360 37240 24360 0 cm_inst.cc_inst.out_notouch_\[96\]
rlabel metal2 44072 24640 44072 24640 0 cm_inst.cc_inst.out_notouch_\[97\]
rlabel metal2 43456 25480 43456 25480 0 cm_inst.cc_inst.out_notouch_\[98\]
rlabel metal3 33936 20776 33936 20776 0 cm_inst.cc_inst.out_notouch_\[99\]
rlabel metal2 18536 4592 18536 4592 0 cm_inst.cc_inst.out_notouch_\[9\]
rlabel metal2 21392 23912 21392 23912 0 cm_inst.page\[0\]
rlabel metal2 25480 14336 25480 14336 0 cm_inst.page\[1\]
rlabel metal2 16968 26208 16968 26208 0 cm_inst.page\[2\]
rlabel metal2 25032 22064 25032 22064 0 cm_inst.page\[3\]
rlabel metal2 18648 24080 18648 24080 0 cm_inst.page\[4\]
rlabel metal2 21896 23968 21896 23968 0 cm_inst.page\[5\]
rlabel metal2 1736 34552 1736 34552 0 in[0]
rlabel metal2 1848 17696 1848 17696 0 in[1]
rlabel metal2 1736 17920 1736 17920 0 in[2]
rlabel metal2 2408 17192 2408 17192 0 in[3]
rlabel metal3 4900 19992 4900 19992 0 in[4]
rlabel metal2 1736 18928 1736 18928 0 in[5]
rlabel metal2 1960 19656 1960 19656 0 in[6]
rlabel metal2 3528 19376 3528 19376 0 in[7]
rlabel metal2 2072 35560 2072 35560 0 net1
rlabel metal2 4312 24360 4312 24360 0 net10
rlabel metal2 14616 29400 14616 29400 0 net100
rlabel metal2 13608 28056 13608 28056 0 net101
rlabel metal2 14896 27160 14896 27160 0 net102
rlabel metal2 13552 37464 13552 37464 0 net103
rlabel metal2 17472 40936 17472 40936 0 net104
rlabel metal2 22120 36400 22120 36400 0 net105
rlabel metal2 25144 36792 25144 36792 0 net106
rlabel metal2 25592 42336 25592 42336 0 net107
rlabel metal3 24080 42728 24080 42728 0 net108
rlabel metal3 13888 37464 13888 37464 0 net109
rlabel metal2 6664 25200 6664 25200 0 net11
rlabel metal2 15064 37128 15064 37128 0 net110
rlabel metal2 29008 26152 29008 26152 0 net111
rlabel metal3 35280 30072 35280 30072 0 net112
rlabel metal2 28392 25928 28392 25928 0 net113
rlabel metal2 45416 29456 45416 29456 0 net114
rlabel metal2 45304 30968 45304 30968 0 net115
rlabel metal2 40040 27776 40040 27776 0 net116
rlabel metal2 45864 31640 45864 31640 0 net117
rlabel metal3 28000 25256 28000 25256 0 net118
rlabel metal3 29400 41944 29400 41944 0 net119
rlabel metal2 4312 23016 4312 23016 0 net12
rlabel metal2 30744 40096 30744 40096 0 net120
rlabel metal2 38920 37184 38920 37184 0 net121
rlabel metal2 39144 36624 39144 36624 0 net122
rlabel metal2 43120 36456 43120 36456 0 net123
rlabel metal3 44548 34104 44548 34104 0 net124
rlabel metal2 34776 35280 34776 35280 0 net125
rlabel metal3 33880 28056 33880 28056 0 net126
rlabel metal2 17752 29568 17752 29568 0 net127
rlabel metal2 12320 21784 12320 21784 0 net128
rlabel metal2 15064 11648 15064 11648 0 net129
rlabel metal2 5096 23072 5096 23072 0 net13
rlabel metal2 15848 13384 15848 13384 0 net130
rlabel metal2 13552 8344 13552 8344 0 net131
rlabel metal2 12600 11200 12600 11200 0 net132
rlabel metal2 19544 3752 19544 3752 0 net133
rlabel metal2 20216 9240 20216 9240 0 net134
rlabel metal2 24920 8288 24920 8288 0 net135
rlabel metal2 24696 7392 24696 7392 0 net136
rlabel metal3 22960 9016 22960 9016 0 net137
rlabel metal2 26040 11424 26040 11424 0 net138
rlabel metal2 24136 9576 24136 9576 0 net139
rlabel metal2 4312 21448 4312 21448 0 net14
rlabel metal2 12936 11480 12936 11480 0 net140
rlabel metal2 12264 16016 12264 16016 0 net141
rlabel metal2 25480 16240 25480 16240 0 net142
rlabel metal2 12712 13832 12712 13832 0 net143
rlabel metal2 31864 8288 31864 8288 0 net144
rlabel metal3 35112 7448 35112 7448 0 net145
rlabel metal2 30632 12040 30632 12040 0 net146
rlabel metal3 32704 11480 32704 11480 0 net147
rlabel metal2 30184 11704 30184 11704 0 net148
rlabel metal3 42112 12152 42112 12152 0 net149
rlabel metal2 4312 28336 4312 28336 0 net15
rlabel metal2 30520 14112 30520 14112 0 net150
rlabel metal3 29288 16184 29288 16184 0 net151
rlabel metal2 34160 17640 34160 17640 0 net152
rlabel metal2 31304 21896 31304 21896 0 net153
rlabel metal2 34440 21560 34440 21560 0 net154
rlabel metal2 36568 17360 36568 17360 0 net155
rlabel metal2 39144 18816 39144 18816 0 net156
rlabel metal2 42056 17808 42056 17808 0 net157
rlabel metal2 39032 23464 39032 23464 0 net158
rlabel metal2 42504 21952 42504 21952 0 net159
rlabel metal2 9576 27496 9576 27496 0 net16
rlabel metal2 44968 24472 44968 24472 0 net160
rlabel metal2 39704 17416 39704 17416 0 net161
rlabel metal2 29624 14112 29624 14112 0 net162
rlabel metal2 13944 13048 13944 13048 0 net163
rlabel metal2 14952 29960 14952 29960 0 net164
rlabel metal2 15064 29792 15064 29792 0 net165
rlabel metal2 13944 29008 13944 29008 0 net166
rlabel metal2 23464 31360 23464 31360 0 net167
rlabel metal3 25928 33096 25928 33096 0 net168
rlabel metal3 23856 33320 23856 33320 0 net169
rlabel metal3 28560 39480 28560 39480 0 net17
rlabel metal2 22568 31920 22568 31920 0 net170
rlabel metal2 14168 28840 14168 28840 0 net171
rlabel metal2 10808 36288 10808 36288 0 net172
rlabel metal3 15008 39592 15008 39592 0 net173
rlabel metal2 21896 35952 21896 35952 0 net174
rlabel metal2 18872 37968 18872 37968 0 net175
rlabel metal3 19712 38136 19712 38136 0 net176
rlabel metal2 23352 42672 23352 42672 0 net177
rlabel metal3 26152 41944 26152 41944 0 net178
rlabel metal2 21672 39928 21672 39928 0 net179
rlabel metal2 35224 20328 35224 20328 0 net18
rlabel metal2 21336 40096 21336 40096 0 net180
rlabel metal2 14616 31080 14616 31080 0 net181
rlabel metal2 31864 29008 31864 29008 0 net182
rlabel metal3 30856 26600 30856 26600 0 net183
rlabel metal2 32312 25088 32312 25088 0 net184
rlabel metal2 39256 26992 39256 26992 0 net185
rlabel metal2 44856 28392 44856 28392 0 net186
rlabel metal2 44744 27160 44744 27160 0 net187
rlabel metal2 44856 30184 44856 30184 0 net188
rlabel metal2 44968 31472 44968 31472 0 net189
rlabel metal2 42280 16520 42280 16520 0 net19
rlabel metal3 29456 42728 29456 42728 0 net190
rlabel metal2 32536 38864 32536 38864 0 net191
rlabel metal2 32648 37128 32648 37128 0 net192
rlabel metal2 39592 37072 39592 37072 0 net193
rlabel metal3 40768 36232 40768 36232 0 net194
rlabel metal2 44856 36064 44856 36064 0 net195
rlabel metal2 37800 38920 37800 38920 0 net196
rlabel metal3 39704 38752 39704 38752 0 net197
rlabel metal2 27944 26768 27944 26768 0 net198
rlabel metal2 16912 30856 16912 30856 0 net199
rlabel metal2 14056 19152 14056 19152 0 net2
rlabel metal3 39144 34664 39144 34664 0 net20
rlabel metal3 14000 12936 14000 12936 0 net200
rlabel metal2 14840 11368 14840 11368 0 net201
rlabel metal2 13496 10696 13496 10696 0 net202
rlabel metal3 12936 11368 12936 11368 0 net203
rlabel metal2 14504 12880 14504 12880 0 net204
rlabel metal2 19880 6496 19880 6496 0 net205
rlabel metal2 19096 6328 19096 6328 0 net206
rlabel metal2 25480 6776 25480 6776 0 net207
rlabel metal2 24920 6720 24920 6720 0 net208
rlabel metal3 22288 8008 22288 8008 0 net209
rlabel metal2 42728 34664 42728 34664 0 net21
rlabel metal3 20776 9800 20776 9800 0 net210
rlabel metal3 20216 15176 20216 15176 0 net211
rlabel metal2 24248 11872 24248 11872 0 net212
rlabel metal2 26264 9856 26264 9856 0 net213
rlabel metal2 22680 11256 22680 11256 0 net214
rlabel metal3 21952 14952 21952 14952 0 net215
rlabel metal2 20272 14280 20272 14280 0 net216
rlabel metal2 14952 12936 14952 12936 0 net217
rlabel metal2 21672 16296 21672 16296 0 net218
rlabel metal2 17528 17584 17528 17584 0 net219
rlabel metal2 36848 21784 36848 21784 0 net22
rlabel metal2 23240 18424 23240 18424 0 net220
rlabel metal3 25368 19880 25368 19880 0 net221
rlabel metal2 10024 16800 10024 16800 0 net222
rlabel metal2 9688 16072 9688 16072 0 net223
rlabel metal2 29512 7840 29512 7840 0 net224
rlabel metal2 35672 7392 35672 7392 0 net225
rlabel metal2 32760 13272 32760 13272 0 net226
rlabel metal3 34496 13720 34496 13720 0 net227
rlabel metal2 29568 6664 29568 6664 0 net228
rlabel metal2 38696 12096 38696 12096 0 net229
rlabel metal2 7280 24920 7280 24920 0 net23
rlabel metal2 42840 12096 42840 12096 0 net230
rlabel metal2 27832 14056 27832 14056 0 net231
rlabel metal2 31080 16576 31080 16576 0 net232
rlabel metal2 34440 16072 34440 16072 0 net233
rlabel metal2 31192 22064 31192 22064 0 net234
rlabel metal2 34664 21168 34664 21168 0 net235
rlabel metal2 28280 21672 28280 21672 0 net236
rlabel metal2 41160 14112 41160 14112 0 net237
rlabel metal2 38976 19880 38976 19880 0 net238
rlabel metal3 41216 16968 41216 16968 0 net239
rlabel metal2 14392 38864 14392 38864 0 net24
rlabel metal2 42504 19488 42504 19488 0 net240
rlabel metal2 38584 23464 38584 23464 0 net241
rlabel metal2 42728 21224 42728 21224 0 net242
rlabel metal2 38136 21840 38136 21840 0 net243
rlabel metal2 29736 18200 29736 18200 0 net244
rlabel metal2 29624 17080 29624 17080 0 net245
rlabel metal2 9688 17864 9688 17864 0 net246
rlabel metal2 13496 31192 13496 31192 0 net247
rlabel metal2 12656 31864 12656 31864 0 net248
rlabel metal2 13496 30128 13496 30128 0 net249
rlabel metal3 24752 39704 24752 39704 0 net25
rlabel metal2 23128 30520 23128 30520 0 net250
rlabel metal2 25480 31416 25480 31416 0 net251
rlabel metal2 24416 32536 24416 32536 0 net252
rlabel metal2 21448 32872 21448 32872 0 net253
rlabel metal2 21224 29680 21224 29680 0 net254
rlabel metal2 14112 30184 14112 30184 0 net255
rlabel metal2 16184 39928 16184 39928 0 net256
rlabel via2 12600 38920 12600 38920 0 net257
rlabel metal2 10136 36400 10136 36400 0 net258
rlabel metal2 12824 41048 12824 41048 0 net259
rlabel metal2 35672 12320 35672 12320 0 net26
rlabel metal2 23464 35672 23464 35672 0 net260
rlabel metal2 26544 36344 26544 36344 0 net261
rlabel metal3 23296 36456 23296 36456 0 net262
rlabel metal3 23072 42504 23072 42504 0 net263
rlabel metal2 22904 43120 22904 43120 0 net264
rlabel metal2 21224 38920 21224 38920 0 net265
rlabel metal3 20580 38920 20580 38920 0 net266
rlabel metal3 12768 31640 12768 31640 0 net267
rlabel metal2 30072 25088 30072 25088 0 net268
rlabel metal2 28616 29064 28616 29064 0 net269
rlabel metal2 34776 17864 34776 17864 0 net27
rlabel metal2 29848 27888 29848 27888 0 net270
rlabel metal2 29232 31192 29232 31192 0 net271
rlabel metal3 32536 33320 32536 33320 0 net272
rlabel metal2 33544 29064 33544 29064 0 net273
rlabel metal3 31920 29960 31920 29960 0 net274
rlabel metal2 38528 28616 38528 28616 0 net275
rlabel metal3 44632 26936 44632 26936 0 net276
rlabel metal2 44184 28448 44184 28448 0 net277
rlabel metal2 45640 30744 45640 30744 0 net278
rlabel metal3 43764 28280 43764 28280 0 net279
rlabel metal2 32200 18928 32200 18928 0 net28
rlabel metal2 38696 28840 38696 28840 0 net280
rlabel metal2 27832 40936 27832 40936 0 net281
rlabel metal2 28280 40040 28280 40040 0 net282
rlabel metal2 30184 35056 30184 35056 0 net283
rlabel metal2 28056 39424 28056 39424 0 net284
rlabel metal2 43288 37184 43288 37184 0 net285
rlabel metal3 40712 37240 40712 37240 0 net286
rlabel metal3 38780 33992 38780 33992 0 net287
rlabel metal2 41104 35784 41104 35784 0 net288
rlabel metal2 40488 35952 40488 35952 0 net289
rlabel metal2 33208 23072 33208 23072 0 net29
rlabel metal2 28504 42560 28504 42560 0 net290
rlabel metal2 29400 28840 29400 28840 0 net291
rlabel metal2 12320 31192 12320 31192 0 net292
rlabel metal2 10472 26600 10472 26600 0 net293
rlabel metal2 4984 6888 4984 6888 0 net294
rlabel metal2 4816 12376 4816 12376 0 net295
rlabel metal2 12600 14616 12600 14616 0 net296
rlabel metal2 8344 14952 8344 14952 0 net297
rlabel metal2 4872 14952 4872 14952 0 net298
rlabel metal2 5656 17864 5656 17864 0 net299
rlabel metal3 12544 16968 12544 16968 0 net3
rlabel metal2 38696 14784 38696 14784 0 net30
rlabel metal2 4760 20356 4760 20356 0 net300
rlabel metal3 5880 20552 5880 20552 0 net301
rlabel metal2 5992 20496 5992 20496 0 net302
rlabel metal2 13496 21280 13496 21280 0 net303
rlabel metal2 7560 21448 7560 21448 0 net304
rlabel metal2 4872 22568 4872 22568 0 net305
rlabel metal2 4760 28000 4760 28000 0 net306
rlabel metal2 7000 26152 7000 26152 0 net307
rlabel metal2 4872 30408 4872 30408 0 net308
rlabel metal2 5432 37520 5432 37520 0 net309
rlabel metal2 40264 23128 40264 23128 0 net31
rlabel metal3 4760 34664 4760 34664 0 net310
rlabel metal2 9688 31780 9688 31780 0 net311
rlabel metal2 5992 30716 5992 30716 0 net312
rlabel metal2 3528 35168 3528 35168 0 net313
rlabel metal2 7896 23632 7896 23632 0 net314
rlabel metal2 7896 27720 7896 27720 0 net315
rlabel metal3 1246 42392 1246 42392 0 net316
rlabel metal3 1246 4760 1246 4760 0 net317
rlabel metal2 46200 42448 46200 42448 0 net318
rlabel metal3 854 43064 854 43064 0 net319
rlabel metal2 40376 19768 40376 19768 0 net32
rlabel metal2 40824 29624 40824 29624 0 net33
rlabel metal2 44968 35056 44968 35056 0 net34
rlabel metal2 41496 29792 41496 29792 0 net35
rlabel metal3 42056 29400 42056 29400 0 net36
rlabel metal2 19096 40320 19096 40320 0 net37
rlabel metal2 22456 10080 22456 10080 0 net38
rlabel metal3 14812 8904 14812 8904 0 net39
rlabel metal2 11592 17472 11592 17472 0 net4
rlabel metal2 14504 22232 14504 22232 0 net40
rlabel metal2 13832 21840 13832 21840 0 net41
rlabel metal2 35168 15960 35168 15960 0 net42
rlabel metal2 34664 16856 34664 16856 0 net43
rlabel metal2 41608 11200 41608 11200 0 net44
rlabel metal2 37016 19992 37016 19992 0 net45
rlabel metal2 33992 23520 33992 23520 0 net46
rlabel metal3 40012 18536 40012 18536 0 net47
rlabel metal2 39928 19600 39928 19600 0 net48
rlabel metal3 39592 23800 39592 23800 0 net49
rlabel metal2 12040 20832 12040 20832 0 net5
rlabel metal2 38920 23856 38920 23856 0 net50
rlabel metal2 33488 20104 33488 20104 0 net51
rlabel metal2 14168 23184 14168 23184 0 net52
rlabel metal2 15176 40432 15176 40432 0 net53
rlabel metal2 15960 40376 15960 40376 0 net54
rlabel metal2 22344 37408 22344 37408 0 net55
rlabel metal2 22512 38920 22512 38920 0 net56
rlabel metal2 22232 39088 22232 39088 0 net57
rlabel metal2 12824 33152 12824 33152 0 net58
rlabel metal2 45640 28784 45640 28784 0 net59
rlabel metal2 6776 18816 6776 18816 0 net6
rlabel metal2 42504 29848 42504 29848 0 net60
rlabel metal2 41608 31528 41608 31528 0 net61
rlabel metal2 35896 38724 35896 38724 0 net62
rlabel metal2 30520 43344 30520 43344 0 net63
rlabel metal2 39480 37240 39480 37240 0 net64
rlabel metal2 44856 34328 44856 34328 0 net65
rlabel metal3 45192 34720 45192 34720 0 net66
rlabel metal2 31024 43512 31024 43512 0 net67
rlabel metal2 32256 23912 32256 23912 0 net68
rlabel metal2 16968 34216 16968 34216 0 net69
rlabel metal2 3192 19768 3192 19768 0 net7
rlabel metal2 16184 23352 16184 23352 0 net70
rlabel metal3 14672 8232 14672 8232 0 net71
rlabel metal2 13496 12208 13496 12208 0 net72
rlabel metal2 23520 7336 23520 7336 0 net73
rlabel metal2 23520 4312 23520 4312 0 net74
rlabel metal3 22176 7448 22176 7448 0 net75
rlabel metal2 21336 7896 21336 7896 0 net76
rlabel metal2 24024 10248 24024 10248 0 net77
rlabel metal2 12376 12208 12376 12208 0 net78
rlabel metal2 26040 16352 26040 16352 0 net79
rlabel metal2 13496 19824 13496 19824 0 net8
rlabel metal2 11256 20916 11256 20916 0 net80
rlabel metal2 11872 22120 11872 22120 0 net81
rlabel metal2 32088 12488 32088 12488 0 net82
rlabel metal3 31136 11368 31136 11368 0 net83
rlabel metal2 33656 10360 33656 10360 0 net84
rlabel metal2 31192 9856 31192 9856 0 net85
rlabel metal2 38024 13160 38024 13160 0 net86
rlabel metal2 37856 11368 37856 11368 0 net87
rlabel metal2 32312 14000 32312 14000 0 net88
rlabel metal3 30408 22456 30408 22456 0 net89
rlabel metal2 4312 25536 4312 25536 0 net9
rlabel metal2 35560 21896 35560 21896 0 net90
rlabel via2 35000 17640 35000 17640 0 net91
rlabel metal2 38864 18536 38864 18536 0 net92
rlabel metal2 42728 14000 42728 14000 0 net93
rlabel metal3 42672 23800 42672 23800 0 net94
rlabel metal2 45752 23520 45752 23520 0 net95
rlabel metal2 45976 24192 45976 24192 0 net96
rlabel metal2 29400 19488 29400 19488 0 net97
rlabel metal2 29064 22624 29064 22624 0 net98
rlabel metal2 12264 22456 12264 22456 0 net99
rlabel metal2 1960 25984 1960 25984 0 out[0]
rlabel metal2 2856 24864 2856 24864 0 out[1]
rlabel metal3 3640 25088 3640 25088 0 out[2]
rlabel metal2 2072 23352 2072 23352 0 out[3]
rlabel metal3 6664 23632 6664 23632 0 out[4]
rlabel metal2 2744 21896 2744 21896 0 out[5]
rlabel metal3 1358 27608 1358 27608 0 out[6]
rlabel metal3 1358 26936 1358 26936 0 out[7]
rlabel metal2 11032 24696 11032 24696 0 ro_inst.counter\[0\]
rlabel metal3 10360 11592 10360 11592 0 ro_inst.counter\[10\]
rlabel metal2 11480 11032 11480 11032 0 ro_inst.counter\[11\]
rlabel metal2 9912 9016 9912 9016 0 ro_inst.counter\[12\]
rlabel metal2 5992 10136 5992 10136 0 ro_inst.counter\[13\]
rlabel metal2 2968 9464 2968 9464 0 ro_inst.counter\[14\]
rlabel metal2 5880 6496 5880 6496 0 ro_inst.counter\[15\]
rlabel metal3 4872 9800 4872 9800 0 ro_inst.counter\[16\]
rlabel metal2 3752 11704 3752 11704 0 ro_inst.counter\[17\]
rlabel metal2 5320 11200 5320 11200 0 ro_inst.counter\[18\]
rlabel metal2 5264 12376 5264 12376 0 ro_inst.counter\[19\]
rlabel metal2 6216 25928 6216 25928 0 ro_inst.counter\[1\]
rlabel metal3 4536 13944 4536 13944 0 ro_inst.counter\[20\]
rlabel metal3 6440 17528 6440 17528 0 ro_inst.counter\[21\]
rlabel metal2 5320 18088 5320 18088 0 ro_inst.counter\[22\]
rlabel metal2 5320 28112 5320 28112 0 ro_inst.counter\[23\]
rlabel metal2 5432 29848 5432 29848 0 ro_inst.counter\[24\]
rlabel metal2 5544 31416 5544 31416 0 ro_inst.counter\[25\]
rlabel metal3 4648 32760 4648 32760 0 ro_inst.counter\[26\]
rlabel metal2 4312 33656 4312 33656 0 ro_inst.counter\[27\]
rlabel metal3 4256 35000 4256 35000 0 ro_inst.counter\[28\]
rlabel metal2 4984 34272 4984 34272 0 ro_inst.counter\[29\]
rlabel metal2 8008 23856 8008 23856 0 ro_inst.counter\[2\]
rlabel metal2 7560 36120 7560 36120 0 ro_inst.counter\[30\]
rlabel metal2 7896 35336 7896 35336 0 ro_inst.counter\[31\]
rlabel metal2 9408 34104 9408 34104 0 ro_inst.counter\[32\]
rlabel metal2 8680 32872 8680 32872 0 ro_inst.counter\[33\]
rlabel metal2 8344 31304 8344 31304 0 ro_inst.counter\[34\]
rlabel metal2 6216 23464 6216 23464 0 ro_inst.counter\[3\]
rlabel metal2 5656 21840 5656 21840 0 ro_inst.counter\[4\]
rlabel metal2 6272 20440 6272 20440 0 ro_inst.counter\[5\]
rlabel metal2 5096 17976 5096 17976 0 ro_inst.counter\[6\]
rlabel metal2 6104 16520 6104 16520 0 ro_inst.counter\[7\]
rlabel metal2 7336 14896 7336 14896 0 ro_inst.counter\[8\]
rlabel metal2 8680 13272 8680 13272 0 ro_inst.counter\[9\]
rlabel metal2 2744 25984 2744 25984 0 ro_inst.counter_n\[0\]
rlabel metal2 8008 11648 8008 11648 0 ro_inst.counter_n\[10\]
rlabel metal2 9744 10584 9744 10584 0 ro_inst.counter_n\[11\]
rlabel metal2 10024 9912 10024 9912 0 ro_inst.counter_n\[12\]
rlabel metal2 6104 10304 6104 10304 0 ro_inst.counter_n\[13\]
rlabel metal2 2072 5880 2072 5880 0 ro_inst.counter_n\[14\]
rlabel metal2 2072 7336 2072 7336 0 ro_inst.counter_n\[15\]
rlabel metal2 4088 11872 4088 11872 0 ro_inst.counter_n\[16\]
rlabel metal2 3584 11368 3584 11368 0 ro_inst.counter_n\[17\]
rlabel metal2 1848 12432 1848 12432 0 ro_inst.counter_n\[18\]
rlabel metal2 2184 12824 2184 12824 0 ro_inst.counter_n\[19\]
rlabel metal3 3920 26936 3920 26936 0 ro_inst.counter_n\[1\]
rlabel metal3 4536 16296 4536 16296 0 ro_inst.counter_n\[20\]
rlabel metal3 4816 17640 4816 17640 0 ro_inst.counter_n\[21\]
rlabel metal2 4984 18872 4984 18872 0 ro_inst.counter_n\[22\]
rlabel metal2 2296 28224 2296 28224 0 ro_inst.counter_n\[23\]
rlabel via2 2296 30184 2296 30184 0 ro_inst.counter_n\[24\]
rlabel metal2 2520 31248 2520 31248 0 ro_inst.counter_n\[25\]
rlabel metal2 2184 32536 2184 32536 0 ro_inst.counter_n\[26\]
rlabel metal2 2184 36456 2184 36456 0 ro_inst.counter_n\[27\]
rlabel metal2 2744 36176 2744 36176 0 ro_inst.counter_n\[28\]
rlabel metal2 3864 35504 3864 35504 0 ro_inst.counter_n\[29\]
rlabel metal2 1960 23800 1960 23800 0 ro_inst.counter_n\[2\]
rlabel metal2 5544 35560 5544 35560 0 ro_inst.counter_n\[30\]
rlabel metal2 6216 35168 6216 35168 0 ro_inst.counter_n\[31\]
rlabel metal2 6664 33600 6664 33600 0 ro_inst.counter_n\[32\]
rlabel metal2 7000 32536 7000 32536 0 ro_inst.counter_n\[33\]
rlabel metal3 7840 31192 7840 31192 0 ro_inst.counter_n\[34\]
rlabel metal2 8568 23352 8568 23352 0 ro_inst.counter_n\[3\]
rlabel metal2 2408 18928 2408 18928 0 ro_inst.counter_n\[4\]
rlabel metal2 2968 19208 2968 19208 0 ro_inst.counter_n\[5\]
rlabel metal2 4984 18144 4984 18144 0 ro_inst.counter_n\[6\]
rlabel metal2 5992 15568 5992 15568 0 ro_inst.counter_n\[7\]
rlabel metal2 5656 14000 5656 14000 0 ro_inst.counter_n\[8\]
rlabel metal2 7336 12040 7336 12040 0 ro_inst.counter_n\[9\]
rlabel metal2 10192 26376 10192 26376 0 ro_inst.enable
rlabel metal2 10024 27664 10024 27664 0 ro_inst.ring\[0\]
rlabel metal2 11536 27048 11536 27048 0 ro_inst.ring\[1\]
rlabel metal2 11536 27272 11536 27272 0 ro_inst.ring\[2\]
rlabel metal2 8120 26544 8120 26544 0 ro_inst.running
rlabel metal2 8680 26880 8680 26880 0 ro_inst.saved_signal
rlabel metal3 8008 26264 8008 26264 0 ro_inst.signal
rlabel metal2 7000 27832 7000 27832 0 ro_inst.slow_clk_n
rlabel metal2 10192 23128 10192 23128 0 ro_sel\[0\]
rlabel metal2 11144 23464 11144 23464 0 ro_sel\[1\]
rlabel metal2 10528 20888 10528 20888 0 ro_sel\[2\]
<< properties >>
string FIXED_BBOX 0 0 48000 48000
<< end >>
