magic
tech gf180mcuD
magscale 1 5
timestamp 1702441481
<< obsm1 >>
rect 672 1415 19400 18454
<< metal2 >>
rect 5376 19600 5432 20000
rect 5712 19600 5768 20000
rect 6048 19600 6104 20000
rect 6384 19600 6440 20000
rect 6720 19600 6776 20000
rect 7056 19600 7112 20000
rect 7392 19600 7448 20000
rect 7728 19600 7784 20000
rect 8064 19600 8120 20000
rect 8400 19600 8456 20000
rect 8736 19600 8792 20000
rect 9072 19600 9128 20000
rect 9408 19600 9464 20000
rect 9744 19600 9800 20000
rect 10080 19600 10136 20000
rect 10416 19600 10472 20000
rect 10752 19600 10808 20000
rect 11088 19600 11144 20000
rect 11424 19600 11480 20000
rect 11760 19600 11816 20000
rect 12096 19600 12152 20000
rect 12432 19600 12488 20000
rect 12768 19600 12824 20000
rect 13104 19600 13160 20000
rect 13440 19600 13496 20000
rect 6048 0 6104 400
rect 6384 0 6440 400
rect 6720 0 6776 400
rect 7056 0 7112 400
rect 7392 0 7448 400
rect 7728 0 7784 400
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 9744 0 9800 400
rect 10080 0 10136 400
rect 10416 0 10472 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 11424 0 11480 400
rect 11760 0 11816 400
rect 12096 0 12152 400
rect 12432 0 12488 400
rect 12768 0 12824 400
rect 13104 0 13160 400
rect 13440 0 13496 400
rect 13776 0 13832 400
rect 14112 0 14168 400
rect 14448 0 14504 400
rect 14784 0 14840 400
rect 15120 0 15176 400
<< obsm2 >>
rect 854 19570 5346 19600
rect 5462 19570 5682 19600
rect 5798 19570 6018 19600
rect 6134 19570 6354 19600
rect 6470 19570 6690 19600
rect 6806 19570 7026 19600
rect 7142 19570 7362 19600
rect 7478 19570 7698 19600
rect 7814 19570 8034 19600
rect 8150 19570 8370 19600
rect 8486 19570 8706 19600
rect 8822 19570 9042 19600
rect 9158 19570 9378 19600
rect 9494 19570 9714 19600
rect 9830 19570 10050 19600
rect 10166 19570 10386 19600
rect 10502 19570 10722 19600
rect 10838 19570 11058 19600
rect 11174 19570 11394 19600
rect 11510 19570 11730 19600
rect 11846 19570 12066 19600
rect 12182 19570 12402 19600
rect 12518 19570 12738 19600
rect 12854 19570 13074 19600
rect 13190 19570 13410 19600
rect 13526 19570 19474 19600
rect 854 430 19474 19570
rect 854 350 6018 430
rect 6134 350 6354 430
rect 6470 350 6690 430
rect 6806 350 7026 430
rect 7142 350 7362 430
rect 7478 350 7698 430
rect 7814 350 8034 430
rect 8150 350 8370 430
rect 8486 350 8706 430
rect 8822 350 9042 430
rect 9158 350 9378 430
rect 9494 350 9714 430
rect 9830 350 10050 430
rect 10166 350 10386 430
rect 10502 350 10722 430
rect 10838 350 11058 430
rect 11174 350 11394 430
rect 11510 350 11730 430
rect 11846 350 12066 430
rect 12182 350 12402 430
rect 12518 350 12738 430
rect 12854 350 13074 430
rect 13190 350 13410 430
rect 13526 350 13746 430
rect 13862 350 14082 430
rect 14198 350 14418 430
rect 14534 350 14754 430
rect 14870 350 15090 430
rect 15206 350 19474 430
<< metal3 >>
rect 19600 15120 20000 15176
rect 19600 14784 20000 14840
rect 0 14448 400 14504
rect 19600 14448 20000 14504
rect 0 14112 400 14168
rect 19600 14112 20000 14168
rect 0 13776 400 13832
rect 19600 13776 20000 13832
rect 0 13440 400 13496
rect 19600 13440 20000 13496
rect 0 13104 400 13160
rect 19600 13104 20000 13160
rect 0 12768 400 12824
rect 19600 12768 20000 12824
rect 0 12432 400 12488
rect 19600 12432 20000 12488
rect 0 12096 400 12152
rect 19600 12096 20000 12152
rect 0 11760 400 11816
rect 19600 11760 20000 11816
rect 0 11424 400 11480
rect 19600 11424 20000 11480
rect 0 11088 400 11144
rect 19600 11088 20000 11144
rect 0 10752 400 10808
rect 19600 10752 20000 10808
rect 0 10416 400 10472
rect 19600 10416 20000 10472
rect 0 10080 400 10136
rect 19600 10080 20000 10136
rect 0 9744 400 9800
rect 19600 9744 20000 9800
rect 0 9408 400 9464
rect 19600 9408 20000 9464
rect 0 9072 400 9128
rect 19600 9072 20000 9128
rect 0 8736 400 8792
rect 19600 8736 20000 8792
rect 0 8400 400 8456
rect 19600 8400 20000 8456
rect 0 8064 400 8120
rect 19600 8064 20000 8120
rect 0 7728 400 7784
rect 19600 7728 20000 7784
rect 0 7392 400 7448
rect 19600 7392 20000 7448
rect 0 7056 400 7112
rect 19600 7056 20000 7112
rect 0 6720 400 6776
rect 19600 6720 20000 6776
rect 0 6384 400 6440
rect 19600 6384 20000 6440
rect 0 6048 400 6104
rect 19600 6048 20000 6104
rect 0 5712 400 5768
rect 19600 5712 20000 5768
rect 19600 5376 20000 5432
rect 19600 5040 20000 5096
<< obsm3 >>
rect 400 15206 19600 18466
rect 400 15090 19570 15206
rect 400 14870 19600 15090
rect 400 14754 19570 14870
rect 400 14534 19600 14754
rect 430 14418 19570 14534
rect 400 14198 19600 14418
rect 430 14082 19570 14198
rect 400 13862 19600 14082
rect 430 13746 19570 13862
rect 400 13526 19600 13746
rect 430 13410 19570 13526
rect 400 13190 19600 13410
rect 430 13074 19570 13190
rect 400 12854 19600 13074
rect 430 12738 19570 12854
rect 400 12518 19600 12738
rect 430 12402 19570 12518
rect 400 12182 19600 12402
rect 430 12066 19570 12182
rect 400 11846 19600 12066
rect 430 11730 19570 11846
rect 400 11510 19600 11730
rect 430 11394 19570 11510
rect 400 11174 19600 11394
rect 430 11058 19570 11174
rect 400 10838 19600 11058
rect 430 10722 19570 10838
rect 400 10502 19600 10722
rect 430 10386 19570 10502
rect 400 10166 19600 10386
rect 430 10050 19570 10166
rect 400 9830 19600 10050
rect 430 9714 19570 9830
rect 400 9494 19600 9714
rect 430 9378 19570 9494
rect 400 9158 19600 9378
rect 430 9042 19570 9158
rect 400 8822 19600 9042
rect 430 8706 19570 8822
rect 400 8486 19600 8706
rect 430 8370 19570 8486
rect 400 8150 19600 8370
rect 430 8034 19570 8150
rect 400 7814 19600 8034
rect 430 7698 19570 7814
rect 400 7478 19600 7698
rect 430 7362 19570 7478
rect 400 7142 19600 7362
rect 430 7026 19570 7142
rect 400 6806 19600 7026
rect 430 6690 19570 6806
rect 400 6470 19600 6690
rect 430 6354 19570 6470
rect 400 6134 19600 6354
rect 430 6018 19570 6134
rect 400 5798 19600 6018
rect 430 5682 19570 5798
rect 400 5462 19600 5682
rect 400 5346 19570 5462
rect 400 5126 19600 5346
rect 400 5010 19570 5126
rect 400 1554 19600 5010
<< metal4 >>
rect 2923 1538 3083 18454
rect 5254 1538 5414 18454
rect 7585 1538 7745 18454
rect 9916 1538 10076 18454
rect 12247 1538 12407 18454
rect 14578 1538 14738 18454
rect 16909 1538 17069 18454
rect 19240 1538 19400 18454
<< obsm4 >>
rect 10150 2137 10346 7607
<< labels >>
rlabel metal2 s 10080 19600 10136 20000 6 out[0]
port 1 nsew signal output
rlabel metal3 s 0 5712 400 5768 6 out[10]
port 2 nsew signal output
rlabel metal3 s 0 6048 400 6104 6 out[11]
port 3 nsew signal output
rlabel metal2 s 5376 19600 5432 20000 6 out[1]
port 4 nsew signal output
rlabel metal2 s 8064 19600 8120 20000 6 out[2]
port 5 nsew signal output
rlabel metal3 s 0 14448 400 14504 6 out[3]
port 6 nsew signal output
rlabel metal2 s 10416 19600 10472 20000 6 out[4]
port 7 nsew signal output
rlabel metal2 s 6048 0 6104 400 6 out[5]
port 8 nsew signal output
rlabel metal2 s 6384 0 6440 400 6 out[6]
port 9 nsew signal output
rlabel metal2 s 9744 0 9800 400 6 out[7]
port 10 nsew signal output
rlabel metal3 s 0 9408 400 9464 6 out[8]
port 11 nsew signal output
rlabel metal3 s 0 8736 400 8792 6 out[9]
port 12 nsew signal output
rlabel metal3 s 19600 15120 20000 15176 6 proj_out[0]
port 13 nsew signal input
rlabel metal3 s 19600 5040 20000 5096 6 proj_out[10]
port 14 nsew signal input
rlabel metal3 s 19600 6720 20000 6776 6 proj_out[11]
port 15 nsew signal input
rlabel metal3 s 19600 12096 20000 12152 6 proj_out[12]
port 16 nsew signal input
rlabel metal2 s 13440 19600 13496 20000 6 proj_out[13]
port 17 nsew signal input
rlabel metal2 s 12096 19600 12152 20000 6 proj_out[14]
port 18 nsew signal input
rlabel metal3 s 19600 13440 20000 13496 6 proj_out[15]
port 19 nsew signal input
rlabel metal3 s 19600 11088 20000 11144 6 proj_out[16]
port 20 nsew signal input
rlabel metal2 s 15120 0 15176 400 6 proj_out[17]
port 21 nsew signal input
rlabel metal2 s 13104 0 13160 400 6 proj_out[18]
port 22 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 proj_out[19]
port 23 nsew signal input
rlabel metal2 s 13104 19600 13160 20000 6 proj_out[1]
port 24 nsew signal input
rlabel metal3 s 19600 9744 20000 9800 6 proj_out[20]
port 25 nsew signal input
rlabel metal3 s 19600 6384 20000 6440 6 proj_out[21]
port 26 nsew signal input
rlabel metal3 s 19600 6048 20000 6104 6 proj_out[22]
port 27 nsew signal input
rlabel metal3 s 19600 8400 20000 8456 6 proj_out[23]
port 28 nsew signal input
rlabel metal3 s 0 13104 400 13160 6 proj_out[24]
port 29 nsew signal input
rlabel metal2 s 7056 19600 7112 20000 6 proj_out[25]
port 30 nsew signal input
rlabel metal2 s 7392 19600 7448 20000 6 proj_out[26]
port 31 nsew signal input
rlabel metal3 s 0 13440 400 13496 6 proj_out[27]
port 32 nsew signal input
rlabel metal2 s 10752 19600 10808 20000 6 proj_out[28]
port 33 nsew signal input
rlabel metal2 s 10416 0 10472 400 6 proj_out[29]
port 34 nsew signal input
rlabel metal2 s 12768 19600 12824 20000 6 proj_out[2]
port 35 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 proj_out[30]
port 36 nsew signal input
rlabel metal2 s 10752 0 10808 400 6 proj_out[31]
port 37 nsew signal input
rlabel metal3 s 0 7056 400 7112 6 proj_out[32]
port 38 nsew signal input
rlabel metal3 s 0 7392 400 7448 6 proj_out[33]
port 39 nsew signal input
rlabel metal3 s 0 8064 400 8120 6 proj_out[34]
port 40 nsew signal input
rlabel metal3 s 0 7728 400 7784 6 proj_out[35]
port 41 nsew signal input
rlabel metal3 s 0 12768 400 12824 6 proj_out[36]
port 42 nsew signal input
rlabel metal2 s 7728 19600 7784 20000 6 proj_out[37]
port 43 nsew signal input
rlabel metal2 s 6384 19600 6440 20000 6 proj_out[38]
port 44 nsew signal input
rlabel metal3 s 0 12432 400 12488 6 proj_out[39]
port 45 nsew signal input
rlabel metal3 s 19600 14112 20000 14168 6 proj_out[3]
port 46 nsew signal input
rlabel metal3 s 19600 10416 20000 10472 6 proj_out[40]
port 47 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 proj_out[41]
port 48 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 proj_out[42]
port 49 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 proj_out[43]
port 50 nsew signal input
rlabel metal3 s 0 9744 400 9800 6 proj_out[44]
port 51 nsew signal input
rlabel metal3 s 0 6720 400 6776 6 proj_out[45]
port 52 nsew signal input
rlabel metal3 s 0 8400 400 8456 6 proj_out[46]
port 53 nsew signal input
rlabel metal3 s 0 6384 400 6440 6 proj_out[47]
port 54 nsew signal input
rlabel metal3 s 19600 13776 20000 13832 6 proj_out[48]
port 55 nsew signal input
rlabel metal2 s 12432 19600 12488 20000 6 proj_out[49]
port 56 nsew signal input
rlabel metal3 s 19600 10752 20000 10808 6 proj_out[4]
port 57 nsew signal input
rlabel metal2 s 11088 19600 11144 20000 6 proj_out[50]
port 58 nsew signal input
rlabel metal3 s 19600 14448 20000 14504 6 proj_out[51]
port 59 nsew signal input
rlabel metal3 s 19600 11760 20000 11816 6 proj_out[52]
port 60 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 proj_out[53]
port 61 nsew signal input
rlabel metal2 s 11424 0 11480 400 6 proj_out[54]
port 62 nsew signal input
rlabel metal2 s 12096 0 12152 400 6 proj_out[55]
port 63 nsew signal input
rlabel metal3 s 19600 10080 20000 10136 6 proj_out[56]
port 64 nsew signal input
rlabel metal3 s 19600 5712 20000 5768 6 proj_out[57]
port 65 nsew signal input
rlabel metal3 s 19600 5376 20000 5432 6 proj_out[58]
port 66 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 proj_out[59]
port 67 nsew signal input
rlabel metal2 s 13776 0 13832 400 6 proj_out[5]
port 68 nsew signal input
rlabel metal3 s 19600 12768 20000 12824 6 proj_out[60]
port 69 nsew signal input
rlabel metal2 s 11424 19600 11480 20000 6 proj_out[61]
port 70 nsew signal input
rlabel metal2 s 11760 19600 11816 20000 6 proj_out[62]
port 71 nsew signal input
rlabel metal3 s 19600 12432 20000 12488 6 proj_out[63]
port 72 nsew signal input
rlabel metal3 s 19600 14784 20000 14840 6 proj_out[64]
port 73 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 proj_out[65]
port 74 nsew signal input
rlabel metal2 s 14784 0 14840 400 6 proj_out[66]
port 75 nsew signal input
rlabel metal2 s 12432 0 12488 400 6 proj_out[67]
port 76 nsew signal input
rlabel metal3 s 19600 9408 20000 9464 6 proj_out[68]
port 77 nsew signal input
rlabel metal3 s 19600 7728 20000 7784 6 proj_out[69]
port 78 nsew signal input
rlabel metal2 s 13440 0 13496 400 6 proj_out[6]
port 79 nsew signal input
rlabel metal3 s 19600 7392 20000 7448 6 proj_out[70]
port 80 nsew signal input
rlabel metal3 s 19600 8064 20000 8120 6 proj_out[71]
port 81 nsew signal input
rlabel metal2 s 9744 19600 9800 20000 6 proj_out[72]
port 82 nsew signal input
rlabel metal2 s 8400 19600 8456 20000 6 proj_out[73]
port 83 nsew signal input
rlabel metal2 s 5712 19600 5768 20000 6 proj_out[74]
port 84 nsew signal input
rlabel metal3 s 0 13776 400 13832 6 proj_out[75]
port 85 nsew signal input
rlabel metal2 s 9408 19600 9464 20000 6 proj_out[76]
port 86 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 proj_out[77]
port 87 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 proj_out[78]
port 88 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 proj_out[79]
port 89 nsew signal input
rlabel metal2 s 14112 0 14168 400 6 proj_out[7]
port 90 nsew signal input
rlabel metal3 s 0 12096 400 12152 6 proj_out[80]
port 91 nsew signal input
rlabel metal3 s 0 10080 400 10136 6 proj_out[81]
port 92 nsew signal input
rlabel metal3 s 0 9072 400 9128 6 proj_out[82]
port 93 nsew signal input
rlabel metal3 s 0 11088 400 11144 6 proj_out[83]
port 94 nsew signal input
rlabel metal2 s 9072 19600 9128 20000 6 proj_out[84]
port 95 nsew signal input
rlabel metal2 s 6720 19600 6776 20000 6 proj_out[85]
port 96 nsew signal input
rlabel metal2 s 6048 19600 6104 20000 6 proj_out[86]
port 97 nsew signal input
rlabel metal3 s 0 11760 400 11816 6 proj_out[87]
port 98 nsew signal input
rlabel metal2 s 8736 19600 8792 20000 6 proj_out[88]
port 99 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 proj_out[89]
port 100 nsew signal input
rlabel metal3 s 19600 9072 20000 9128 6 proj_out[8]
port 101 nsew signal input
rlabel metal2 s 9408 0 9464 400 6 proj_out[90]
port 102 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 proj_out[91]
port 103 nsew signal input
rlabel metal3 s 0 14112 400 14168 6 proj_out[92]
port 104 nsew signal input
rlabel metal3 s 0 10416 400 10472 6 proj_out[93]
port 105 nsew signal input
rlabel metal3 s 0 10752 400 10808 6 proj_out[94]
port 106 nsew signal input
rlabel metal3 s 0 11424 400 11480 6 proj_out[95]
port 107 nsew signal input
rlabel metal3 s 19600 7056 20000 7112 6 proj_out[9]
port 108 nsew signal input
rlabel metal3 s 19600 11424 20000 11480 6 sel[0]
port 109 nsew signal input
rlabel metal3 s 19600 13104 20000 13160 6 sel[1]
port 110 nsew signal input
rlabel metal3 s 19600 8736 20000 8792 6 sel[2]
port 111 nsew signal input
rlabel metal4 s 2923 1538 3083 18454 6 vdd
port 112 nsew power bidirectional
rlabel metal4 s 7585 1538 7745 18454 6 vdd
port 112 nsew power bidirectional
rlabel metal4 s 12247 1538 12407 18454 6 vdd
port 112 nsew power bidirectional
rlabel metal4 s 16909 1538 17069 18454 6 vdd
port 112 nsew power bidirectional
rlabel metal4 s 5254 1538 5414 18454 6 vss
port 113 nsew ground bidirectional
rlabel metal4 s 9916 1538 10076 18454 6 vss
port 113 nsew ground bidirectional
rlabel metal4 s 14578 1538 14738 18454 6 vss
port 113 nsew ground bidirectional
rlabel metal4 s 19240 1538 19400 18454 6 vss
port 113 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 717866
string GDS_FILE /home/htamas/progs/gfmpw1-multi.v2/openlane/output_mux/runs/23_12_13_05_22/results/signoff/output_mux.magic.gds
string GDS_START 169908
<< end >>

